magic
tech sky130A
magscale 1 2
timestamp 1650815115
<< viali >>
rect 2329 37417 2363 37451
rect 3065 37417 3099 37451
rect 7665 37417 7699 37451
rect 9505 37417 9539 37451
rect 10241 37417 10275 37451
rect 11713 37417 11747 37451
rect 22385 37417 22419 37451
rect 27445 37417 27479 37451
rect 28181 37417 28215 37451
rect 30021 37417 30055 37451
rect 33333 37417 33367 37451
rect 35173 37417 35207 37451
rect 37841 37417 37875 37451
rect 40417 37417 40451 37451
rect 41245 37417 41279 37451
rect 4445 37349 4479 37383
rect 5365 37349 5399 37383
rect 7021 37349 7055 37383
rect 12633 37349 12667 37383
rect 21097 37349 21131 37383
rect 25697 37349 25731 37383
rect 32505 37349 32539 37383
rect 35817 37349 35851 37383
rect 8309 37281 8343 37315
rect 10977 37281 11011 37315
rect 14105 37281 14139 37315
rect 19257 37281 19291 37315
rect 23305 37281 23339 37315
rect 24777 37281 24811 37315
rect 31401 37281 31435 37315
rect 33977 37281 34011 37315
rect 36553 37281 36587 37315
rect 1409 37213 1443 37247
rect 2237 37213 2271 37247
rect 2973 37213 3007 37247
rect 4261 37213 4295 37247
rect 5181 37213 5215 37247
rect 6837 37213 6871 37247
rect 7573 37213 7607 37247
rect 9413 37213 9447 37247
rect 10149 37213 10183 37247
rect 11621 37213 11655 37247
rect 12449 37213 12483 37247
rect 13369 37213 13403 37247
rect 14381 37213 14415 37247
rect 15393 37213 15427 37247
rect 16681 37213 16715 37247
rect 16957 37213 16991 37247
rect 17969 37213 18003 37247
rect 19533 37213 19567 37247
rect 20913 37213 20947 37247
rect 23489 37213 23523 37247
rect 24961 37213 24995 37247
rect 25881 37213 25915 37247
rect 27537 37213 27571 37247
rect 28273 37213 28307 37247
rect 28825 37213 28859 37247
rect 30113 37213 30147 37247
rect 30849 37213 30883 37247
rect 32689 37213 32723 37247
rect 33425 37213 33459 37247
rect 35265 37213 35299 37247
rect 36001 37213 36035 37247
rect 38117 37213 38151 37247
rect 38669 37213 38703 37247
rect 40325 37213 40359 37247
rect 42441 37213 42475 37247
rect 43177 37213 43211 37247
rect 43913 37213 43947 37247
rect 22293 37145 22327 37179
rect 41521 37145 41555 37179
rect 1593 37077 1627 37111
rect 13185 37077 13219 37111
rect 15577 37077 15611 37111
rect 18153 37077 18187 37111
rect 30757 37077 30791 37111
rect 38853 37077 38887 37111
rect 42625 37077 42659 37111
rect 43361 37077 43395 37111
rect 44097 37077 44131 37111
rect 1501 36873 1535 36907
rect 2237 36873 2271 36907
rect 3157 36873 3191 36907
rect 4445 36873 4479 36907
rect 4997 36873 5031 36907
rect 5641 36873 5675 36907
rect 6837 36873 6871 36907
rect 8033 36873 8067 36907
rect 9229 36873 9263 36907
rect 9965 36873 9999 36907
rect 10793 36873 10827 36907
rect 12357 36873 12391 36907
rect 13277 36873 13311 36907
rect 14105 36873 14139 36907
rect 16681 36873 16715 36907
rect 18889 36873 18923 36907
rect 21097 36873 21131 36907
rect 21925 36873 21959 36907
rect 22661 36873 22695 36907
rect 23857 36873 23891 36907
rect 24961 36873 24995 36907
rect 26249 36873 26283 36907
rect 27445 36873 27479 36907
rect 27997 36873 28031 36907
rect 28733 36873 28767 36907
rect 29929 36873 29963 36907
rect 30665 36873 30699 36907
rect 31401 36873 31435 36907
rect 32321 36873 32355 36907
rect 33057 36873 33091 36907
rect 33885 36873 33919 36907
rect 34713 36873 34747 36907
rect 35817 36873 35851 36907
rect 36645 36873 36679 36907
rect 38209 36873 38243 36907
rect 38761 36873 38795 36907
rect 39589 36873 39623 36907
rect 40785 36873 40819 36907
rect 42625 36873 42659 36907
rect 43361 36873 43395 36907
rect 44097 36873 44131 36907
rect 1685 36737 1719 36771
rect 2421 36737 2455 36771
rect 3341 36737 3375 36771
rect 4261 36737 4295 36771
rect 5825 36737 5859 36771
rect 7021 36737 7055 36771
rect 8217 36737 8251 36771
rect 9413 36737 9447 36771
rect 10149 36737 10183 36771
rect 10977 36737 11011 36771
rect 11805 36737 11839 36771
rect 12541 36737 12575 36771
rect 13461 36737 13495 36771
rect 14289 36737 14323 36771
rect 15301 36737 15335 36771
rect 17233 36737 17267 36771
rect 19073 36737 19107 36771
rect 19625 36737 19659 36771
rect 20913 36737 20947 36771
rect 22109 36737 22143 36771
rect 22845 36737 22879 36771
rect 23673 36737 23707 36771
rect 25145 36737 25179 36771
rect 26065 36737 26099 36771
rect 27261 36737 27295 36771
rect 28549 36737 28583 36771
rect 29745 36737 29779 36771
rect 30481 36737 30515 36771
rect 31217 36737 31251 36771
rect 32137 36737 32171 36771
rect 32873 36737 32907 36771
rect 33701 36737 33735 36771
rect 34529 36737 34563 36771
rect 36001 36737 36035 36771
rect 36461 36737 36495 36771
rect 37473 36737 37507 36771
rect 38025 36737 38059 36771
rect 39405 36737 39439 36771
rect 40601 36737 40635 36771
rect 41613 36737 41647 36771
rect 42441 36737 42475 36771
rect 43177 36737 43211 36771
rect 43913 36737 43947 36771
rect 15577 36669 15611 36703
rect 16037 36669 16071 36703
rect 17509 36669 17543 36703
rect 19901 36669 19935 36703
rect 11621 36601 11655 36635
rect 37289 36601 37323 36635
rect 41521 36533 41555 36567
rect 1501 36329 1535 36363
rect 2329 36329 2363 36363
rect 3893 36329 3927 36363
rect 4813 36329 4847 36363
rect 6009 36329 6043 36363
rect 7205 36329 7239 36363
rect 7849 36329 7883 36363
rect 9045 36329 9079 36363
rect 9689 36329 9723 36363
rect 10241 36329 10275 36363
rect 11345 36329 11379 36363
rect 12357 36329 12391 36363
rect 13461 36329 13495 36363
rect 14565 36329 14599 36363
rect 15761 36329 15795 36363
rect 16865 36329 16899 36363
rect 17785 36329 17819 36363
rect 18521 36329 18555 36363
rect 20085 36329 20119 36363
rect 20729 36329 20763 36363
rect 21741 36329 21775 36363
rect 22937 36329 22971 36363
rect 23581 36329 23615 36363
rect 24593 36329 24627 36363
rect 25421 36329 25455 36363
rect 25973 36329 26007 36363
rect 26709 36329 26743 36363
rect 27905 36329 27939 36363
rect 28549 36329 28583 36363
rect 30481 36329 30515 36363
rect 31493 36329 31527 36363
rect 33149 36329 33183 36363
rect 33977 36329 34011 36363
rect 35173 36329 35207 36363
rect 35725 36329 35759 36363
rect 36277 36329 36311 36363
rect 37105 36329 37139 36363
rect 38209 36329 38243 36363
rect 40049 36329 40083 36363
rect 41153 36329 41187 36363
rect 41705 36329 41739 36363
rect 42349 36329 42383 36363
rect 43085 36329 43119 36363
rect 44097 36329 44131 36363
rect 1685 36125 1719 36159
rect 2513 36125 2547 36159
rect 3157 36125 3191 36159
rect 4077 36125 4111 36159
rect 4997 36125 5031 36159
rect 6193 36125 6227 36159
rect 7389 36125 7423 36159
rect 9229 36125 9263 36159
rect 12541 36125 12575 36159
rect 14381 36125 14415 36159
rect 15577 36125 15611 36159
rect 17049 36125 17083 36159
rect 17601 36125 17635 36159
rect 18337 36125 18371 36159
rect 19533 36125 19567 36159
rect 20269 36125 20303 36159
rect 21925 36125 21959 36159
rect 23121 36125 23155 36159
rect 24409 36125 24443 36159
rect 25237 36125 25271 36159
rect 26525 36125 26559 36159
rect 27721 36125 27755 36159
rect 29837 36125 29871 36159
rect 31309 36125 31343 36159
rect 33793 36125 33827 36159
rect 34989 36125 35023 36159
rect 38025 36125 38059 36159
rect 38761 36125 38795 36159
rect 39865 36125 39899 36159
rect 40969 36125 41003 36159
rect 43913 36125 43947 36159
rect 2973 35989 3007 36023
rect 10885 35989 10919 36023
rect 19349 35989 19383 36023
rect 29653 35989 29687 36023
rect 32045 35989 32079 36023
rect 38945 35989 38979 36023
rect 2973 35785 3007 35819
rect 4169 35785 4203 35819
rect 4905 35785 4939 35819
rect 17141 35785 17175 35819
rect 19073 35785 19107 35819
rect 19625 35785 19659 35819
rect 22109 35785 22143 35819
rect 24593 35785 24627 35819
rect 40141 35785 40175 35819
rect 41337 35785 41371 35819
rect 44097 35785 44131 35819
rect 1409 35717 1443 35751
rect 3525 35717 3559 35751
rect 22661 35717 22695 35751
rect 1685 35649 1719 35683
rect 2513 35649 2547 35683
rect 33517 35649 33551 35683
rect 43913 35649 43947 35683
rect 1593 35581 1627 35615
rect 30113 35581 30147 35615
rect 2329 35513 2363 35547
rect 6469 35513 6503 35547
rect 10149 35513 10183 35547
rect 27629 35513 27663 35547
rect 1593 35445 1627 35479
rect 1869 35445 1903 35479
rect 8401 35445 8435 35479
rect 9505 35445 9539 35479
rect 10977 35445 11011 35479
rect 11989 35445 12023 35479
rect 12633 35445 12667 35479
rect 13185 35445 13219 35479
rect 14473 35445 14507 35479
rect 23213 35445 23247 35479
rect 23673 35445 23707 35479
rect 25237 35445 25271 35479
rect 25973 35445 26007 35479
rect 27077 35445 27111 35479
rect 29561 35445 29595 35479
rect 31033 35445 31067 35479
rect 32689 35445 32723 35479
rect 34345 35445 34379 35479
rect 34897 35445 34931 35479
rect 36277 35445 36311 35479
rect 37841 35445 37875 35479
rect 38577 35445 38611 35479
rect 39221 35445 39255 35479
rect 40601 35445 40635 35479
rect 42441 35445 42475 35479
rect 43361 35445 43395 35479
rect 1593 35241 1627 35275
rect 2053 35241 2087 35275
rect 2697 35241 2731 35275
rect 26433 35241 26467 35275
rect 37933 35241 37967 35275
rect 22109 35173 22143 35207
rect 1409 35037 1443 35071
rect 2237 35037 2271 35071
rect 4445 34969 4479 35003
rect 3893 34901 3927 34935
rect 4997 34901 5031 34935
rect 23305 34901 23339 34935
rect 24409 34901 24443 34935
rect 25053 34901 25087 34935
rect 30389 34901 30423 34935
rect 31125 34901 31159 34935
rect 33609 34901 33643 34935
rect 38669 34901 38703 34935
rect 39865 34901 39899 34935
rect 40785 34901 40819 34935
rect 42993 34901 43027 34935
rect 43729 34901 43763 34935
rect 2697 34697 2731 34731
rect 1409 34561 1443 34595
rect 2053 34561 2087 34595
rect 3249 34561 3283 34595
rect 43729 34493 43763 34527
rect 1593 34357 1627 34391
rect 1501 34153 1535 34187
rect 2053 34153 2087 34187
rect 2513 33813 2547 33847
rect 43729 33813 43763 33847
rect 1593 33473 1627 33507
rect 2053 33473 2087 33507
rect 1409 33269 1443 33303
rect 1409 32385 1443 32419
rect 2053 32385 2087 32419
rect 1593 32181 1627 32215
rect 1685 31977 1719 32011
rect 1593 31841 1627 31875
rect 1409 31773 1443 31807
rect 1685 31773 1719 31807
rect 1869 31637 1903 31671
rect 1593 31433 1627 31467
rect 1409 31297 1443 31331
rect 2053 31297 2087 31331
rect 1409 30209 1443 30243
rect 2053 30209 2087 30243
rect 43361 30209 43395 30243
rect 43913 30209 43947 30243
rect 1593 30005 1627 30039
rect 44097 30005 44131 30039
rect 1593 28509 1627 28543
rect 2053 28509 2087 28543
rect 1409 28373 1443 28407
rect 1409 28101 1443 28135
rect 1685 28033 1719 28067
rect 1593 27965 1627 27999
rect 1593 27829 1627 27863
rect 1869 27829 1903 27863
rect 8861 27829 8895 27863
rect 1593 27625 1627 27659
rect 2559 27557 2593 27591
rect 2697 27557 2731 27591
rect 2789 27489 2823 27523
rect 1409 27421 1443 27455
rect 2421 27421 2455 27455
rect 3065 27285 3099 27319
rect 8401 27285 8435 27319
rect 9045 27285 9079 27319
rect 9597 27285 9631 27319
rect 11161 27285 11195 27319
rect 1409 27081 1443 27115
rect 8033 27081 8067 27115
rect 9321 27081 9355 27115
rect 11529 26809 11563 26843
rect 12633 26809 12667 26843
rect 1961 26741 1995 26775
rect 2513 26741 2547 26775
rect 8585 26741 8619 26775
rect 9873 26741 9907 26775
rect 10333 26741 10367 26775
rect 10885 26741 10919 26775
rect 12173 26741 12207 26775
rect 1593 26537 1627 26571
rect 7021 26537 7055 26571
rect 10425 26537 10459 26571
rect 9505 26469 9539 26503
rect 12633 26469 12667 26503
rect 1409 26333 1443 26367
rect 2053 26333 2087 26367
rect 3157 26333 3191 26367
rect 11989 26333 12023 26367
rect 3801 26265 3835 26299
rect 7665 26265 7699 26299
rect 9045 26265 9079 26299
rect 10885 26265 10919 26299
rect 11529 26265 11563 26299
rect 13093 26265 13127 26299
rect 2605 26197 2639 26231
rect 8309 26197 8343 26231
rect 6929 25993 6963 26027
rect 10425 25993 10459 26027
rect 12081 25993 12115 26027
rect 1961 25789 1995 25823
rect 8309 25789 8343 25823
rect 13461 25789 13495 25823
rect 5825 25721 5859 25755
rect 1501 25653 1535 25687
rect 2881 25653 2915 25687
rect 3433 25653 3467 25687
rect 3985 25653 4019 25687
rect 7665 25653 7699 25687
rect 8769 25653 8803 25687
rect 9321 25653 9355 25687
rect 9873 25653 9907 25687
rect 11529 25653 11563 25687
rect 13001 25653 13035 25687
rect 14105 25653 14139 25687
rect 4445 25449 4479 25483
rect 5549 25449 5583 25483
rect 9137 25449 9171 25483
rect 10333 25449 10367 25483
rect 11161 25449 11195 25483
rect 11713 25449 11747 25483
rect 6101 25381 6135 25415
rect 9781 25381 9815 25415
rect 12817 25313 12851 25347
rect 13369 25313 13403 25347
rect 1409 25245 1443 25279
rect 3801 25245 3835 25279
rect 7941 25245 7975 25279
rect 8953 25245 8987 25279
rect 9597 25245 9631 25279
rect 14105 25245 14139 25279
rect 2513 25177 2547 25211
rect 1593 25109 1627 25143
rect 3065 25109 3099 25143
rect 4905 25109 4939 25143
rect 6653 25109 6687 25143
rect 7205 25109 7239 25143
rect 7757 25109 7791 25143
rect 12265 25109 12299 25143
rect 14749 25109 14783 25143
rect 9229 24837 9263 24871
rect 12725 24837 12759 24871
rect 3525 24769 3559 24803
rect 7297 24769 7331 24803
rect 7941 24769 7975 24803
rect 8585 24769 8619 24803
rect 9781 24769 9815 24803
rect 10609 24769 10643 24803
rect 1869 24701 1903 24735
rect 14933 24701 14967 24735
rect 15485 24701 15519 24735
rect 2973 24633 3007 24667
rect 4169 24633 4203 24667
rect 10425 24633 10459 24667
rect 11529 24633 11563 24667
rect 16773 24633 16807 24667
rect 2421 24565 2455 24599
rect 4721 24565 4755 24599
rect 5181 24565 5215 24599
rect 5825 24565 5859 24599
rect 6561 24565 6595 24599
rect 7113 24565 7147 24599
rect 7757 24565 7791 24599
rect 8401 24565 8435 24599
rect 9137 24565 9171 24599
rect 9965 24565 9999 24599
rect 12173 24565 12207 24599
rect 13277 24565 13311 24599
rect 13737 24565 13771 24599
rect 14381 24565 14415 24599
rect 15945 24565 15979 24599
rect 17233 24565 17267 24599
rect 1685 24361 1719 24395
rect 1869 24361 1903 24395
rect 11529 24361 11563 24395
rect 12541 24361 12575 24395
rect 14749 24361 14783 24395
rect 16313 24361 16347 24395
rect 17417 24361 17451 24395
rect 19349 24361 19383 24395
rect 22109 24361 22143 24395
rect 7757 24293 7791 24327
rect 9413 24293 9447 24327
rect 13093 24293 13127 24327
rect 1593 24225 1627 24259
rect 9045 24225 9079 24259
rect 9505 24225 9539 24259
rect 14197 24225 14231 24259
rect 1685 24157 1719 24191
rect 7205 24157 7239 24191
rect 10701 24157 10735 24191
rect 11345 24157 11379 24191
rect 11989 24157 12023 24191
rect 15301 24157 15335 24191
rect 1409 24089 1443 24123
rect 8125 24089 8159 24123
rect 10057 24089 10091 24123
rect 10241 24089 10275 24123
rect 17969 24089 18003 24123
rect 18613 24089 18647 24123
rect 2421 24021 2455 24055
rect 2881 24021 2915 24055
rect 3801 24021 3835 24055
rect 4353 24021 4387 24055
rect 4905 24021 4939 24055
rect 5549 24021 5583 24055
rect 6469 24021 6503 24055
rect 7021 24021 7055 24055
rect 7665 24021 7699 24055
rect 10885 24021 10919 24055
rect 15761 24021 15795 24055
rect 16865 24021 16899 24055
rect 1409 23817 1443 23851
rect 9873 23817 9907 23851
rect 14289 23817 14323 23851
rect 15301 23817 15335 23851
rect 17049 23817 17083 23851
rect 18705 23817 18739 23851
rect 19901 23817 19935 23851
rect 3341 23749 3375 23783
rect 4169 23749 4203 23783
rect 7757 23749 7791 23783
rect 8217 23749 8251 23783
rect 9413 23749 9447 23783
rect 10701 23749 10735 23783
rect 11713 23749 11747 23783
rect 17601 23749 17635 23783
rect 22293 23749 22327 23783
rect 22477 23749 22511 23783
rect 1593 23681 1627 23715
rect 5825 23681 5859 23715
rect 6837 23681 6871 23715
rect 8493 23681 8527 23715
rect 10517 23681 10551 23715
rect 10793 23681 10827 23715
rect 12265 23681 12299 23715
rect 13093 23681 13127 23715
rect 13553 23681 13587 23715
rect 32597 23681 32631 23715
rect 8309 23613 8343 23647
rect 2329 23545 2363 23579
rect 4721 23545 4755 23579
rect 5641 23545 5675 23579
rect 7297 23545 7331 23579
rect 7481 23545 7515 23579
rect 9781 23545 9815 23579
rect 10517 23545 10551 23579
rect 11529 23545 11563 23579
rect 12909 23545 12943 23579
rect 2881 23477 2915 23511
rect 6653 23477 6687 23511
rect 8309 23477 8343 23511
rect 8677 23477 8711 23511
rect 12449 23477 12483 23511
rect 13737 23477 13771 23511
rect 15853 23477 15887 23511
rect 18245 23477 18279 23511
rect 19349 23477 19383 23511
rect 32689 23477 32723 23511
rect 1593 23273 1627 23307
rect 3249 23273 3283 23307
rect 5641 23273 5675 23307
rect 9137 23273 9171 23307
rect 11253 23273 11287 23307
rect 15577 23273 15611 23307
rect 16773 23273 16807 23307
rect 17601 23273 17635 23307
rect 18613 23273 18647 23307
rect 20729 23273 20763 23307
rect 6469 23205 6503 23239
rect 8953 23205 8987 23239
rect 10241 23205 10275 23239
rect 11069 23205 11103 23239
rect 11713 23205 11747 23239
rect 18061 23205 18095 23239
rect 21557 23205 21591 23239
rect 28733 23205 28767 23239
rect 3893 23137 3927 23171
rect 7757 23137 7791 23171
rect 9229 23137 9263 23171
rect 9873 23137 9907 23171
rect 10793 23137 10827 23171
rect 19257 23137 19291 23171
rect 19533 23137 19567 23171
rect 30205 23137 30239 23171
rect 1409 23069 1443 23103
rect 5181 23069 5215 23103
rect 5825 23069 5859 23103
rect 7573 23069 7607 23103
rect 9137 23069 9171 23103
rect 11989 23069 12023 23103
rect 12633 23069 12667 23103
rect 13185 23069 13219 23103
rect 14105 23069 14139 23103
rect 17417 23069 17451 23103
rect 30941 23069 30975 23103
rect 4445 23001 4479 23035
rect 6745 23001 6779 23035
rect 9413 23001 9447 23035
rect 11713 23001 11747 23035
rect 12449 23001 12483 23035
rect 14749 23001 14783 23035
rect 20637 23001 20671 23035
rect 21373 23001 21407 23035
rect 22109 23001 22143 23035
rect 28549 23001 28583 23035
rect 30021 23001 30055 23035
rect 30757 23001 30791 23035
rect 31493 23001 31527 23035
rect 31677 23001 31711 23035
rect 2145 22933 2179 22967
rect 2697 22933 2731 22967
rect 4997 22933 5031 22967
rect 6285 22933 6319 22967
rect 7205 22933 7239 22967
rect 7665 22933 7699 22967
rect 10333 22933 10367 22967
rect 11897 22933 11931 22967
rect 13369 22933 13403 22967
rect 14289 22933 14323 22967
rect 16313 22933 16347 22967
rect 22201 22933 22235 22967
rect 27997 22933 28031 22967
rect 32321 22933 32355 22967
rect 2697 22729 2731 22763
rect 3525 22729 3559 22763
rect 4721 22729 4755 22763
rect 5825 22729 5859 22763
rect 7573 22729 7607 22763
rect 11989 22729 12023 22763
rect 12541 22729 12575 22763
rect 14841 22729 14875 22763
rect 15853 22729 15887 22763
rect 22385 22729 22419 22763
rect 29837 22729 29871 22763
rect 7113 22661 7147 22695
rect 10977 22661 11011 22695
rect 11529 22661 11563 22695
rect 12725 22661 12759 22695
rect 14013 22661 14047 22695
rect 16773 22661 16807 22695
rect 21189 22661 21223 22695
rect 22293 22661 22327 22695
rect 1593 22593 1627 22627
rect 2053 22593 2087 22627
rect 2881 22593 2915 22627
rect 4261 22593 4295 22627
rect 4905 22593 4939 22627
rect 7205 22593 7239 22627
rect 8585 22593 8619 22627
rect 8861 22593 8895 22627
rect 10149 22593 10183 22627
rect 10609 22593 10643 22627
rect 10793 22593 10827 22627
rect 12449 22593 12483 22627
rect 13461 22593 13495 22627
rect 14657 22593 14691 22627
rect 15301 22593 15335 22627
rect 17877 22593 17911 22627
rect 19165 22593 19199 22627
rect 19441 22593 19475 22627
rect 20177 22593 20211 22627
rect 5365 22525 5399 22559
rect 6929 22525 6963 22559
rect 13185 22525 13219 22559
rect 13369 22525 13403 22559
rect 18153 22525 18187 22559
rect 19901 22525 19935 22559
rect 5733 22457 5767 22491
rect 9919 22457 9953 22491
rect 11897 22457 11931 22491
rect 14197 22457 14231 22491
rect 1409 22389 1443 22423
rect 4077 22389 4111 22423
rect 12725 22389 12759 22423
rect 13461 22389 13495 22423
rect 30573 22389 30607 22423
rect 31309 22389 31343 22423
rect 6929 22185 6963 22219
rect 10977 22185 11011 22219
rect 22109 22185 22143 22219
rect 4629 22117 4663 22151
rect 5641 22117 5675 22151
rect 11713 22117 11747 22151
rect 12725 22117 12759 22151
rect 3801 22049 3835 22083
rect 4813 22049 4847 22083
rect 5733 22049 5767 22083
rect 6285 22049 6319 22083
rect 10333 22049 10367 22083
rect 15393 22049 15427 22083
rect 18521 22049 18555 22083
rect 19533 22049 19567 22083
rect 20545 22049 20579 22083
rect 1409 21981 1443 22015
rect 2237 21981 2271 22015
rect 2881 21981 2915 22015
rect 7941 21981 7975 22015
rect 8217 21981 8251 22015
rect 9505 21981 9539 22015
rect 9781 21981 9815 22015
rect 12357 21981 12391 22015
rect 13277 21981 13311 22015
rect 13369 21981 13403 22015
rect 14105 21981 14139 22015
rect 14289 21981 14323 22015
rect 15669 21981 15703 22015
rect 16865 21981 16899 22015
rect 17141 21981 17175 22015
rect 20821 21981 20855 22015
rect 4353 21913 4387 21947
rect 5273 21913 5307 21947
rect 11437 21913 11471 21947
rect 13553 21913 13587 21947
rect 18337 21913 18371 21947
rect 19349 21913 19383 21947
rect 21281 21913 21315 21947
rect 1593 21845 1627 21879
rect 2053 21845 2087 21879
rect 2697 21845 2731 21879
rect 6469 21845 6503 21879
rect 6561 21845 6595 21879
rect 10517 21845 10551 21879
rect 10609 21845 10643 21879
rect 11897 21845 11931 21879
rect 12817 21845 12851 21879
rect 13277 21845 13311 21879
rect 17601 21845 17635 21879
rect 1685 21641 1719 21675
rect 2973 21641 3007 21675
rect 13185 21641 13219 21675
rect 27721 21641 27755 21675
rect 6469 21573 6503 21607
rect 6653 21573 6687 21607
rect 8861 21573 8895 21607
rect 13645 21573 13679 21607
rect 22937 21573 22971 21607
rect 1501 21505 1535 21539
rect 2329 21505 2363 21539
rect 2789 21505 2823 21539
rect 3525 21505 3559 21539
rect 3709 21505 3743 21539
rect 5457 21505 5491 21539
rect 9505 21505 9539 21539
rect 10977 21505 11011 21539
rect 11897 21505 11931 21539
rect 13829 21505 13863 21539
rect 15485 21505 15519 21539
rect 16957 21505 16991 21539
rect 19073 21505 19107 21539
rect 20637 21505 20671 21539
rect 4169 21437 4203 21471
rect 4629 21437 4663 21471
rect 5549 21437 5583 21471
rect 5641 21437 5675 21471
rect 8033 21437 8067 21471
rect 9045 21437 9079 21471
rect 11989 21437 12023 21471
rect 12081 21437 12115 21471
rect 12725 21437 12759 21471
rect 15761 21437 15795 21471
rect 16681 21437 16715 21471
rect 20913 21437 20947 21471
rect 2145 21369 2179 21403
rect 4353 21369 4387 21403
rect 11529 21369 11563 21403
rect 13093 21369 13127 21403
rect 5089 21301 5123 21335
rect 9735 21301 9769 21335
rect 10793 21301 10827 21335
rect 14381 21301 14415 21335
rect 18061 21301 18095 21335
rect 18521 21301 18555 21335
rect 21833 21301 21867 21335
rect 22385 21301 22419 21335
rect 23489 21301 23523 21335
rect 24133 21301 24167 21335
rect 3249 21097 3283 21131
rect 4537 21097 4571 21131
rect 8401 21097 8435 21131
rect 13277 21097 13311 21131
rect 15853 21097 15887 21131
rect 25237 21097 25271 21131
rect 26617 21097 26651 21131
rect 28089 21097 28123 21131
rect 1685 21029 1719 21063
rect 2329 21029 2363 21063
rect 3157 21029 3191 21063
rect 15669 21029 15703 21063
rect 16589 21029 16623 21063
rect 17509 21029 17543 21063
rect 17693 21029 17727 21063
rect 18153 21029 18187 21063
rect 27537 21029 27571 21063
rect 4997 20961 5031 20995
rect 5181 20961 5215 20995
rect 6285 20961 6319 20995
rect 11805 20961 11839 20995
rect 12725 20961 12759 20995
rect 14657 20961 14691 20995
rect 14933 20961 14967 20995
rect 16313 20961 16347 20995
rect 16773 20961 16807 20995
rect 27169 20961 27203 20995
rect 27629 20961 27663 20995
rect 1501 20893 1535 20927
rect 2145 20893 2179 20927
rect 6561 20893 6595 20927
rect 7021 20893 7055 20927
rect 8953 20893 8987 20927
rect 10793 20893 10827 20927
rect 12081 20893 12115 20927
rect 12817 20893 12851 20927
rect 12909 20893 12943 20927
rect 18337 20893 18371 20927
rect 20361 20893 20395 20927
rect 2789 20825 2823 20859
rect 3801 20825 3835 20859
rect 3985 20825 4019 20859
rect 4905 20825 4939 20859
rect 7288 20825 7322 20859
rect 9137 20825 9171 20859
rect 15393 20825 15427 20859
rect 17233 20825 17267 20859
rect 19349 20825 19383 20859
rect 23121 20825 23155 20859
rect 19901 20757 19935 20791
rect 20913 20757 20947 20791
rect 21465 20757 21499 20791
rect 22109 20757 22143 20791
rect 22661 20757 22695 20791
rect 23673 20757 23707 20791
rect 24501 20757 24535 20791
rect 29561 20757 29595 20791
rect 3249 20553 3283 20587
rect 6561 20553 6595 20587
rect 18981 20553 19015 20587
rect 20453 20553 20487 20587
rect 21005 20553 21039 20587
rect 22661 20553 22695 20587
rect 24225 20553 24259 20587
rect 25789 20553 25823 20587
rect 28365 20553 28399 20587
rect 29745 20553 29779 20587
rect 2145 20485 2179 20519
rect 15669 20485 15703 20519
rect 17601 20485 17635 20519
rect 18521 20485 18555 20519
rect 19441 20485 19475 20519
rect 22753 20485 22787 20519
rect 24961 20485 24995 20519
rect 27537 20485 27571 20519
rect 1409 20417 1443 20451
rect 4261 20417 4295 20451
rect 5549 20417 5583 20451
rect 5825 20417 5859 20451
rect 6653 20417 6687 20451
rect 9781 20417 9815 20451
rect 10977 20417 11011 20451
rect 13461 20417 13495 20451
rect 14933 20417 14967 20451
rect 24133 20417 24167 20451
rect 25697 20417 25731 20451
rect 28917 20417 28951 20451
rect 29101 20417 29135 20451
rect 2789 20349 2823 20383
rect 4537 20349 4571 20383
rect 7205 20349 7239 20383
rect 8861 20349 8895 20383
rect 9045 20349 9079 20383
rect 9505 20349 9539 20383
rect 12081 20349 12115 20383
rect 12357 20349 12391 20383
rect 13737 20349 13771 20383
rect 15209 20349 15243 20383
rect 2329 20281 2363 20315
rect 3157 20281 3191 20315
rect 10793 20281 10827 20315
rect 16037 20281 16071 20315
rect 17325 20281 17359 20315
rect 18245 20281 18279 20315
rect 19165 20281 19199 20315
rect 21833 20281 21867 20315
rect 1593 20213 1627 20247
rect 16129 20213 16163 20247
rect 17141 20213 17175 20247
rect 18061 20213 18095 20247
rect 19901 20213 19935 20247
rect 23305 20213 23339 20247
rect 24869 20213 24903 20247
rect 27445 20213 27479 20247
rect 33609 20213 33643 20247
rect 2053 20009 2087 20043
rect 3249 20009 3283 20043
rect 18705 20009 18739 20043
rect 25697 20009 25731 20043
rect 32781 20009 32815 20043
rect 1961 19941 1995 19975
rect 16957 19941 16991 19975
rect 17969 19941 18003 19975
rect 19901 19941 19935 19975
rect 27077 19941 27111 19975
rect 30665 19941 30699 19975
rect 36093 19941 36127 19975
rect 1593 19873 1627 19907
rect 2697 19873 2731 19907
rect 4537 19873 4571 19907
rect 5825 19873 5859 19907
rect 7297 19873 7331 19907
rect 10793 19873 10827 19907
rect 11805 19873 11839 19907
rect 13277 19873 13311 19907
rect 14381 19873 14415 19907
rect 15945 19873 15979 19907
rect 16221 19873 16255 19907
rect 20913 19873 20947 19907
rect 22201 19873 22235 19907
rect 27813 19873 27847 19907
rect 35357 19873 35391 19907
rect 4813 19805 4847 19839
rect 6101 19805 6135 19839
rect 6561 19805 6595 19839
rect 8953 19805 8987 19839
rect 12081 19805 12115 19839
rect 13553 19805 13587 19839
rect 14105 19805 14139 19839
rect 19717 19805 19751 19839
rect 20637 19805 20671 19839
rect 21925 19805 21959 19839
rect 23305 19805 23339 19839
rect 24869 19805 24903 19839
rect 26249 19805 26283 19839
rect 28549 19805 28583 19839
rect 30021 19805 30055 19839
rect 33977 19805 34011 19839
rect 2789 19737 2823 19771
rect 6745 19737 6779 19771
rect 9137 19737 9171 19771
rect 17233 19737 17267 19771
rect 17693 19737 17727 19771
rect 23489 19737 23523 19771
rect 25053 19737 25087 19771
rect 25605 19737 25639 19771
rect 26893 19737 26927 19771
rect 27629 19737 27663 19771
rect 30205 19737 30239 19771
rect 30849 19737 30883 19771
rect 32689 19737 32723 19771
rect 33793 19737 33827 19771
rect 35173 19737 35207 19771
rect 35909 19737 35943 19771
rect 2881 19669 2915 19703
rect 16773 19669 16807 19703
rect 18153 19669 18187 19703
rect 28641 19669 28675 19703
rect 31401 19669 31435 19703
rect 32045 19669 32079 19703
rect 2053 19465 2087 19499
rect 2513 19465 2547 19499
rect 3985 19465 4019 19499
rect 5825 19465 5859 19499
rect 13967 19465 14001 19499
rect 18613 19465 18647 19499
rect 19717 19465 19751 19499
rect 28733 19465 28767 19499
rect 29469 19465 29503 19499
rect 33149 19465 33183 19499
rect 4712 19397 4746 19431
rect 8493 19397 8527 19431
rect 9137 19397 9171 19431
rect 10793 19397 10827 19431
rect 20269 19397 20303 19431
rect 21097 19397 21131 19431
rect 25329 19397 25363 19431
rect 26065 19397 26099 19431
rect 1409 19329 1443 19363
rect 2421 19329 2455 19363
rect 3617 19329 3651 19363
rect 4445 19329 4479 19363
rect 6837 19329 6871 19363
rect 8677 19329 8711 19363
rect 10977 19329 11011 19363
rect 11796 19329 11830 19363
rect 15209 19329 15243 19363
rect 15945 19329 15979 19363
rect 16681 19329 16715 19363
rect 16948 19329 16982 19363
rect 18797 19329 18831 19363
rect 22109 19329 22143 19363
rect 24593 19329 24627 19363
rect 27445 19329 27479 19363
rect 28181 19329 28215 19363
rect 28825 19329 28859 19363
rect 29561 19329 29595 19363
rect 33057 19329 33091 19363
rect 34253 19329 34287 19363
rect 2697 19261 2731 19295
rect 3341 19261 3375 19295
rect 3525 19261 3559 19295
rect 11529 19261 11563 19295
rect 14197 19261 14231 19295
rect 15485 19261 15519 19295
rect 19257 19261 19291 19295
rect 20453 19261 20487 19295
rect 21833 19261 21867 19295
rect 23213 19261 23247 19295
rect 25513 19261 25547 19295
rect 26249 19261 26283 19295
rect 34437 19261 34471 19295
rect 16129 19193 16163 19227
rect 18061 19193 18095 19227
rect 19533 19193 19567 19227
rect 23765 19193 23799 19227
rect 27629 19193 27663 19227
rect 1593 19125 1627 19159
rect 12909 19125 12943 19159
rect 21005 19125 21039 19159
rect 24685 19125 24719 19159
rect 30205 19125 30239 19159
rect 32413 19125 32447 19159
rect 34897 19125 34931 19159
rect 35633 19125 35667 19159
rect 2053 18921 2087 18955
rect 3249 18921 3283 18955
rect 21557 18921 21591 18955
rect 22201 18921 22235 18955
rect 24409 18921 24443 18955
rect 24961 18921 24995 18955
rect 27261 18921 27295 18955
rect 18153 18853 18187 18887
rect 19625 18853 19659 18887
rect 20453 18853 20487 18887
rect 1869 18785 1903 18819
rect 2697 18785 2731 18819
rect 2789 18785 2823 18819
rect 6101 18785 6135 18819
rect 6561 18785 6595 18819
rect 8217 18785 8251 18819
rect 10609 18785 10643 18819
rect 11713 18785 11747 18819
rect 14105 18785 14139 18819
rect 15945 18785 15979 18819
rect 16221 18785 16255 18819
rect 16865 18785 16899 18819
rect 19717 18785 19751 18819
rect 1777 18717 1811 18751
rect 2053 18717 2087 18751
rect 2881 18717 2915 18751
rect 4261 18717 4295 18751
rect 8401 18717 8435 18751
rect 11253 18717 11287 18751
rect 14381 18717 14415 18751
rect 20269 18717 20303 18751
rect 21097 18717 21131 18751
rect 21741 18717 21775 18751
rect 22385 18717 22419 18751
rect 23029 18717 23063 18751
rect 5917 18649 5951 18683
rect 11069 18649 11103 18683
rect 11980 18649 12014 18683
rect 17877 18649 17911 18683
rect 19257 18649 19291 18683
rect 25605 18649 25639 18683
rect 27169 18649 27203 18683
rect 1593 18581 1627 18615
rect 13093 18581 13127 18615
rect 16957 18581 16991 18615
rect 17049 18581 17083 18615
rect 17417 18581 17451 18615
rect 18337 18581 18371 18615
rect 20913 18581 20947 18615
rect 22845 18581 22879 18615
rect 23581 18581 23615 18615
rect 26617 18581 26651 18615
rect 33977 18581 34011 18615
rect 2329 18377 2363 18411
rect 16037 18377 16071 18411
rect 16681 18377 16715 18411
rect 18245 18377 18279 18411
rect 22385 18377 22419 18411
rect 22937 18377 22971 18411
rect 23581 18377 23615 18411
rect 24777 18377 24811 18411
rect 25789 18377 25823 18411
rect 29285 18377 29319 18411
rect 4712 18309 4746 18343
rect 8309 18309 8343 18343
rect 21189 18309 21223 18343
rect 22293 18309 22327 18343
rect 28365 18309 28399 18343
rect 29193 18309 29227 18343
rect 30205 18309 30239 18343
rect 3709 18241 3743 18275
rect 3985 18241 4019 18275
rect 4445 18241 4479 18275
rect 11529 18241 11563 18275
rect 14105 18241 14139 18275
rect 14372 18241 14406 18275
rect 17049 18241 17083 18275
rect 17141 18241 17175 18275
rect 18337 18241 18371 18275
rect 19993 18241 20027 18275
rect 20913 18241 20947 18275
rect 21005 18241 21039 18275
rect 23121 18241 23155 18275
rect 24225 18241 24259 18275
rect 25329 18241 25363 18275
rect 27629 18241 27663 18275
rect 28181 18241 28215 18275
rect 30021 18241 30055 18275
rect 2145 18173 2179 18207
rect 2237 18173 2271 18207
rect 6929 18173 6963 18207
rect 8493 18173 8527 18207
rect 9045 18173 9079 18207
rect 10609 18173 10643 18207
rect 10793 18173 10827 18207
rect 11713 18173 11747 18207
rect 12449 18173 12483 18207
rect 17233 18173 17267 18207
rect 18429 18173 18463 18207
rect 19533 18173 19567 18207
rect 20453 18173 20487 18207
rect 26341 18173 26375 18207
rect 5825 18105 5859 18139
rect 19165 18105 19199 18139
rect 20361 18105 20395 18139
rect 1501 18037 1535 18071
rect 2697 18037 2731 18071
rect 15485 18037 15519 18071
rect 17877 18037 17911 18071
rect 19073 18037 19107 18071
rect 21189 18037 21223 18071
rect 27077 18037 27111 18071
rect 1593 17833 1627 17867
rect 3801 17833 3835 17867
rect 17141 17833 17175 17867
rect 18521 17833 18555 17867
rect 20913 17833 20947 17867
rect 24409 17833 24443 17867
rect 25605 17833 25639 17867
rect 26065 17833 26099 17867
rect 27813 17833 27847 17867
rect 28273 17833 28307 17867
rect 6101 17765 6135 17799
rect 15485 17765 15519 17799
rect 19625 17765 19659 17799
rect 20177 17765 20211 17799
rect 21649 17765 21683 17799
rect 22569 17765 22603 17799
rect 23489 17765 23523 17799
rect 1593 17697 1627 17731
rect 2973 17697 3007 17731
rect 3893 17697 3927 17731
rect 4721 17697 4755 17731
rect 6561 17697 6595 17731
rect 7021 17697 7055 17731
rect 12449 17697 12483 17731
rect 12909 17697 12943 17731
rect 14105 17697 14139 17731
rect 16129 17697 16163 17731
rect 17785 17697 17819 17731
rect 22385 17697 22419 17731
rect 23305 17697 23339 17731
rect 1409 17629 1443 17663
rect 1685 17629 1719 17663
rect 3249 17629 3283 17663
rect 4077 17629 4111 17663
rect 10793 17629 10827 17663
rect 13093 17629 13127 17663
rect 14361 17629 14395 17663
rect 20177 17629 20211 17663
rect 20453 17629 20487 17663
rect 21189 17629 21223 17663
rect 21833 17629 21867 17663
rect 26617 17629 26651 17663
rect 27169 17629 27203 17663
rect 3801 17561 3835 17595
rect 4988 17561 5022 17595
rect 6745 17561 6779 17595
rect 8953 17561 8987 17595
rect 10609 17561 10643 17595
rect 16313 17561 16347 17595
rect 18505 17561 18539 17595
rect 18705 17561 18739 17595
rect 19257 17561 19291 17595
rect 20913 17561 20947 17595
rect 22845 17561 22879 17595
rect 23765 17561 23799 17595
rect 1869 17493 1903 17527
rect 4261 17493 4295 17527
rect 16221 17493 16255 17527
rect 16681 17493 16715 17527
rect 17509 17493 17543 17527
rect 17601 17493 17635 17527
rect 18337 17493 18371 17527
rect 19717 17493 19751 17527
rect 20361 17493 20395 17527
rect 21097 17493 21131 17527
rect 24961 17493 24995 17527
rect 29009 17493 29043 17527
rect 29837 17493 29871 17527
rect 1777 17289 1811 17323
rect 3985 17289 4019 17323
rect 5825 17289 5859 17323
rect 23121 17289 23155 17323
rect 2872 17221 2906 17255
rect 4690 17221 4724 17255
rect 9137 17221 9171 17255
rect 10793 17221 10827 17255
rect 11529 17221 11563 17255
rect 13185 17221 13219 17255
rect 14350 17221 14384 17255
rect 18429 17221 18463 17255
rect 19349 17221 19383 17255
rect 20637 17221 20671 17255
rect 26157 17221 26191 17255
rect 28089 17221 28123 17255
rect 1685 17153 1719 17187
rect 2605 17153 2639 17187
rect 4445 17153 4479 17187
rect 6469 17153 6503 17187
rect 7113 17153 7147 17187
rect 7380 17153 7414 17187
rect 14105 17153 14139 17187
rect 16681 17153 16715 17187
rect 16957 17153 16991 17187
rect 18113 17153 18147 17187
rect 18245 17153 18279 17187
rect 19073 17153 19107 17187
rect 21281 17153 21315 17187
rect 22017 17153 22051 17187
rect 22109 17153 22143 17187
rect 22293 17153 22327 17187
rect 28641 17153 28675 17187
rect 1501 17085 1535 17119
rect 8953 17085 8987 17119
rect 13369 17085 13403 17119
rect 16037 17085 16071 17119
rect 19257 17085 19291 17119
rect 20177 17085 20211 17119
rect 23581 17085 23615 17119
rect 24685 17085 24719 17119
rect 25605 17085 25639 17119
rect 2145 17017 2179 17051
rect 8493 17017 8527 17051
rect 17969 17017 18003 17051
rect 18889 17017 18923 17051
rect 20269 17017 20303 17051
rect 21097 17017 21131 17051
rect 23305 17017 23339 17051
rect 25053 17017 25087 17051
rect 6561 16949 6595 16983
rect 15485 16949 15519 16983
rect 18429 16949 18463 16983
rect 19349 16949 19383 16983
rect 22293 16949 22327 16983
rect 24041 16949 24075 16983
rect 25145 16949 25179 16983
rect 26985 16949 27019 16983
rect 27629 16949 27663 16983
rect 1777 16745 1811 16779
rect 19441 16745 19475 16779
rect 20637 16745 20671 16779
rect 25881 16745 25915 16779
rect 28181 16745 28215 16779
rect 28641 16745 28675 16779
rect 1961 16677 1995 16711
rect 14197 16677 14231 16711
rect 21373 16677 21407 16711
rect 22385 16677 22419 16711
rect 23489 16677 23523 16711
rect 25421 16677 25455 16711
rect 27077 16677 27111 16711
rect 29561 16677 29595 16711
rect 1685 16609 1719 16643
rect 2421 16609 2455 16643
rect 4353 16609 4387 16643
rect 6469 16609 6503 16643
rect 6929 16609 6963 16643
rect 9045 16609 9079 16643
rect 9781 16609 9815 16643
rect 11345 16609 11379 16643
rect 11805 16609 11839 16643
rect 14657 16609 14691 16643
rect 16589 16609 16623 16643
rect 16865 16609 16899 16643
rect 17877 16609 17911 16643
rect 18153 16609 18187 16643
rect 19625 16609 19659 16643
rect 20453 16609 20487 16643
rect 21557 16609 21591 16643
rect 24501 16609 24535 16643
rect 27629 16609 27663 16643
rect 1777 16541 1811 16575
rect 4629 16541 4663 16575
rect 6213 16541 6247 16575
rect 7196 16541 7230 16575
rect 12081 16541 12115 16575
rect 14924 16541 14958 16575
rect 19441 16541 19475 16575
rect 19717 16541 19751 16575
rect 20361 16541 20395 16575
rect 23305 16541 23339 16575
rect 1501 16473 1535 16507
rect 11161 16473 11195 16507
rect 20637 16473 20671 16507
rect 21097 16473 21131 16507
rect 22017 16473 22051 16507
rect 25237 16473 25271 16507
rect 2651 16405 2685 16439
rect 5089 16405 5123 16439
rect 8309 16405 8343 16439
rect 13185 16405 13219 16439
rect 16037 16405 16071 16439
rect 19257 16405 19291 16439
rect 20177 16405 20211 16439
rect 22477 16405 22511 16439
rect 26433 16405 26467 16439
rect 1685 16201 1719 16235
rect 2145 16201 2179 16235
rect 3985 16201 4019 16235
rect 11621 16201 11655 16235
rect 15761 16201 15795 16235
rect 16681 16201 16715 16235
rect 21833 16201 21867 16235
rect 23673 16201 23707 16235
rect 25053 16201 25087 16235
rect 25605 16201 25639 16235
rect 27629 16201 27663 16235
rect 30389 16201 30423 16235
rect 2850 16133 2884 16167
rect 12756 16133 12790 16167
rect 17794 16133 17828 16167
rect 20177 16133 20211 16167
rect 23213 16133 23247 16167
rect 26157 16133 26191 16167
rect 1777 16065 1811 16099
rect 2605 16065 2639 16099
rect 4445 16065 4479 16099
rect 4712 16065 4746 16099
rect 6469 16065 6503 16099
rect 6561 16065 6595 16099
rect 8421 16065 8455 16099
rect 8677 16065 8711 16099
rect 9137 16065 9171 16099
rect 13001 16065 13035 16099
rect 14677 16065 14711 16099
rect 14933 16065 14967 16099
rect 15669 16065 15703 16099
rect 18061 16065 18095 16099
rect 18889 16065 18923 16099
rect 19901 16065 19935 16099
rect 19993 16065 20027 16099
rect 20821 16065 20855 16099
rect 23857 16065 23891 16099
rect 24501 16065 24535 16099
rect 26985 16065 27019 16099
rect 1593 15997 1627 16031
rect 10793 15997 10827 16031
rect 10977 15997 11011 16031
rect 15485 15997 15519 16031
rect 18613 15997 18647 16031
rect 18797 15997 18831 16031
rect 20637 15997 20671 16031
rect 21097 15997 21131 16031
rect 22293 15997 22327 16031
rect 22753 15997 22787 16031
rect 29193 15997 29227 16031
rect 5825 15929 5859 15963
rect 16129 15929 16163 15963
rect 19257 15929 19291 15963
rect 19717 15929 19751 15963
rect 21925 15929 21959 15963
rect 22937 15929 22971 15963
rect 24317 15929 24351 15963
rect 29745 15929 29779 15963
rect 6745 15861 6779 15895
rect 7297 15861 7331 15895
rect 13553 15861 13587 15895
rect 20177 15861 20211 15895
rect 21005 15861 21039 15895
rect 28089 15861 28123 15895
rect 28641 15861 28675 15895
rect 1777 15657 1811 15691
rect 14197 15657 14231 15691
rect 19717 15657 19751 15691
rect 20637 15657 20671 15691
rect 21373 15657 21407 15691
rect 21557 15657 21591 15691
rect 23673 15657 23707 15691
rect 25789 15657 25823 15691
rect 26341 15657 26375 15691
rect 26801 15657 26835 15691
rect 27353 15657 27387 15691
rect 29561 15657 29595 15691
rect 30113 15657 30147 15691
rect 1961 15589 1995 15623
rect 8309 15589 8343 15623
rect 19257 15589 19291 15623
rect 22293 15589 22327 15623
rect 22937 15589 22971 15623
rect 24409 15589 24443 15623
rect 1593 15521 1627 15555
rect 2421 15521 2455 15555
rect 4629 15521 4663 15555
rect 9229 15521 9263 15555
rect 10885 15521 10919 15555
rect 11069 15521 11103 15555
rect 13277 15521 13311 15555
rect 17877 15521 17911 15555
rect 19625 15521 19659 15555
rect 21281 15521 21315 15555
rect 22477 15521 22511 15555
rect 27905 15521 27939 15555
rect 1777 15453 1811 15487
rect 2697 15453 2731 15487
rect 4353 15453 4387 15487
rect 5089 15453 5123 15487
rect 6929 15453 6963 15487
rect 7196 15453 7230 15487
rect 11529 15453 11563 15487
rect 15577 15453 15611 15487
rect 16037 15453 16071 15487
rect 18153 15453 18187 15487
rect 19441 15453 19475 15487
rect 20361 15453 20395 15487
rect 20453 15453 20487 15487
rect 21373 15453 21407 15487
rect 23213 15453 23247 15487
rect 23857 15453 23891 15487
rect 24593 15453 24627 15487
rect 25237 15453 25271 15487
rect 1501 15385 1535 15419
rect 5356 15385 5390 15419
rect 15332 15385 15366 15419
rect 16282 15385 16316 15419
rect 19717 15385 19751 15419
rect 20637 15385 20671 15419
rect 21097 15385 21131 15419
rect 22017 15385 22051 15419
rect 22937 15385 22971 15419
rect 23121 15385 23155 15419
rect 6469 15317 6503 15351
rect 17417 15317 17451 15351
rect 20177 15317 20211 15351
rect 25053 15317 25087 15351
rect 28457 15317 28491 15351
rect 20177 15113 20211 15147
rect 21189 15113 21223 15147
rect 25697 15113 25731 15147
rect 26341 15113 26375 15147
rect 26985 15113 27019 15147
rect 30389 15113 30423 15147
rect 12756 15045 12790 15079
rect 16948 15045 16982 15079
rect 19809 15045 19843 15079
rect 21833 15045 21867 15079
rect 25237 15045 25271 15079
rect 29745 15045 29779 15079
rect 3157 14977 3191 15011
rect 3433 14977 3467 15011
rect 4445 14977 4479 15011
rect 4712 14977 4746 15011
rect 6377 14977 6411 15011
rect 7021 14977 7055 15011
rect 7288 14977 7322 15011
rect 13001 14977 13035 15011
rect 14096 14977 14130 15011
rect 15853 14977 15887 15011
rect 15945 14977 15979 15011
rect 16681 14977 16715 15011
rect 18521 14977 18555 15011
rect 19993 14977 20027 15011
rect 20085 14977 20119 15011
rect 21005 14977 21039 15011
rect 21281 14977 21315 15011
rect 22017 14977 22051 15011
rect 22293 14977 22327 15011
rect 23397 14977 23431 15011
rect 25881 14977 25915 15011
rect 27629 14977 27663 15011
rect 2421 14909 2455 14943
rect 2697 14909 2731 14943
rect 8953 14909 8987 14943
rect 10609 14909 10643 14943
rect 10793 14909 10827 14943
rect 13829 14909 13863 14943
rect 20361 14909 20395 14943
rect 24317 14909 24351 14943
rect 28089 14909 28123 14943
rect 11621 14841 11655 14875
rect 18061 14841 18095 14875
rect 22201 14841 22235 14875
rect 23121 14841 23155 14875
rect 24041 14841 24075 14875
rect 24869 14841 24903 14875
rect 29193 14841 29227 14875
rect 5825 14773 5859 14807
rect 6561 14773 6595 14807
rect 8401 14773 8435 14807
rect 15209 14773 15243 14807
rect 16129 14773 16163 14807
rect 18751 14773 18785 14807
rect 20821 14773 20855 14807
rect 22937 14773 22971 14807
rect 23857 14773 23891 14807
rect 24777 14773 24811 14807
rect 28641 14773 28675 14807
rect 1501 14569 1535 14603
rect 1961 14569 1995 14603
rect 13185 14569 13219 14603
rect 19901 14569 19935 14603
rect 22385 14569 22419 14603
rect 24409 14569 24443 14603
rect 25789 14569 25823 14603
rect 26893 14569 26927 14603
rect 27445 14569 27479 14603
rect 28457 14569 28491 14603
rect 29653 14569 29687 14603
rect 3019 14501 3053 14535
rect 6561 14501 6595 14535
rect 12633 14501 12667 14535
rect 15485 14501 15519 14535
rect 17417 14501 17451 14535
rect 20361 14501 20395 14535
rect 20729 14501 20763 14535
rect 22201 14501 22235 14535
rect 23029 14501 23063 14535
rect 1869 14433 1903 14467
rect 4445 14433 4479 14467
rect 4721 14433 4755 14467
rect 7021 14433 7055 14467
rect 18429 14433 18463 14467
rect 21649 14433 21683 14467
rect 25145 14433 25179 14467
rect 1685 14365 1719 14399
rect 3249 14365 3283 14399
rect 5181 14365 5215 14399
rect 5448 14365 5482 14399
rect 8953 14365 8987 14399
rect 10793 14365 10827 14399
rect 11253 14365 11287 14399
rect 11520 14365 11554 14399
rect 14105 14365 14139 14399
rect 16037 14365 16071 14399
rect 18705 14365 18739 14399
rect 19257 14365 19291 14399
rect 19487 14365 19521 14399
rect 19717 14365 19751 14399
rect 20545 14365 20579 14399
rect 20821 14365 20855 14399
rect 21465 14365 21499 14399
rect 21741 14365 21775 14399
rect 23213 14365 23247 14399
rect 23397 14365 23431 14399
rect 24593 14365 24627 14399
rect 25053 14365 25087 14399
rect 25237 14365 25271 14399
rect 1961 14297 1995 14331
rect 7288 14297 7322 14331
rect 10609 14297 10643 14331
rect 13369 14297 13403 14331
rect 13553 14297 13587 14331
rect 14350 14297 14384 14331
rect 16304 14297 16338 14331
rect 21281 14297 21315 14331
rect 22569 14297 22603 14331
rect 30113 14297 30147 14331
rect 8401 14229 8435 14263
rect 22359 14229 22393 14263
rect 26341 14229 26375 14263
rect 27905 14229 27939 14263
rect 30665 14229 30699 14263
rect 2513 14025 2547 14059
rect 5825 14025 5859 14059
rect 7757 14025 7791 14059
rect 22661 14025 22695 14059
rect 23495 14025 23529 14059
rect 23581 14025 23615 14059
rect 28089 14025 28123 14059
rect 28641 14025 28675 14059
rect 29285 14025 29319 14059
rect 30849 14025 30883 14059
rect 8401 13957 8435 13991
rect 11774 13957 11808 13991
rect 13829 13957 13863 13991
rect 16948 13957 16982 13991
rect 21833 13957 21867 13991
rect 22033 13957 22067 13991
rect 22937 13957 22971 13991
rect 25329 13957 25363 13991
rect 25881 13957 25915 13991
rect 27537 13957 27571 13991
rect 1409 13889 1443 13923
rect 2145 13889 2179 13923
rect 2329 13889 2363 13923
rect 2697 13889 2731 13923
rect 4445 13889 4479 13923
rect 4712 13889 4746 13923
rect 6377 13889 6411 13923
rect 6644 13889 6678 13923
rect 8217 13889 8251 13923
rect 10701 13889 10735 13923
rect 10793 13889 10827 13923
rect 10977 13889 11011 13923
rect 14657 13889 14691 13923
rect 14924 13889 14958 13923
rect 16681 13889 16715 13923
rect 18613 13889 18647 13923
rect 18889 13889 18923 13923
rect 19717 13889 19751 13923
rect 20453 13889 20487 13923
rect 20545 13889 20579 13923
rect 20729 13889 20763 13923
rect 22683 13889 22717 13923
rect 23397 13889 23431 13923
rect 23682 13879 23716 13913
rect 24133 13889 24167 13923
rect 24317 13889 24351 13923
rect 24869 13889 24903 13923
rect 30297 13889 30331 13923
rect 3709 13821 3743 13855
rect 3985 13821 4019 13855
rect 10057 13821 10091 13855
rect 11529 13821 11563 13855
rect 13921 13821 13955 13855
rect 14013 13821 14047 13855
rect 18705 13821 18739 13855
rect 18797 13821 18831 13855
rect 19993 13821 20027 13855
rect 26985 13821 27019 13855
rect 29745 13821 29779 13855
rect 1593 13753 1627 13787
rect 10517 13753 10551 13787
rect 12909 13753 12943 13787
rect 16037 13753 16071 13787
rect 18061 13753 18095 13787
rect 19533 13753 19567 13787
rect 19901 13753 19935 13787
rect 22753 13753 22787 13787
rect 2237 13685 2271 13719
rect 10885 13685 10919 13719
rect 13461 13685 13495 13719
rect 19073 13685 19107 13719
rect 20913 13685 20947 13719
rect 22017 13685 22051 13719
rect 22201 13685 22235 13719
rect 24133 13685 24167 13719
rect 1685 13481 1719 13515
rect 4077 13481 4111 13515
rect 4261 13481 4295 13515
rect 6101 13481 6135 13515
rect 19257 13481 19291 13515
rect 22109 13481 22143 13515
rect 22661 13481 22695 13515
rect 23397 13481 23431 13515
rect 25053 13481 25087 13515
rect 26065 13481 26099 13515
rect 27261 13481 27295 13515
rect 28273 13481 28307 13515
rect 30113 13481 30147 13515
rect 13553 13413 13587 13447
rect 18337 13413 18371 13447
rect 26709 13413 26743 13447
rect 28917 13413 28951 13447
rect 1501 13345 1535 13379
rect 2697 13345 2731 13379
rect 2789 13345 2823 13379
rect 3893 13345 3927 13379
rect 6561 13345 6595 13379
rect 19717 13345 19751 13379
rect 21097 13345 21131 13379
rect 25513 13345 25547 13379
rect 1685 13277 1719 13311
rect 2881 13277 2915 13311
rect 3801 13277 3835 13311
rect 4077 13277 4111 13311
rect 4721 13277 4755 13311
rect 10793 13277 10827 13311
rect 11253 13277 11287 13311
rect 13369 13277 13403 13311
rect 14105 13277 14139 13311
rect 15945 13277 15979 13311
rect 17969 13277 18003 13311
rect 19441 13277 19475 13311
rect 19625 13277 19659 13311
rect 20361 13277 20395 13311
rect 20637 13277 20671 13311
rect 21281 13277 21315 13311
rect 22937 13277 22971 13311
rect 23581 13277 23615 13311
rect 24501 13277 24535 13311
rect 1409 13209 1443 13243
rect 4966 13209 5000 13243
rect 6745 13209 6779 13243
rect 8401 13209 8435 13243
rect 8953 13209 8987 13243
rect 10609 13209 10643 13243
rect 11498 13209 11532 13243
rect 13185 13209 13219 13243
rect 14372 13209 14406 13243
rect 16190 13209 16224 13243
rect 18061 13209 18095 13243
rect 21465 13209 21499 13243
rect 22017 13209 22051 13243
rect 22661 13209 22695 13243
rect 22845 13209 22879 13243
rect 27721 13209 27755 13243
rect 1869 13141 1903 13175
rect 3249 13141 3283 13175
rect 12633 13141 12667 13175
rect 15485 13141 15519 13175
rect 17325 13141 17359 13175
rect 17785 13141 17819 13175
rect 18153 13141 18187 13175
rect 20177 13141 20211 13175
rect 20545 13141 20579 13175
rect 29561 13141 29595 13175
rect 30665 13141 30699 13175
rect 1869 12937 1903 12971
rect 3525 12937 3559 12971
rect 7849 12937 7883 12971
rect 15531 12937 15565 12971
rect 16681 12937 16715 12971
rect 19599 12937 19633 12971
rect 23029 12937 23063 12971
rect 25973 12937 26007 12971
rect 28181 12937 28215 12971
rect 28733 12937 28767 12971
rect 29285 12937 29319 12971
rect 3617 12869 3651 12903
rect 8493 12869 8527 12903
rect 14596 12869 14630 12903
rect 18521 12869 18555 12903
rect 19809 12869 19843 12903
rect 20269 12869 20303 12903
rect 20485 12869 20519 12903
rect 21189 12869 21223 12903
rect 22385 12869 22419 12903
rect 25513 12869 25547 12903
rect 1409 12801 1443 12835
rect 1593 12801 1627 12835
rect 1685 12801 1719 12835
rect 2513 12801 2547 12835
rect 2789 12801 2823 12835
rect 4445 12801 4479 12835
rect 4712 12801 4746 12835
rect 6469 12801 6503 12835
rect 6736 12801 6770 12835
rect 8309 12801 8343 12835
rect 10793 12801 10827 12835
rect 12734 12801 12768 12835
rect 13001 12801 13035 12835
rect 14841 12801 14875 12835
rect 15301 12801 15335 12835
rect 17794 12801 17828 12835
rect 18705 12801 18739 12835
rect 18981 12801 19015 12835
rect 21097 12801 21131 12835
rect 21281 12801 21315 12835
rect 22201 12801 22235 12835
rect 23673 12801 23707 12835
rect 23857 12801 23891 12835
rect 24409 12801 24443 12835
rect 2697 12733 2731 12767
rect 3341 12733 3375 12767
rect 8769 12733 8803 12767
rect 10609 12733 10643 12767
rect 18061 12733 18095 12767
rect 24961 12733 24995 12767
rect 29745 12733 29779 12767
rect 2329 12665 2363 12699
rect 11621 12665 11655 12699
rect 23489 12665 23523 12699
rect 27537 12665 27571 12699
rect 1593 12597 1627 12631
rect 2513 12597 2547 12631
rect 3985 12597 4019 12631
rect 5825 12597 5859 12631
rect 10977 12597 11011 12631
rect 13461 12597 13495 12631
rect 18889 12597 18923 12631
rect 19441 12597 19475 12631
rect 19625 12597 19659 12631
rect 20453 12597 20487 12631
rect 20637 12597 20671 12631
rect 27077 12597 27111 12631
rect 2605 12393 2639 12427
rect 15485 12393 15519 12427
rect 17877 12393 17911 12427
rect 21557 12393 21591 12427
rect 25605 12393 25639 12427
rect 26157 12393 26191 12427
rect 28273 12393 28307 12427
rect 1869 12325 1903 12359
rect 16497 12325 16531 12359
rect 17325 12325 17359 12359
rect 20269 12325 20303 12359
rect 21005 12325 21039 12359
rect 27813 12325 27847 12359
rect 2513 12257 2547 12291
rect 4537 12257 4571 12291
rect 4721 12257 4755 12291
rect 8953 12257 8987 12291
rect 9137 12257 9171 12291
rect 10425 12257 10459 12291
rect 11253 12257 11287 12291
rect 12725 12257 12759 12291
rect 18245 12257 18279 12291
rect 19625 12257 19659 12291
rect 29561 12257 29595 12291
rect 2421 12189 2455 12223
rect 2697 12189 2731 12223
rect 5825 12189 5859 12223
rect 6101 12189 6135 12223
rect 8401 12189 8435 12223
rect 14105 12189 14139 12223
rect 16129 12189 16163 12223
rect 16313 12189 16347 12223
rect 17141 12189 17175 12223
rect 17417 12189 17451 12223
rect 18061 12189 18095 12223
rect 18337 12189 18371 12223
rect 19441 12189 19475 12223
rect 20085 12189 20119 12223
rect 20821 12189 20855 12223
rect 21557 12189 21591 12223
rect 21741 12189 21775 12223
rect 22569 12189 22603 12223
rect 23213 12189 23247 12223
rect 23397 12189 23431 12223
rect 28825 12189 28859 12223
rect 1501 12121 1535 12155
rect 6561 12121 6595 12155
rect 8217 12121 8251 12155
rect 11437 12121 11471 12155
rect 14372 12121 14406 12155
rect 16957 12121 16991 12155
rect 19257 12121 19291 12155
rect 24409 12121 24443 12155
rect 25053 12121 25087 12155
rect 30113 12121 30147 12155
rect 1961 12053 1995 12087
rect 2881 12053 2915 12087
rect 4077 12053 4111 12087
rect 4445 12053 4479 12087
rect 15945 12053 15979 12087
rect 16221 12053 16255 12087
rect 22753 12053 22787 12087
rect 23305 12053 23339 12087
rect 26617 12053 26651 12087
rect 27261 12053 27295 12087
rect 3709 11849 3743 11883
rect 5365 11849 5399 11883
rect 13369 11849 13403 11883
rect 15761 11849 15795 11883
rect 18521 11849 18555 11883
rect 20269 11849 20303 11883
rect 21833 11849 21867 11883
rect 22661 11849 22695 11883
rect 27537 11849 27571 11883
rect 28089 11849 28123 11883
rect 28641 11849 28675 11883
rect 1685 11781 1719 11815
rect 10333 11781 10367 11815
rect 11796 11781 11830 11815
rect 14504 11781 14538 11815
rect 15485 11781 15519 11815
rect 19501 11781 19535 11815
rect 19717 11781 19751 11815
rect 22017 11781 22051 11815
rect 22845 11781 22879 11815
rect 24041 11781 24075 11815
rect 25697 11781 25731 11815
rect 26341 11781 26375 11815
rect 3249 11713 3283 11747
rect 3433 11713 3467 11747
rect 3525 11713 3559 11747
rect 4169 11713 4203 11747
rect 4438 11713 4472 11747
rect 5457 11713 5491 11747
rect 7104 11713 7138 11747
rect 10517 11713 10551 11747
rect 15393 11713 15427 11747
rect 15577 11713 15611 11747
rect 16681 11713 16715 11747
rect 16865 11713 16899 11747
rect 17601 11713 17635 11747
rect 18705 11713 18739 11747
rect 18889 11713 18923 11747
rect 20177 11713 20211 11747
rect 20361 11713 20395 11747
rect 21005 11713 21039 11747
rect 21189 11713 21223 11747
rect 22201 11713 22235 11747
rect 23029 11713 23063 11747
rect 29745 11713 29779 11747
rect 2329 11645 2363 11679
rect 2789 11645 2823 11679
rect 4353 11645 4387 11679
rect 5273 11645 5307 11679
rect 6837 11645 6871 11679
rect 9045 11645 9079 11679
rect 11529 11645 11563 11679
rect 14749 11645 14783 11679
rect 15209 11645 15243 11679
rect 17141 11645 17175 11679
rect 29193 11645 29227 11679
rect 1869 11577 1903 11611
rect 2697 11577 2731 11611
rect 8217 11577 8251 11611
rect 12909 11577 12943 11611
rect 17049 11577 17083 11611
rect 17877 11577 17911 11611
rect 19349 11577 19383 11611
rect 20821 11577 20855 11611
rect 3249 11509 3283 11543
rect 4445 11509 4479 11543
rect 4629 11509 4663 11543
rect 5825 11509 5859 11543
rect 18061 11509 18095 11543
rect 19533 11509 19567 11543
rect 23581 11509 23615 11543
rect 24593 11509 24627 11543
rect 25237 11509 25271 11543
rect 26985 11509 27019 11543
rect 1685 11305 1719 11339
rect 4629 11305 4663 11339
rect 12633 11305 12667 11339
rect 13093 11305 13127 11339
rect 13553 11305 13587 11339
rect 17325 11305 17359 11339
rect 20085 11305 20119 11339
rect 21005 11305 21039 11339
rect 22569 11305 22603 11339
rect 23489 11305 23523 11339
rect 24409 11305 24443 11339
rect 27261 11305 27295 11339
rect 3157 11237 3191 11271
rect 5089 11237 5123 11271
rect 15485 11237 15519 11271
rect 27813 11237 27847 11271
rect 28365 11237 28399 11271
rect 29009 11237 29043 11271
rect 3249 11169 3283 11203
rect 5549 11169 5583 11203
rect 5733 11169 5767 11203
rect 6561 11169 6595 11203
rect 7849 11169 7883 11203
rect 9137 11169 9171 11203
rect 9413 11169 9447 11203
rect 13185 11169 13219 11203
rect 15117 11169 15151 11203
rect 16037 11169 16071 11203
rect 18061 11169 18095 11203
rect 21649 11169 21683 11203
rect 25053 11169 25087 11203
rect 26709 11169 26743 11203
rect 1869 11101 1903 11135
rect 4353 11101 4387 11135
rect 4445 11101 4479 11135
rect 5457 11101 5491 11135
rect 6285 11101 6319 11135
rect 7573 11101 7607 11135
rect 8953 11101 8987 11135
rect 11253 11101 11287 11135
rect 13369 11101 13403 11135
rect 14381 11101 14415 11135
rect 14473 11101 14507 11135
rect 15301 11101 15335 11135
rect 15577 11101 15611 11135
rect 16129 11101 16163 11135
rect 16313 11101 16347 11135
rect 18429 11101 18463 11135
rect 19533 11101 19567 11135
rect 22017 11101 22051 11135
rect 23673 11101 23707 11135
rect 2789 11033 2823 11067
rect 4629 11033 4663 11067
rect 11498 11033 11532 11067
rect 13093 11033 13127 11067
rect 14289 11033 14323 11067
rect 14657 11033 14691 11067
rect 16957 11033 16991 11067
rect 17141 11033 17175 11067
rect 18245 11033 18279 11067
rect 19349 11033 19383 11067
rect 20269 11033 20303 11067
rect 20453 11033 20487 11067
rect 21097 11033 21131 11067
rect 21833 11033 21867 11067
rect 22753 11033 22787 11067
rect 22937 11033 22971 11067
rect 23857 11033 23891 11067
rect 24777 11033 24811 11067
rect 25697 11033 25731 11067
rect 26249 11033 26283 11067
rect 4169 10965 4203 10999
rect 14105 10965 14139 10999
rect 16497 10965 16531 10999
rect 24869 10965 24903 10999
rect 2329 10761 2363 10795
rect 3801 10761 3835 10795
rect 5825 10761 5859 10795
rect 9597 10761 9631 10795
rect 14565 10761 14599 10795
rect 14933 10761 14967 10795
rect 19717 10761 19751 10795
rect 20729 10761 20763 10795
rect 22385 10761 22419 10795
rect 23397 10761 23431 10795
rect 25053 10761 25087 10795
rect 27537 10761 27571 10795
rect 28181 10761 28215 10795
rect 4445 10693 4479 10727
rect 6469 10693 6503 10727
rect 13553 10693 13587 10727
rect 18245 10693 18279 10727
rect 19257 10693 19291 10727
rect 25697 10693 25731 10727
rect 1409 10625 1443 10659
rect 1593 10625 1627 10659
rect 2145 10625 2179 10659
rect 3249 10625 3283 10659
rect 3893 10625 3927 10659
rect 5365 10625 5399 10659
rect 5641 10625 5675 10659
rect 6377 10625 6411 10659
rect 8585 10625 8619 10659
rect 10721 10625 10755 10659
rect 11796 10625 11830 10659
rect 13737 10625 13771 10659
rect 14749 10625 14783 10659
rect 15025 10625 15059 10659
rect 15761 10625 15795 10659
rect 18337 10625 18371 10659
rect 26985 10625 27019 10659
rect 5549 10557 5583 10591
rect 7021 10557 7055 10591
rect 8309 10557 8343 10591
rect 10977 10557 11011 10591
rect 11529 10557 11563 10591
rect 13461 10557 13495 10591
rect 15485 10557 15519 10591
rect 17233 10557 17267 10591
rect 17693 10557 17727 10591
rect 20177 10557 20211 10591
rect 24593 10557 24627 10591
rect 1593 10489 1627 10523
rect 4813 10489 4847 10523
rect 12909 10489 12943 10523
rect 14013 10489 14047 10523
rect 17417 10489 17451 10523
rect 18889 10489 18923 10523
rect 19901 10489 19935 10523
rect 3065 10421 3099 10455
rect 4905 10421 4939 10455
rect 5641 10421 5675 10455
rect 7251 10421 7285 10455
rect 15577 10421 15611 10455
rect 15945 10421 15979 10455
rect 16681 10421 16715 10455
rect 18797 10421 18831 10455
rect 21189 10421 21223 10455
rect 21925 10421 21959 10455
rect 24041 10421 24075 10455
rect 26249 10421 26283 10455
rect 1593 10217 1627 10251
rect 1869 10217 1903 10251
rect 5549 10217 5583 10251
rect 6009 10217 6043 10251
rect 8953 10217 8987 10251
rect 9413 10217 9447 10251
rect 14105 10217 14139 10251
rect 14473 10217 14507 10251
rect 17233 10217 17267 10251
rect 18153 10217 18187 10251
rect 22661 10217 22695 10251
rect 23305 10217 23339 10251
rect 25053 10217 25087 10251
rect 26249 10217 26283 10251
rect 43361 10217 43395 10251
rect 2605 10149 2639 10183
rect 4169 10149 4203 10183
rect 4997 10149 5031 10183
rect 7205 10149 7239 10183
rect 9873 10149 9907 10183
rect 13093 10149 13127 10183
rect 15301 10149 15335 10183
rect 15485 10149 15519 10183
rect 17417 10149 17451 10183
rect 19533 10149 19567 10183
rect 19717 10149 19751 10183
rect 25605 10149 25639 10183
rect 26893 10149 26927 10183
rect 1593 10081 1627 10115
rect 5641 10081 5675 10115
rect 6561 10081 6595 10115
rect 7757 10081 7791 10115
rect 7941 10081 7975 10115
rect 9137 10081 9171 10115
rect 16405 10081 16439 10115
rect 1685 10013 1719 10047
rect 2421 10013 2455 10047
rect 3065 10013 3099 10047
rect 3249 10013 3283 10047
rect 5825 10013 5859 10047
rect 6745 10013 6779 10047
rect 8953 10013 8987 10047
rect 9229 10013 9263 10047
rect 11253 10013 11287 10047
rect 11713 10013 11747 10047
rect 14289 10013 14323 10047
rect 14565 10013 14599 10047
rect 15025 10013 15059 10047
rect 17693 10013 17727 10047
rect 19257 10013 19291 10047
rect 21649 10013 21683 10047
rect 24593 10013 24627 10047
rect 27077 10013 27111 10047
rect 28089 10013 28123 10047
rect 29009 10013 29043 10047
rect 29561 10013 29595 10047
rect 43913 10013 43947 10047
rect 1409 9945 1443 9979
rect 3985 9945 4019 9979
rect 4629 9945 4663 9979
rect 5549 9945 5583 9979
rect 6837 9945 6871 9979
rect 11008 9945 11042 9979
rect 11958 9945 11992 9979
rect 16589 9945 16623 9979
rect 16773 9945 16807 9979
rect 18337 9945 18371 9979
rect 18521 9945 18555 9979
rect 20453 9945 20487 9979
rect 20591 9945 20625 9979
rect 20729 9945 20763 9979
rect 21023 9945 21057 9979
rect 3157 9877 3191 9911
rect 5089 9877 5123 9911
rect 8033 9877 8067 9911
rect 8401 9877 8435 9911
rect 22109 9877 22143 9911
rect 23765 9877 23799 9911
rect 24409 9877 24443 9911
rect 27905 9877 27939 9911
rect 28825 9877 28859 9911
rect 44097 9877 44131 9911
rect 7021 9673 7055 9707
rect 8769 9673 8803 9707
rect 19165 9673 19199 9707
rect 27261 9673 27295 9707
rect 28181 9673 28215 9707
rect 7481 9605 7515 9639
rect 13001 9605 13035 9639
rect 14473 9605 14507 9639
rect 15945 9605 15979 9639
rect 16681 9605 16715 9639
rect 17969 9605 18003 9639
rect 21097 9605 21131 9639
rect 22009 9605 22043 9639
rect 24225 9605 24259 9639
rect 24777 9605 24811 9639
rect 25973 9605 26007 9639
rect 1777 9537 1811 9571
rect 2421 9537 2455 9571
rect 3341 9537 3375 9571
rect 4169 9537 4203 9571
rect 4905 9537 4939 9571
rect 5641 9537 5675 9571
rect 6561 9537 6595 9571
rect 6837 9537 6871 9571
rect 7797 9537 7831 9571
rect 9597 9537 9631 9571
rect 13185 9537 13219 9571
rect 14105 9537 14139 9571
rect 15117 9537 15151 9571
rect 15301 9537 15335 9571
rect 15761 9537 15795 9571
rect 16129 9537 16163 9571
rect 16865 9537 16899 9571
rect 20913 9537 20947 9571
rect 22182 9537 22216 9571
rect 23305 9537 23339 9571
rect 6745 9469 6779 9503
rect 7665 9469 7699 9503
rect 8861 9469 8895 9503
rect 9045 9469 9079 9503
rect 9873 9469 9907 9503
rect 11529 9469 11563 9503
rect 11805 9469 11839 9503
rect 12909 9469 12943 9503
rect 14197 9469 14231 9503
rect 14289 9469 14323 9503
rect 18061 9469 18095 9503
rect 18245 9469 18279 9503
rect 18889 9469 18923 9503
rect 19073 9469 19107 9503
rect 19993 9469 20027 9503
rect 2605 9401 2639 9435
rect 3525 9401 3559 9435
rect 3985 9401 4019 9435
rect 5825 9401 5859 9435
rect 7941 9401 7975 9435
rect 14933 9401 14967 9435
rect 17049 9401 17083 9435
rect 17601 9401 17635 9435
rect 20269 9401 20303 9435
rect 26157 9401 26191 9435
rect 1961 9333 1995 9367
rect 5089 9333 5123 9367
rect 6561 9333 6595 9367
rect 7481 9333 7515 9367
rect 8401 9333 8435 9367
rect 10885 9333 10919 9367
rect 13461 9333 13495 9367
rect 19533 9333 19567 9367
rect 20453 9333 20487 9367
rect 21281 9333 21315 9367
rect 21833 9333 21867 9367
rect 22661 9333 22695 9367
rect 24869 9333 24903 9367
rect 1409 9129 1443 9163
rect 2053 9129 2087 9163
rect 2697 9129 2731 9163
rect 4445 9129 4479 9163
rect 5825 9129 5859 9163
rect 7941 9129 7975 9163
rect 8401 9129 8435 9163
rect 9137 9129 9171 9163
rect 11989 9129 12023 9163
rect 13185 9129 13219 9163
rect 14105 9129 14139 9163
rect 14749 9129 14783 9163
rect 16497 9129 16531 9163
rect 19349 9129 19383 9163
rect 19809 9129 19843 9163
rect 24409 9129 24443 9163
rect 25789 9129 25823 9163
rect 26985 9129 27019 9163
rect 4997 9061 5031 9095
rect 7113 9061 7147 9095
rect 9597 9061 9631 9095
rect 15945 9061 15979 9095
rect 16037 9061 16071 9095
rect 19993 9061 20027 9095
rect 21097 9061 21131 9095
rect 21189 9061 21223 9095
rect 23121 9061 23155 9095
rect 8033 8993 8067 9027
rect 9229 8993 9263 9027
rect 10333 8993 10367 9027
rect 12633 8993 12667 9027
rect 17049 8993 17083 9027
rect 18429 8993 18463 9027
rect 22569 8993 22603 9027
rect 1593 8925 1627 8959
rect 2237 8925 2271 8959
rect 2881 8925 2915 8959
rect 4261 8925 4295 8959
rect 5181 8925 5215 8959
rect 5641 8925 5675 8959
rect 6285 8925 6319 8959
rect 6469 8925 6503 8959
rect 6561 8925 6595 8959
rect 8210 8925 8244 8959
rect 9413 8925 9447 8959
rect 10057 8925 10091 8959
rect 14289 8925 14323 8959
rect 14933 8925 14967 8959
rect 21649 8925 21683 8959
rect 22017 8925 22051 8959
rect 7481 8857 7515 8891
rect 7941 8857 7975 8891
rect 9137 8857 9171 8891
rect 11437 8857 11471 8891
rect 11713 8857 11747 8891
rect 12725 8857 12759 8891
rect 12909 8857 12943 8891
rect 15117 8857 15151 8891
rect 15577 8857 15611 8891
rect 16865 8857 16899 8891
rect 18061 8857 18095 8891
rect 18245 8857 18279 8891
rect 20269 8857 20303 8891
rect 20729 8857 20763 8891
rect 21833 8857 21867 8891
rect 23673 8857 23707 8891
rect 27629 8857 27663 8891
rect 6561 8789 6595 8823
rect 7021 8789 7055 8823
rect 11529 8789 11563 8823
rect 16957 8789 16991 8823
rect 23765 8789 23799 8823
rect 25053 8789 25087 8823
rect 27721 8789 27755 8823
rect 1593 8585 1627 8619
rect 2053 8585 2087 8619
rect 2697 8585 2731 8619
rect 3433 8585 3467 8619
rect 4537 8585 4571 8619
rect 5181 8585 5215 8619
rect 7389 8585 7423 8619
rect 8953 8585 8987 8619
rect 9321 8585 9355 8619
rect 10609 8585 10643 8619
rect 11621 8585 11655 8619
rect 15761 8585 15795 8619
rect 19349 8585 19383 8619
rect 25513 8585 25547 8619
rect 6653 8517 6687 8551
rect 6837 8517 6871 8551
rect 7573 8517 7607 8551
rect 12817 8517 12851 8551
rect 13033 8517 13067 8551
rect 13645 8517 13679 8551
rect 13861 8517 13895 8551
rect 14565 8517 14599 8551
rect 14749 8517 14783 8551
rect 19809 8517 19843 8551
rect 22569 8517 22603 8551
rect 1409 8449 1443 8483
rect 2237 8449 2271 8483
rect 2881 8449 2915 8483
rect 4353 8449 4387 8483
rect 4997 8449 5031 8483
rect 5825 8449 5859 8483
rect 7297 8449 7331 8483
rect 10149 8449 10183 8483
rect 10333 8449 10367 8483
rect 10425 8449 10459 8483
rect 11989 8449 12023 8483
rect 16681 8449 16715 8483
rect 17601 8449 17635 8483
rect 18337 8449 18371 8483
rect 18521 8449 18555 8483
rect 18705 8449 18739 8483
rect 23305 8449 23339 8483
rect 24409 8449 24443 8483
rect 8033 8381 8067 8415
rect 9413 8381 9447 8415
rect 9597 8381 9631 8415
rect 12081 8381 12115 8415
rect 12265 8381 12299 8415
rect 15853 8381 15887 8415
rect 16037 8381 16071 8415
rect 17141 8381 17175 8415
rect 20269 8381 20303 8415
rect 20729 8381 20763 8415
rect 25973 8381 26007 8415
rect 7573 8313 7607 8347
rect 8401 8313 8435 8347
rect 13185 8313 13219 8347
rect 14013 8313 14047 8347
rect 15393 8313 15427 8347
rect 16957 8313 16991 8347
rect 19533 8313 19567 8347
rect 20545 8313 20579 8347
rect 21281 8313 21315 8347
rect 22753 8313 22787 8347
rect 23857 8313 23891 8347
rect 5641 8245 5675 8279
rect 8493 8245 8527 8279
rect 10149 8245 10183 8279
rect 13001 8245 13035 8279
rect 13829 8245 13863 8279
rect 21925 8245 21959 8279
rect 24961 8245 24995 8279
rect 2053 8041 2087 8075
rect 2605 8041 2639 8075
rect 3249 8041 3283 8075
rect 3801 8041 3835 8075
rect 6193 8041 6227 8075
rect 6653 8041 6687 8075
rect 9137 8041 9171 8075
rect 10149 8041 10183 8075
rect 12633 8041 12667 8075
rect 17785 8041 17819 8075
rect 18613 8041 18647 8075
rect 25053 8041 25087 8075
rect 25605 8041 25639 8075
rect 8217 7973 8251 8007
rect 9229 7905 9263 7939
rect 10517 7905 10551 7939
rect 11989 7905 12023 7939
rect 13185 7905 13219 7939
rect 22385 7905 22419 7939
rect 6009 7837 6043 7871
rect 6837 7837 6871 7871
rect 7297 7837 7331 7871
rect 9413 7837 9447 7871
rect 10333 7837 10367 7871
rect 10609 7837 10643 7871
rect 13093 7837 13127 7871
rect 14289 7837 14323 7871
rect 15025 7837 15059 7871
rect 15669 7837 15703 7871
rect 16313 7837 16347 7871
rect 16957 7837 16991 7871
rect 17141 7837 17175 7871
rect 17969 7837 18003 7871
rect 19809 7837 19843 7871
rect 20085 7837 20119 7871
rect 21005 7837 21039 7871
rect 21465 7837 21499 7871
rect 22661 7837 22695 7871
rect 1593 7769 1627 7803
rect 4905 7769 4939 7803
rect 7941 7769 7975 7803
rect 9137 7769 9171 7803
rect 11897 7769 11931 7803
rect 14105 7769 14139 7803
rect 17325 7769 17359 7803
rect 18153 7769 18187 7803
rect 4353 7701 4387 7735
rect 5549 7701 5583 7735
rect 7481 7701 7515 7735
rect 8401 7701 8435 7735
rect 9597 7701 9631 7735
rect 11437 7701 11471 7735
rect 11805 7701 11839 7735
rect 13001 7701 13035 7735
rect 14841 7701 14875 7735
rect 15485 7701 15519 7735
rect 16129 7701 16163 7735
rect 20821 7701 20855 7735
rect 21649 7701 21683 7735
rect 23765 7701 23799 7735
rect 24409 7701 24443 7735
rect 1593 7497 1627 7531
rect 2145 7497 2179 7531
rect 4077 7497 4111 7531
rect 4997 7497 5031 7531
rect 6469 7497 6503 7531
rect 8125 7497 8159 7531
rect 8861 7497 8895 7531
rect 9321 7497 9355 7531
rect 14473 7497 14507 7531
rect 2697 7429 2731 7463
rect 3249 7429 3283 7463
rect 5825 7429 5859 7463
rect 8585 7429 8619 7463
rect 10425 7429 10459 7463
rect 12817 7429 12851 7463
rect 13001 7429 13035 7463
rect 14841 7429 14875 7463
rect 17049 7429 17083 7463
rect 17233 7429 17267 7463
rect 1409 7361 1443 7395
rect 6929 7361 6963 7395
rect 7941 7361 7975 7395
rect 8769 7361 8803 7395
rect 8861 7361 8895 7395
rect 9781 7361 9815 7395
rect 10609 7361 10643 7395
rect 11897 7361 11931 7395
rect 13645 7361 13679 7395
rect 15853 7361 15887 7395
rect 18889 7361 18923 7395
rect 19349 7361 19383 7395
rect 20821 7361 20855 7395
rect 22109 7361 22143 7395
rect 23397 7361 23431 7395
rect 10333 7293 10367 7327
rect 11989 7293 12023 7327
rect 12173 7293 12207 7327
rect 14933 7293 14967 7327
rect 15117 7293 15151 7327
rect 16957 7293 16991 7327
rect 18613 7293 18647 7327
rect 19625 7293 19659 7327
rect 22385 7293 22419 7327
rect 23673 7293 23707 7327
rect 9505 7225 9539 7259
rect 10885 7225 10919 7259
rect 7113 7157 7147 7191
rect 11529 7157 11563 7191
rect 13461 7157 13495 7191
rect 15669 7157 15703 7191
rect 17509 7157 17543 7191
rect 20637 7157 20671 7191
rect 24777 7157 24811 7191
rect 8401 6953 8435 6987
rect 10701 6953 10735 6987
rect 12633 6953 12667 6987
rect 14105 6953 14139 6987
rect 9321 6885 9355 6919
rect 19901 6885 19935 6919
rect 4445 6817 4479 6851
rect 5181 6817 5215 6851
rect 5733 6817 5767 6851
rect 6837 6817 6871 6851
rect 9597 6817 9631 6851
rect 11989 6817 12023 6851
rect 14749 6817 14783 6851
rect 15301 6817 15335 6851
rect 22201 6817 22235 6851
rect 43729 6817 43763 6851
rect 1409 6749 1443 6783
rect 6285 6749 6319 6783
rect 7297 6749 7331 6783
rect 8217 6749 8251 6783
rect 13461 6749 13495 6783
rect 17417 6749 17451 6783
rect 18429 6749 18463 6783
rect 18705 6749 18739 6783
rect 20637 6749 20671 6783
rect 21557 6749 21591 6783
rect 22477 6749 22511 6783
rect 23673 6749 23707 6783
rect 24593 6749 24627 6783
rect 2605 6681 2639 6715
rect 3801 6681 3835 6715
rect 10685 6681 10719 6715
rect 10885 6681 10919 6715
rect 11805 6681 11839 6715
rect 12725 6681 12759 6715
rect 19349 6681 19383 6715
rect 19625 6681 19659 6715
rect 1593 6613 1627 6647
rect 3065 6613 3099 6647
rect 7481 6613 7515 6647
rect 9137 6613 9171 6647
rect 10517 6613 10551 6647
rect 11345 6613 11379 6647
rect 11713 6613 11747 6647
rect 13277 6613 13311 6647
rect 15761 6613 15795 6647
rect 16681 6613 16715 6647
rect 17233 6613 17267 6647
rect 19441 6613 19475 6647
rect 20453 6613 20487 6647
rect 21741 6613 21775 6647
rect 23489 6613 23523 6647
rect 24409 6613 24443 6647
rect 25145 6613 25179 6647
rect 25605 6613 25639 6647
rect 1869 6409 1903 6443
rect 2789 6409 2823 6443
rect 3893 6409 3927 6443
rect 4353 6409 4387 6443
rect 5825 6409 5859 6443
rect 7205 6409 7239 6443
rect 8309 6409 8343 6443
rect 8953 6409 8987 6443
rect 9597 6409 9631 6443
rect 12265 6409 12299 6443
rect 13001 6409 13035 6443
rect 14841 6409 14875 6443
rect 15945 6409 15979 6443
rect 17325 6409 17359 6443
rect 10517 6341 10551 6375
rect 11805 6341 11839 6375
rect 18153 6341 18187 6375
rect 19717 6341 19751 6375
rect 21925 6341 21959 6375
rect 23581 6341 23615 6375
rect 1409 6273 1443 6307
rect 1593 6273 1627 6307
rect 1685 6273 1719 6307
rect 3249 6273 3283 6307
rect 6745 6273 6779 6307
rect 7849 6273 7883 6307
rect 8493 6273 8527 6307
rect 9137 6273 9171 6307
rect 9781 6273 9815 6307
rect 10333 6273 10367 6307
rect 10609 6273 10643 6307
rect 11621 6273 11655 6307
rect 12449 6273 12483 6307
rect 12909 6273 12943 6307
rect 13093 6273 13127 6307
rect 13541 6273 13575 6307
rect 13737 6273 13771 6307
rect 18337 6273 18371 6307
rect 19625 6273 19659 6307
rect 13645 6205 13679 6239
rect 15393 6205 15427 6239
rect 18061 6205 18095 6239
rect 19809 6205 19843 6239
rect 20821 6205 20855 6239
rect 5273 6137 5307 6171
rect 14197 6137 14231 6171
rect 16773 6137 16807 6171
rect 18613 6137 18647 6171
rect 20177 6137 20211 6171
rect 24133 6137 24167 6171
rect 1593 6069 1627 6103
rect 10333 6069 10367 6103
rect 22385 6069 22419 6103
rect 22937 6069 22971 6103
rect 24593 6069 24627 6103
rect 25237 6069 25271 6103
rect 25697 6069 25731 6103
rect 26249 6069 26283 6103
rect 43085 6069 43119 6103
rect 43637 6069 43671 6103
rect 44189 6069 44223 6103
rect 1409 5865 1443 5899
rect 2697 5865 2731 5899
rect 3801 5865 3835 5899
rect 6653 5865 6687 5899
rect 7849 5865 7883 5899
rect 8401 5865 8435 5899
rect 9229 5865 9263 5899
rect 10609 5865 10643 5899
rect 11253 5865 11287 5899
rect 12265 5865 12299 5899
rect 13553 5865 13587 5899
rect 14841 5865 14875 5899
rect 16405 5865 16439 5899
rect 16957 5865 16991 5899
rect 18153 5865 18187 5899
rect 18705 5865 18739 5899
rect 19349 5865 19383 5899
rect 19901 5865 19935 5899
rect 21005 5865 21039 5899
rect 23121 5865 23155 5899
rect 26617 5865 26651 5899
rect 27169 5865 27203 5899
rect 27813 5865 27847 5899
rect 2145 5797 2179 5831
rect 3157 5797 3191 5831
rect 26065 5797 26099 5831
rect 13001 5729 13035 5763
rect 14197 5729 14231 5763
rect 20361 5729 20395 5763
rect 24961 5729 24995 5763
rect 1593 5661 1627 5695
rect 9873 5661 9907 5695
rect 10425 5661 10459 5695
rect 10609 5661 10643 5695
rect 11069 5661 11103 5695
rect 11253 5661 11287 5695
rect 14473 5661 14507 5695
rect 17601 5661 17635 5695
rect 43913 5661 43947 5695
rect 4905 5593 4939 5627
rect 7297 5593 7331 5627
rect 14381 5593 14415 5627
rect 15853 5593 15887 5627
rect 16129 5593 16163 5627
rect 22569 5593 22603 5627
rect 24409 5593 24443 5627
rect 5457 5525 5491 5559
rect 5917 5525 5951 5559
rect 9689 5525 9723 5559
rect 11805 5525 11839 5559
rect 13093 5525 13127 5559
rect 13185 5525 13219 5559
rect 15945 5525 15979 5559
rect 21557 5525 21591 5559
rect 22109 5525 22143 5559
rect 23673 5525 23707 5559
rect 25513 5525 25547 5559
rect 41705 5525 41739 5559
rect 42257 5525 42291 5559
rect 42901 5525 42935 5559
rect 43453 5525 43487 5559
rect 44097 5525 44131 5559
rect 1593 5321 1627 5355
rect 2145 5321 2179 5355
rect 4169 5321 4203 5355
rect 6377 5321 6411 5355
rect 8033 5321 8067 5355
rect 9781 5321 9815 5355
rect 10333 5321 10367 5355
rect 11529 5321 11563 5355
rect 15577 5321 15611 5355
rect 16129 5321 16163 5355
rect 16773 5321 16807 5355
rect 17877 5321 17911 5355
rect 18889 5321 18923 5355
rect 28089 5321 28123 5355
rect 41429 5321 41463 5355
rect 2789 5253 2823 5287
rect 8585 5253 8619 5287
rect 14473 5253 14507 5287
rect 18337 5253 18371 5287
rect 19533 5253 19567 5287
rect 43913 5253 43947 5287
rect 1409 5185 1443 5219
rect 9597 5185 9631 5219
rect 12449 5185 12483 5219
rect 14657 5185 14691 5219
rect 21833 5185 21867 5219
rect 24593 5185 24627 5219
rect 44097 5185 44131 5219
rect 10793 5117 10827 5151
rect 14381 5117 14415 5151
rect 20545 5117 20579 5151
rect 23489 5117 23523 5151
rect 27537 5117 27571 5151
rect 3433 5049 3467 5083
rect 21097 5049 21131 5083
rect 22937 5049 22971 5083
rect 4721 4981 4755 5015
rect 5273 4981 5307 5015
rect 5825 4981 5859 5015
rect 7389 4981 7423 5015
rect 9045 4981 9079 5015
rect 13001 4981 13035 5015
rect 13553 4981 13587 5015
rect 14933 4981 14967 5015
rect 17233 4981 17267 5015
rect 19993 4981 20027 5015
rect 22385 4981 22419 5015
rect 24041 4981 24075 5015
rect 25145 4981 25179 5015
rect 25697 4981 25731 5015
rect 26341 4981 26375 5015
rect 26985 4981 27019 5015
rect 42625 4981 42659 5015
rect 43453 4981 43487 5015
rect 2697 4777 2731 4811
rect 4629 4777 4663 4811
rect 5181 4777 5215 4811
rect 9137 4777 9171 4811
rect 9689 4777 9723 4811
rect 10517 4777 10551 4811
rect 11253 4777 11287 4811
rect 13185 4777 13219 4811
rect 14749 4777 14783 4811
rect 15209 4777 15243 4811
rect 16681 4777 16715 4811
rect 17785 4777 17819 4811
rect 18337 4777 18371 4811
rect 19349 4777 19383 4811
rect 23673 4777 23707 4811
rect 28825 4777 28859 4811
rect 35909 4777 35943 4811
rect 37933 4777 37967 4811
rect 40785 4777 40819 4811
rect 1593 4709 1627 4743
rect 2237 4709 2271 4743
rect 12725 4709 12759 4743
rect 22109 4709 22143 4743
rect 28273 4709 28307 4743
rect 43913 4709 43947 4743
rect 3893 4641 3927 4675
rect 7297 4641 7331 4675
rect 8401 4641 8435 4675
rect 24409 4641 24443 4675
rect 1409 4573 1443 4607
rect 2053 4573 2087 4607
rect 6837 4573 6871 4607
rect 11713 4573 11747 4607
rect 16129 4573 16163 4607
rect 19809 4573 19843 4607
rect 39129 4573 39163 4607
rect 43177 4573 43211 4607
rect 5733 4505 5767 4539
rect 17233 4505 17267 4539
rect 20913 4505 20947 4539
rect 22569 4505 22603 4539
rect 42165 4505 42199 4539
rect 44097 4505 44131 4539
rect 6285 4437 6319 4471
rect 14197 4437 14231 4471
rect 20361 4437 20395 4471
rect 21465 4437 21499 4471
rect 23121 4437 23155 4471
rect 24961 4437 24995 4471
rect 25513 4437 25547 4471
rect 26157 4437 26191 4471
rect 26617 4437 26651 4471
rect 27261 4437 27295 4471
rect 27721 4437 27755 4471
rect 33793 4437 33827 4471
rect 34805 4437 34839 4471
rect 35357 4437 35391 4471
rect 36553 4437 36587 4471
rect 37289 4437 37323 4471
rect 38669 4437 38703 4471
rect 39865 4437 39899 4471
rect 41429 4437 41463 4471
rect 42717 4437 42751 4471
rect 43361 4437 43395 4471
rect 5825 4233 5859 4267
rect 9505 4233 9539 4267
rect 3985 4165 4019 4199
rect 10057 4165 10091 4199
rect 10701 4165 10735 4199
rect 11621 4165 11655 4199
rect 12633 4165 12667 4199
rect 14381 4165 14415 4199
rect 43361 4165 43395 4199
rect 44097 4165 44131 4199
rect 7757 4097 7791 4131
rect 8401 4097 8435 4131
rect 13185 4097 13219 4131
rect 13829 4097 13863 4131
rect 16681 4097 16715 4131
rect 17417 4097 17451 4131
rect 18429 4097 18463 4131
rect 19533 4097 19567 4131
rect 19993 4097 20027 4131
rect 26249 4097 26283 4131
rect 27537 4097 27571 4131
rect 42441 4097 42475 4131
rect 43177 4097 43211 4131
rect 43913 4097 43947 4131
rect 7297 4029 7331 4063
rect 15393 4029 15427 4063
rect 21833 4029 21867 4063
rect 33609 4029 33643 4063
rect 37841 4029 37875 4063
rect 2053 3961 2087 3995
rect 4721 3961 4755 3995
rect 8585 3961 8619 3995
rect 12173 3961 12207 3995
rect 19349 3961 19383 3995
rect 22385 3961 22419 3995
rect 23581 3961 23615 3995
rect 41889 3961 41923 3995
rect 1409 3893 1443 3927
rect 2697 3893 2731 3927
rect 3341 3893 3375 3927
rect 5181 3893 5215 3927
rect 6745 3893 6779 3927
rect 7941 3893 7975 3927
rect 14841 3893 14875 3927
rect 15945 3893 15979 3927
rect 18613 3893 18647 3927
rect 20545 3893 20579 3927
rect 21097 3893 21131 3927
rect 22937 3893 22971 3927
rect 24041 3893 24075 3927
rect 24593 3893 24627 3927
rect 25145 3893 25179 3927
rect 25697 3893 25731 3927
rect 27353 3893 27387 3927
rect 27997 3893 28031 3927
rect 28733 3893 28767 3927
rect 29377 3893 29411 3927
rect 30021 3893 30055 3927
rect 30757 3893 30791 3927
rect 31217 3893 31251 3927
rect 32321 3893 32355 3927
rect 33149 3893 33183 3927
rect 34621 3893 34655 3927
rect 35357 3893 35391 3927
rect 36093 3893 36127 3927
rect 36553 3893 36587 3927
rect 37289 3893 37323 3927
rect 38853 3893 38887 3927
rect 39773 3893 39807 3927
rect 40233 3893 40267 3927
rect 40785 3893 40819 3927
rect 42625 3893 42659 3927
rect 6653 3689 6687 3723
rect 9505 3689 9539 3723
rect 9965 3689 9999 3723
rect 10793 3689 10827 3723
rect 11437 3689 11471 3723
rect 11897 3689 11931 3723
rect 13369 3689 13403 3723
rect 14105 3689 14139 3723
rect 16589 3689 16623 3723
rect 18337 3689 18371 3723
rect 19441 3689 19475 3723
rect 20545 3689 20579 3723
rect 21281 3689 21315 3723
rect 37473 3689 37507 3723
rect 2697 3621 2731 3655
rect 3985 3621 4019 3655
rect 6009 3621 6043 3655
rect 12725 3621 12759 3655
rect 14749 3621 14783 3655
rect 15577 3621 15611 3655
rect 25053 3621 25087 3655
rect 27261 3621 27295 3655
rect 28181 3621 28215 3655
rect 43177 3621 43211 3655
rect 43913 3621 43947 3655
rect 1961 3553 1995 3587
rect 7665 3553 7699 3587
rect 2237 3485 2271 3519
rect 3801 3485 3835 3519
rect 4445 3485 4479 3519
rect 5825 3485 5859 3519
rect 6469 3485 6503 3519
rect 7941 3485 7975 3519
rect 9321 3485 9355 3519
rect 10609 3485 10643 3519
rect 11253 3485 11287 3519
rect 12081 3485 12115 3519
rect 12909 3485 12943 3519
rect 14289 3485 14323 3519
rect 15761 3485 15795 3519
rect 16773 3485 16807 3519
rect 18153 3485 18187 3519
rect 19257 3485 19291 3519
rect 20361 3485 20395 3519
rect 21465 3485 21499 3519
rect 22385 3485 22419 3519
rect 23397 3485 23431 3519
rect 24593 3485 24627 3519
rect 25237 3485 25271 3519
rect 26525 3485 26559 3519
rect 27997 3485 28031 3519
rect 28917 3485 28951 3519
rect 29561 3485 29595 3519
rect 30297 3485 30331 3519
rect 31033 3485 31067 3519
rect 31953 3485 31987 3519
rect 32965 3485 32999 3519
rect 33885 3485 33919 3519
rect 34805 3485 34839 3519
rect 35725 3485 35759 3519
rect 36645 3485 36679 3519
rect 38117 3485 38151 3519
rect 39129 3485 39163 3519
rect 39865 3485 39899 3519
rect 41613 3485 41647 3519
rect 42349 3485 42383 3519
rect 5365 3417 5399 3451
rect 27077 3417 27111 3451
rect 37565 3417 37599 3451
rect 43361 3417 43395 3451
rect 44097 3417 44131 3451
rect 4629 3349 4663 3383
rect 17233 3349 17267 3383
rect 22201 3349 22235 3383
rect 23213 3349 23247 3383
rect 24409 3349 24443 3383
rect 25697 3349 25731 3383
rect 26341 3349 26375 3383
rect 28733 3349 28767 3383
rect 29745 3349 29779 3383
rect 30481 3349 30515 3383
rect 31217 3349 31251 3383
rect 32137 3349 32171 3383
rect 33149 3349 33183 3383
rect 34069 3349 34103 3383
rect 34989 3349 35023 3383
rect 35909 3349 35943 3383
rect 36829 3349 36863 3383
rect 38301 3349 38335 3383
rect 38945 3349 38979 3383
rect 40049 3349 40083 3383
rect 40693 3349 40727 3383
rect 41797 3349 41831 3383
rect 42533 3349 42567 3383
rect 4169 3145 4203 3179
rect 14381 3145 14415 3179
rect 15025 3145 15059 3179
rect 17785 3145 17819 3179
rect 18245 3145 18279 3179
rect 20177 3145 20211 3179
rect 21005 3145 21039 3179
rect 21925 3145 21959 3179
rect 22845 3145 22879 3179
rect 23765 3145 23799 3179
rect 24593 3145 24627 3179
rect 27077 3145 27111 3179
rect 32597 3145 32631 3179
rect 34069 3145 34103 3179
rect 35541 3145 35575 3179
rect 37381 3145 37415 3179
rect 44005 3145 44039 3179
rect 26065 3077 26099 3111
rect 26249 3077 26283 3111
rect 27629 3077 27663 3111
rect 27813 3077 27847 3111
rect 30297 3077 30331 3111
rect 31033 3077 31067 3111
rect 33425 3077 33459 3111
rect 34713 3077 34747 3111
rect 37473 3077 37507 3111
rect 38025 3077 38059 3111
rect 39497 3077 39531 3111
rect 40233 3077 40267 3111
rect 42809 3077 42843 3111
rect 44097 3077 44131 3111
rect 1961 3009 1995 3043
rect 3249 3009 3283 3043
rect 3985 3009 4019 3043
rect 4629 3009 4663 3043
rect 5549 3009 5583 3043
rect 7573 3009 7607 3043
rect 8585 3009 8619 3043
rect 9321 3009 9355 3043
rect 10517 3009 10551 3043
rect 10793 3009 10827 3043
rect 11805 3009 11839 3043
rect 12265 3009 12299 3043
rect 12909 3009 12943 3043
rect 13553 3009 13587 3043
rect 14565 3009 14599 3043
rect 15209 3009 15243 3043
rect 15945 3009 15979 3043
rect 17141 3009 17175 3043
rect 17601 3009 17635 3043
rect 19073 3009 19107 3043
rect 19993 3009 20027 3043
rect 21189 3009 21223 3043
rect 22109 3009 22143 3043
rect 23029 3009 23063 3043
rect 23949 3009 23983 3043
rect 24777 3009 24811 3043
rect 25513 3009 25547 3043
rect 28825 3009 28859 3043
rect 30113 3009 30147 3043
rect 30849 3009 30883 3043
rect 32689 3009 32723 3043
rect 34161 3009 34195 3043
rect 34897 3009 34931 3043
rect 35633 3009 35667 3043
rect 36553 3009 36587 3043
rect 38209 3009 38243 3043
rect 38945 3009 38979 3043
rect 39681 3009 39715 3043
rect 40417 3009 40451 3043
rect 40969 3009 41003 3043
rect 42993 3009 43027 3043
rect 2237 2941 2271 2975
rect 3525 2941 3559 2975
rect 7297 2941 7331 2975
rect 8861 2941 8895 2975
rect 36369 2941 36403 2975
rect 5733 2873 5767 2907
rect 13093 2873 13127 2907
rect 16129 2873 16163 2907
rect 33241 2873 33275 2907
rect 38761 2873 38795 2907
rect 4813 2805 4847 2839
rect 9505 2805 9539 2839
rect 11621 2805 11655 2839
rect 12449 2805 12483 2839
rect 13737 2805 13771 2839
rect 16957 2805 16991 2839
rect 18889 2805 18923 2839
rect 25329 2805 25363 2839
rect 28365 2805 28399 2839
rect 29055 2805 29089 2839
rect 41153 2805 41187 2839
rect 41797 2805 41831 2839
rect 4261 2601 4295 2635
rect 9137 2601 9171 2635
rect 32597 2601 32631 2635
rect 38025 2601 38059 2635
rect 2697 2533 2731 2567
rect 5733 2533 5767 2567
rect 8401 2533 8435 2567
rect 17785 2533 17819 2567
rect 28411 2533 28445 2567
rect 29791 2533 29825 2567
rect 34713 2533 34747 2567
rect 36185 2533 36219 2567
rect 38945 2533 38979 2567
rect 1961 2465 1995 2499
rect 7297 2465 7331 2499
rect 10149 2465 10183 2499
rect 10425 2465 10459 2499
rect 25973 2465 26007 2499
rect 30849 2465 30883 2499
rect 43545 2465 43579 2499
rect 2237 2397 2271 2431
rect 4905 2397 4939 2431
rect 5549 2397 5583 2431
rect 7021 2397 7055 2431
rect 8217 2397 8251 2431
rect 8953 2397 8987 2431
rect 11805 2397 11839 2431
rect 12541 2397 12575 2431
rect 13369 2397 13403 2431
rect 14381 2397 14415 2431
rect 15209 2397 15243 2431
rect 15669 2397 15703 2431
rect 16957 2397 16991 2431
rect 18521 2397 18555 2431
rect 19993 2397 20027 2431
rect 20913 2397 20947 2431
rect 21833 2397 21867 2431
rect 22845 2397 22879 2431
rect 23765 2397 23799 2431
rect 24409 2397 24443 2431
rect 25789 2397 25823 2431
rect 28181 2397 28215 2431
rect 29561 2397 29595 2431
rect 33241 2397 33275 2431
rect 33425 2397 33459 2431
rect 36369 2397 36403 2431
rect 39865 2397 39899 2431
rect 42993 2397 43027 2431
rect 2881 2329 2915 2363
rect 4353 2329 4387 2363
rect 10885 2329 10919 2363
rect 17601 2329 17635 2363
rect 27445 2329 27479 2363
rect 27629 2329 27663 2363
rect 31033 2329 31067 2363
rect 32689 2329 32723 2363
rect 34897 2329 34931 2363
rect 35633 2329 35667 2363
rect 37473 2329 37507 2363
rect 38117 2329 38151 2363
rect 39129 2329 39163 2363
rect 40969 2329 41003 2363
rect 41705 2329 41739 2363
rect 43729 2329 43763 2363
rect 11621 2261 11655 2295
rect 12357 2261 12391 2295
rect 13185 2261 13219 2295
rect 14197 2261 14231 2295
rect 15025 2261 15059 2295
rect 15853 2261 15887 2295
rect 16773 2261 16807 2295
rect 18337 2261 18371 2295
rect 19809 2261 19843 2295
rect 20729 2261 20763 2295
rect 22017 2261 22051 2295
rect 22661 2261 22695 2295
rect 23581 2261 23615 2295
rect 24593 2261 24627 2295
rect 25145 2261 25179 2295
rect 33977 2261 34011 2295
rect 35541 2261 35575 2295
rect 40049 2261 40083 2295
rect 40877 2261 40911 2295
rect 41613 2261 41647 2295
rect 42901 2261 42935 2295
<< metal1 >>
rect 21818 38020 21824 38072
rect 21876 38060 21882 38072
rect 30006 38060 30012 38072
rect 21876 38032 30012 38060
rect 21876 38020 21882 38032
rect 30006 38020 30012 38032
rect 30064 38020 30070 38072
rect 12710 37952 12716 38004
rect 12768 37992 12774 38004
rect 24946 37992 24952 38004
rect 12768 37964 24952 37992
rect 12768 37952 12774 37964
rect 24946 37952 24952 37964
rect 25004 37952 25010 38004
rect 9490 37884 9496 37936
rect 9548 37924 9554 37936
rect 20254 37924 20260 37936
rect 9548 37896 20260 37924
rect 9548 37884 9554 37896
rect 20254 37884 20260 37896
rect 20312 37884 20318 37936
rect 20898 37884 20904 37936
rect 20956 37924 20962 37936
rect 28166 37924 28172 37936
rect 20956 37896 28172 37924
rect 20956 37884 20962 37896
rect 28166 37884 28172 37896
rect 28224 37884 28230 37936
rect 2774 37816 2780 37868
rect 2832 37856 2838 37868
rect 11146 37856 11152 37868
rect 2832 37828 11152 37856
rect 2832 37816 2838 37828
rect 11146 37816 11152 37828
rect 11204 37816 11210 37868
rect 18046 37816 18052 37868
rect 18104 37856 18110 37868
rect 27430 37856 27436 37868
rect 18104 37828 27436 37856
rect 18104 37816 18110 37828
rect 27430 37816 27436 37828
rect 27488 37816 27494 37868
rect 27706 37816 27712 37868
rect 27764 37856 27770 37868
rect 35802 37856 35808 37868
rect 27764 37828 35808 37856
rect 27764 37816 27770 37828
rect 35802 37816 35808 37828
rect 35860 37816 35866 37868
rect 3050 37748 3056 37800
rect 3108 37788 3114 37800
rect 10318 37788 10324 37800
rect 3108 37760 10324 37788
rect 3108 37748 3114 37760
rect 10318 37748 10324 37760
rect 10376 37748 10382 37800
rect 10410 37748 10416 37800
rect 10468 37788 10474 37800
rect 23842 37788 23848 37800
rect 10468 37760 23848 37788
rect 10468 37748 10474 37760
rect 23842 37748 23848 37760
rect 23900 37748 23906 37800
rect 29822 37748 29828 37800
rect 29880 37788 29886 37800
rect 37826 37788 37832 37800
rect 29880 37760 37832 37788
rect 29880 37748 29886 37760
rect 37826 37748 37832 37760
rect 37884 37748 37890 37800
rect 3970 37680 3976 37732
rect 4028 37720 4034 37732
rect 12434 37720 12440 37732
rect 4028 37692 12440 37720
rect 4028 37680 4034 37692
rect 12434 37680 12440 37692
rect 12492 37680 12498 37732
rect 17770 37680 17776 37732
rect 17828 37720 17834 37732
rect 22554 37720 22560 37732
rect 17828 37692 22560 37720
rect 17828 37680 17834 37692
rect 22554 37680 22560 37692
rect 22612 37680 22618 37732
rect 25314 37680 25320 37732
rect 25372 37720 25378 37732
rect 33318 37720 33324 37732
rect 25372 37692 33324 37720
rect 25372 37680 25378 37692
rect 33318 37680 33324 37692
rect 33376 37680 33382 37732
rect 7650 37612 7656 37664
rect 7708 37652 7714 37664
rect 21450 37652 21456 37664
rect 7708 37624 21456 37652
rect 7708 37612 7714 37624
rect 21450 37612 21456 37624
rect 21508 37612 21514 37664
rect 24302 37612 24308 37664
rect 24360 37652 24366 37664
rect 34698 37652 34704 37664
rect 24360 37624 34704 37652
rect 24360 37612 24366 37624
rect 34698 37612 34704 37624
rect 34756 37612 34762 37664
rect 1104 37562 44896 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 44896 37562
rect 1104 37488 44896 37510
rect 2317 37451 2375 37457
rect 2317 37417 2329 37451
rect 2363 37448 2375 37451
rect 2774 37448 2780 37460
rect 2363 37420 2780 37448
rect 2363 37417 2375 37420
rect 2317 37411 2375 37417
rect 2774 37408 2780 37420
rect 2832 37408 2838 37460
rect 3050 37448 3056 37460
rect 3011 37420 3056 37448
rect 3050 37408 3056 37420
rect 3108 37408 3114 37460
rect 3510 37408 3516 37460
rect 3568 37448 3574 37460
rect 5166 37448 5172 37460
rect 3568 37420 5172 37448
rect 3568 37408 3574 37420
rect 5166 37408 5172 37420
rect 5224 37408 5230 37460
rect 7650 37448 7656 37460
rect 7611 37420 7656 37448
rect 7650 37408 7656 37420
rect 7708 37408 7714 37460
rect 9490 37448 9496 37460
rect 9451 37420 9496 37448
rect 9490 37408 9496 37420
rect 9548 37408 9554 37460
rect 10229 37451 10287 37457
rect 10229 37417 10241 37451
rect 10275 37448 10287 37451
rect 10410 37448 10416 37460
rect 10275 37420 10416 37448
rect 10275 37417 10287 37420
rect 10229 37411 10287 37417
rect 10410 37408 10416 37420
rect 10468 37408 10474 37460
rect 11701 37451 11759 37457
rect 11701 37417 11713 37451
rect 11747 37448 11759 37451
rect 22373 37451 22431 37457
rect 11747 37420 21220 37448
rect 11747 37417 11759 37420
rect 11701 37411 11759 37417
rect 4433 37383 4491 37389
rect 4433 37349 4445 37383
rect 4479 37380 4491 37383
rect 4706 37380 4712 37392
rect 4479 37352 4712 37380
rect 4479 37349 4491 37352
rect 4433 37343 4491 37349
rect 4706 37340 4712 37352
rect 4764 37340 4770 37392
rect 5350 37380 5356 37392
rect 5311 37352 5356 37380
rect 5350 37340 5356 37352
rect 5408 37340 5414 37392
rect 7009 37383 7067 37389
rect 7009 37349 7021 37383
rect 7055 37380 7067 37383
rect 8110 37380 8116 37392
rect 7055 37352 8116 37380
rect 7055 37349 7067 37352
rect 7009 37343 7067 37349
rect 8110 37340 8116 37352
rect 8168 37340 8174 37392
rect 12621 37383 12679 37389
rect 12621 37349 12633 37383
rect 12667 37380 12679 37383
rect 12710 37380 12716 37392
rect 12667 37352 12716 37380
rect 12667 37349 12679 37352
rect 12621 37343 12679 37349
rect 12710 37340 12716 37352
rect 12768 37340 12774 37392
rect 21082 37380 21088 37392
rect 21043 37352 21088 37380
rect 21082 37340 21088 37352
rect 21140 37340 21146 37392
rect 21192 37380 21220 37420
rect 22373 37417 22385 37451
rect 22419 37448 22431 37451
rect 27430 37448 27436 37460
rect 22419 37420 26234 37448
rect 27391 37420 27436 37448
rect 22419 37417 22431 37420
rect 22373 37411 22431 37417
rect 22462 37380 22468 37392
rect 21192 37352 22468 37380
rect 22462 37340 22468 37352
rect 22520 37340 22526 37392
rect 22554 37340 22560 37392
rect 22612 37380 22618 37392
rect 25685 37383 25743 37389
rect 25685 37380 25697 37383
rect 22612 37352 25697 37380
rect 22612 37340 22618 37352
rect 25685 37349 25697 37352
rect 25731 37349 25743 37383
rect 26206 37380 26234 37420
rect 27430 37408 27436 37420
rect 27488 37408 27494 37460
rect 28166 37448 28172 37460
rect 28127 37420 28172 37448
rect 28166 37408 28172 37420
rect 28224 37408 28230 37460
rect 30006 37448 30012 37460
rect 29967 37420 30012 37448
rect 30006 37408 30012 37420
rect 30064 37408 30070 37460
rect 33318 37448 33324 37460
rect 33279 37420 33324 37448
rect 33318 37408 33324 37420
rect 33376 37408 33382 37460
rect 34698 37408 34704 37460
rect 34756 37448 34762 37460
rect 35161 37451 35219 37457
rect 35161 37448 35173 37451
rect 34756 37420 35173 37448
rect 34756 37408 34762 37420
rect 35161 37417 35173 37420
rect 35207 37417 35219 37451
rect 37826 37448 37832 37460
rect 37787 37420 37832 37448
rect 35161 37411 35219 37417
rect 37826 37408 37832 37420
rect 37884 37408 37890 37460
rect 40402 37448 40408 37460
rect 40363 37420 40408 37448
rect 40402 37408 40408 37420
rect 40460 37408 40466 37460
rect 41230 37448 41236 37460
rect 41191 37420 41236 37448
rect 41230 37408 41236 37420
rect 41288 37408 41294 37460
rect 29730 37380 29736 37392
rect 26206 37352 29736 37380
rect 25685 37343 25743 37349
rect 29730 37340 29736 37352
rect 29788 37340 29794 37392
rect 32493 37383 32551 37389
rect 32493 37380 32505 37383
rect 29840 37352 32505 37380
rect 3694 37272 3700 37324
rect 3752 37312 3758 37324
rect 5074 37312 5080 37324
rect 3752 37284 5080 37312
rect 3752 37272 3758 37284
rect 5074 37272 5080 37284
rect 5132 37272 5138 37324
rect 8297 37315 8355 37321
rect 8297 37312 8309 37315
rect 6840 37284 8309 37312
rect 198 37204 204 37256
rect 256 37244 262 37256
rect 1397 37247 1455 37253
rect 1397 37244 1409 37247
rect 256 37216 1409 37244
rect 256 37204 262 37216
rect 1397 37213 1409 37216
rect 1443 37213 1455 37247
rect 1397 37207 1455 37213
rect 1412 37176 1440 37207
rect 1486 37204 1492 37256
rect 1544 37244 1550 37256
rect 2222 37244 2228 37256
rect 1544 37216 2228 37244
rect 1544 37204 1550 37216
rect 2222 37204 2228 37216
rect 2280 37204 2286 37256
rect 2774 37204 2780 37256
rect 2832 37244 2838 37256
rect 2961 37247 3019 37253
rect 2961 37244 2973 37247
rect 2832 37216 2973 37244
rect 2832 37204 2838 37216
rect 2961 37213 2973 37216
rect 3007 37213 3019 37247
rect 2961 37207 3019 37213
rect 3786 37204 3792 37256
rect 3844 37244 3850 37256
rect 4249 37247 4307 37253
rect 4249 37244 4261 37247
rect 3844 37216 4261 37244
rect 3844 37204 3850 37216
rect 4249 37213 4261 37216
rect 4295 37244 4307 37247
rect 4798 37244 4804 37256
rect 4295 37216 4804 37244
rect 4295 37213 4307 37216
rect 4249 37207 4307 37213
rect 4798 37204 4804 37216
rect 4856 37204 4862 37256
rect 4982 37204 4988 37256
rect 5040 37244 5046 37256
rect 5169 37247 5227 37253
rect 5169 37244 5181 37247
rect 5040 37216 5181 37244
rect 5040 37204 5046 37216
rect 5169 37213 5181 37216
rect 5215 37213 5227 37247
rect 5169 37207 5227 37213
rect 6178 37204 6184 37256
rect 6236 37244 6242 37256
rect 6840 37253 6868 37284
rect 8297 37281 8309 37284
rect 8343 37281 8355 37315
rect 8297 37275 8355 37281
rect 10965 37315 11023 37321
rect 10965 37281 10977 37315
rect 11011 37312 11023 37315
rect 12250 37312 12256 37324
rect 11011 37284 12256 37312
rect 11011 37281 11023 37284
rect 10965 37275 11023 37281
rect 12250 37272 12256 37284
rect 12308 37312 12314 37324
rect 12308 37284 12480 37312
rect 12308 37272 12314 37284
rect 6825 37247 6883 37253
rect 6825 37244 6837 37247
rect 6236 37216 6837 37244
rect 6236 37204 6242 37216
rect 6825 37213 6837 37216
rect 6871 37213 6883 37247
rect 6825 37207 6883 37213
rect 7374 37204 7380 37256
rect 7432 37244 7438 37256
rect 7561 37247 7619 37253
rect 7561 37244 7573 37247
rect 7432 37216 7573 37244
rect 7432 37204 7438 37216
rect 7561 37213 7573 37216
rect 7607 37213 7619 37247
rect 7561 37207 7619 37213
rect 8662 37204 8668 37256
rect 8720 37244 8726 37256
rect 9401 37247 9459 37253
rect 9401 37244 9413 37247
rect 8720 37216 9413 37244
rect 8720 37204 8726 37216
rect 9401 37213 9413 37216
rect 9447 37244 9459 37247
rect 9582 37244 9588 37256
rect 9447 37216 9588 37244
rect 9447 37213 9459 37216
rect 9401 37207 9459 37213
rect 9582 37204 9588 37216
rect 9640 37204 9646 37256
rect 9858 37204 9864 37256
rect 9916 37244 9922 37256
rect 10137 37247 10195 37253
rect 10137 37244 10149 37247
rect 9916 37216 10149 37244
rect 9916 37204 9922 37216
rect 10137 37213 10149 37216
rect 10183 37213 10195 37247
rect 10137 37207 10195 37213
rect 11054 37204 11060 37256
rect 11112 37244 11118 37256
rect 12452 37253 12480 37284
rect 13446 37272 13452 37324
rect 13504 37312 13510 37324
rect 14093 37315 14151 37321
rect 14093 37312 14105 37315
rect 13504 37284 14105 37312
rect 13504 37272 13510 37284
rect 14093 37281 14105 37284
rect 14139 37281 14151 37315
rect 14093 37275 14151 37281
rect 18322 37272 18328 37324
rect 18380 37312 18386 37324
rect 19058 37312 19064 37324
rect 18380 37284 19064 37312
rect 18380 37272 18386 37284
rect 19058 37272 19064 37284
rect 19116 37312 19122 37324
rect 19245 37315 19303 37321
rect 19245 37312 19257 37315
rect 19116 37284 19257 37312
rect 19116 37272 19122 37284
rect 19245 37281 19257 37284
rect 19291 37281 19303 37315
rect 19245 37275 19303 37281
rect 20070 37272 20076 37324
rect 20128 37312 20134 37324
rect 23293 37315 23351 37321
rect 23293 37312 23305 37315
rect 20128 37284 23305 37312
rect 20128 37272 20134 37284
rect 23293 37281 23305 37284
rect 23339 37281 23351 37315
rect 24762 37312 24768 37324
rect 24723 37284 24768 37312
rect 23293 37275 23351 37281
rect 24762 37272 24768 37284
rect 24820 37272 24826 37324
rect 26878 37272 26884 37324
rect 26936 37312 26942 37324
rect 29840 37312 29868 37352
rect 32493 37349 32505 37352
rect 32539 37349 32551 37383
rect 35802 37380 35808 37392
rect 35763 37352 35808 37380
rect 32493 37343 32551 37349
rect 35802 37340 35808 37352
rect 35860 37340 35866 37392
rect 31389 37315 31447 37321
rect 31389 37312 31401 37315
rect 26936 37284 29868 37312
rect 30116 37284 31401 37312
rect 26936 37272 26942 37284
rect 11609 37247 11667 37253
rect 11609 37244 11621 37247
rect 11112 37216 11621 37244
rect 11112 37204 11118 37216
rect 11609 37213 11621 37216
rect 11655 37213 11667 37247
rect 11609 37207 11667 37213
rect 12437 37247 12495 37253
rect 12437 37213 12449 37247
rect 12483 37213 12495 37247
rect 13354 37244 13360 37256
rect 13315 37216 13360 37244
rect 12437 37207 12495 37213
rect 13354 37204 13360 37216
rect 13412 37204 13418 37256
rect 14369 37247 14427 37253
rect 14369 37213 14381 37247
rect 14415 37213 14427 37247
rect 15378 37244 15384 37256
rect 15339 37216 15384 37244
rect 14369 37207 14427 37213
rect 2406 37176 2412 37188
rect 1412 37148 2412 37176
rect 2406 37136 2412 37148
rect 2464 37136 2470 37188
rect 14384 37176 14412 37207
rect 15378 37204 15384 37216
rect 15436 37204 15442 37256
rect 15930 37204 15936 37256
rect 15988 37244 15994 37256
rect 16666 37244 16672 37256
rect 15988 37216 16672 37244
rect 15988 37204 15994 37216
rect 16666 37204 16672 37216
rect 16724 37204 16730 37256
rect 16945 37247 17003 37253
rect 16945 37213 16957 37247
rect 16991 37213 17003 37247
rect 16945 37207 17003 37213
rect 16114 37176 16120 37188
rect 14384 37148 16120 37176
rect 16114 37136 16120 37148
rect 16172 37136 16178 37188
rect 16574 37136 16580 37188
rect 16632 37176 16638 37188
rect 16960 37176 16988 37207
rect 17034 37204 17040 37256
rect 17092 37244 17098 37256
rect 17957 37247 18015 37253
rect 17957 37244 17969 37247
rect 17092 37216 17969 37244
rect 17092 37204 17098 37216
rect 17957 37213 17969 37216
rect 18003 37213 18015 37247
rect 17957 37207 18015 37213
rect 19521 37247 19579 37253
rect 19521 37213 19533 37247
rect 19567 37213 19579 37247
rect 19521 37207 19579 37213
rect 16632 37148 16988 37176
rect 16632 37136 16638 37148
rect 18598 37136 18604 37188
rect 18656 37176 18662 37188
rect 19536 37176 19564 37207
rect 20714 37204 20720 37256
rect 20772 37244 20778 37256
rect 20901 37247 20959 37253
rect 20901 37244 20913 37247
rect 20772 37216 20913 37244
rect 20772 37204 20778 37216
rect 20901 37213 20913 37216
rect 20947 37213 20959 37247
rect 20901 37207 20959 37213
rect 23198 37204 23204 37256
rect 23256 37244 23262 37256
rect 23382 37244 23388 37256
rect 23256 37216 23388 37244
rect 23256 37204 23262 37216
rect 23382 37204 23388 37216
rect 23440 37244 23446 37256
rect 23477 37247 23535 37253
rect 23477 37244 23489 37247
rect 23440 37216 23489 37244
rect 23440 37204 23446 37216
rect 23477 37213 23489 37216
rect 23523 37213 23535 37247
rect 23477 37207 23535 37213
rect 24394 37204 24400 37256
rect 24452 37244 24458 37256
rect 24949 37247 25007 37253
rect 24949 37244 24961 37247
rect 24452 37216 24961 37244
rect 24452 37204 24458 37216
rect 24949 37213 24961 37216
rect 24995 37213 25007 37247
rect 24949 37207 25007 37213
rect 25590 37204 25596 37256
rect 25648 37244 25654 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 25648 37216 25881 37244
rect 25648 37204 25654 37216
rect 25869 37213 25881 37216
rect 25915 37213 25927 37247
rect 25869 37207 25927 37213
rect 26786 37204 26792 37256
rect 26844 37244 26850 37256
rect 27522 37244 27528 37256
rect 26844 37216 27528 37244
rect 26844 37204 26850 37216
rect 27522 37204 27528 37216
rect 27580 37204 27586 37256
rect 27982 37204 27988 37256
rect 28040 37244 28046 37256
rect 28261 37247 28319 37253
rect 28261 37244 28273 37247
rect 28040 37216 28273 37244
rect 28040 37204 28046 37216
rect 28261 37213 28273 37216
rect 28307 37244 28319 37247
rect 28813 37247 28871 37253
rect 28813 37244 28825 37247
rect 28307 37216 28825 37244
rect 28307 37213 28319 37216
rect 28261 37207 28319 37213
rect 28813 37213 28825 37216
rect 28859 37213 28871 37247
rect 28813 37207 28871 37213
rect 29178 37204 29184 37256
rect 29236 37244 29242 37256
rect 30116 37253 30144 37284
rect 31389 37281 31401 37284
rect 31435 37281 31447 37315
rect 33965 37315 34023 37321
rect 33965 37312 33977 37315
rect 31389 37275 31447 37281
rect 32692 37284 33977 37312
rect 30101 37247 30159 37253
rect 30101 37244 30113 37247
rect 29236 37216 30113 37244
rect 29236 37204 29242 37216
rect 30101 37213 30113 37216
rect 30147 37213 30159 37247
rect 30101 37207 30159 37213
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30837 37247 30895 37253
rect 30837 37244 30849 37247
rect 30432 37216 30849 37244
rect 30432 37204 30438 37216
rect 30837 37213 30849 37216
rect 30883 37213 30895 37247
rect 30837 37207 30895 37213
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32692 37253 32720 37284
rect 33965 37281 33977 37284
rect 34011 37281 34023 37315
rect 36541 37315 36599 37321
rect 36541 37312 36553 37315
rect 33965 37275 34023 37281
rect 35268 37284 36553 37312
rect 32677 37247 32735 37253
rect 32677 37244 32689 37247
rect 31812 37216 32689 37244
rect 31812 37204 31818 37216
rect 32677 37213 32689 37216
rect 32723 37213 32735 37247
rect 32677 37207 32735 37213
rect 32858 37204 32864 37256
rect 32916 37244 32922 37256
rect 33134 37244 33140 37256
rect 32916 37216 33140 37244
rect 32916 37204 32922 37216
rect 33134 37204 33140 37216
rect 33192 37244 33198 37256
rect 33413 37247 33471 37253
rect 33413 37244 33425 37247
rect 33192 37216 33425 37244
rect 33192 37204 33198 37216
rect 33413 37213 33425 37216
rect 33459 37213 33471 37247
rect 33413 37207 33471 37213
rect 34054 37204 34060 37256
rect 34112 37244 34118 37256
rect 35268 37253 35296 37284
rect 36541 37281 36553 37284
rect 36587 37281 36599 37315
rect 36541 37275 36599 37281
rect 35253 37247 35311 37253
rect 35253 37244 35265 37247
rect 34112 37216 35265 37244
rect 34112 37204 34118 37216
rect 35253 37213 35265 37216
rect 35299 37213 35311 37247
rect 35253 37207 35311 37213
rect 35342 37204 35348 37256
rect 35400 37244 35406 37256
rect 35710 37244 35716 37256
rect 35400 37216 35716 37244
rect 35400 37204 35406 37216
rect 35710 37204 35716 37216
rect 35768 37244 35774 37256
rect 35989 37247 36047 37253
rect 35989 37244 36001 37247
rect 35768 37216 36001 37244
rect 35768 37204 35774 37216
rect 35989 37213 36001 37216
rect 36035 37213 36047 37247
rect 35989 37207 36047 37213
rect 37642 37204 37648 37256
rect 37700 37244 37706 37256
rect 38105 37247 38163 37253
rect 38105 37244 38117 37247
rect 37700 37216 38117 37244
rect 37700 37204 37706 37216
rect 38105 37213 38117 37216
rect 38151 37244 38163 37247
rect 38378 37244 38384 37256
rect 38151 37216 38384 37244
rect 38151 37213 38163 37216
rect 38105 37207 38163 37213
rect 38378 37204 38384 37216
rect 38436 37204 38442 37256
rect 38562 37204 38568 37256
rect 38620 37244 38626 37256
rect 38657 37247 38715 37253
rect 38657 37244 38669 37247
rect 38620 37216 38669 37244
rect 38620 37204 38626 37216
rect 38657 37213 38669 37216
rect 38703 37213 38715 37247
rect 38657 37207 38715 37213
rect 38930 37204 38936 37256
rect 38988 37244 38994 37256
rect 40126 37244 40132 37256
rect 38988 37216 40132 37244
rect 38988 37204 38994 37216
rect 40126 37204 40132 37216
rect 40184 37244 40190 37256
rect 40313 37247 40371 37253
rect 40313 37244 40325 37247
rect 40184 37216 40325 37244
rect 40184 37204 40190 37216
rect 40313 37213 40325 37216
rect 40359 37213 40371 37247
rect 40313 37207 40371 37213
rect 42334 37204 42340 37256
rect 42392 37244 42398 37256
rect 42429 37247 42487 37253
rect 42429 37244 42441 37247
rect 42392 37216 42441 37244
rect 42392 37204 42398 37216
rect 42429 37213 42441 37216
rect 42475 37213 42487 37247
rect 42429 37207 42487 37213
rect 43070 37204 43076 37256
rect 43128 37244 43134 37256
rect 43165 37247 43223 37253
rect 43165 37244 43177 37247
rect 43128 37216 43177 37244
rect 43128 37204 43134 37216
rect 43165 37213 43177 37216
rect 43211 37213 43223 37247
rect 43165 37207 43223 37213
rect 43438 37204 43444 37256
rect 43496 37244 43502 37256
rect 43901 37247 43959 37253
rect 43901 37244 43913 37247
rect 43496 37216 43913 37244
rect 43496 37204 43502 37216
rect 43901 37213 43913 37216
rect 43947 37213 43959 37247
rect 43901 37207 43959 37213
rect 18656 37148 19564 37176
rect 18656 37136 18662 37148
rect 22094 37136 22100 37188
rect 22152 37176 22158 37188
rect 22281 37179 22339 37185
rect 22281 37176 22293 37179
rect 22152 37148 22293 37176
rect 22152 37136 22158 37148
rect 22281 37145 22293 37148
rect 22327 37145 22339 37179
rect 22281 37139 22339 37145
rect 40218 37136 40224 37188
rect 40276 37176 40282 37188
rect 41506 37176 41512 37188
rect 40276 37148 41512 37176
rect 40276 37136 40282 37148
rect 41506 37136 41512 37148
rect 41564 37136 41570 37188
rect 1581 37111 1639 37117
rect 1581 37077 1593 37111
rect 1627 37108 1639 37111
rect 2590 37108 2596 37120
rect 1627 37080 2596 37108
rect 1627 37077 1639 37080
rect 1581 37071 1639 37077
rect 2590 37068 2596 37080
rect 2648 37068 2654 37120
rect 12618 37068 12624 37120
rect 12676 37108 12682 37120
rect 13173 37111 13231 37117
rect 13173 37108 13185 37111
rect 12676 37080 13185 37108
rect 12676 37068 12682 37080
rect 13173 37077 13185 37080
rect 13219 37077 13231 37111
rect 13173 37071 13231 37077
rect 15194 37068 15200 37120
rect 15252 37108 15258 37120
rect 15565 37111 15623 37117
rect 15565 37108 15577 37111
rect 15252 37080 15577 37108
rect 15252 37068 15258 37080
rect 15565 37077 15577 37080
rect 15611 37077 15623 37111
rect 15565 37071 15623 37077
rect 16298 37068 16304 37120
rect 16356 37108 16362 37120
rect 18141 37111 18199 37117
rect 18141 37108 18153 37111
rect 16356 37080 18153 37108
rect 16356 37068 16362 37080
rect 18141 37077 18153 37080
rect 18187 37077 18199 37111
rect 30742 37108 30748 37120
rect 30703 37080 30748 37108
rect 18141 37071 18199 37077
rect 30742 37068 30748 37080
rect 30800 37068 30806 37120
rect 38838 37108 38844 37120
rect 38799 37080 38844 37108
rect 38838 37068 38844 37080
rect 38896 37068 38902 37120
rect 41690 37068 41696 37120
rect 41748 37108 41754 37120
rect 42613 37111 42671 37117
rect 42613 37108 42625 37111
rect 41748 37080 42625 37108
rect 41748 37068 41754 37080
rect 42613 37077 42625 37080
rect 42659 37077 42671 37111
rect 42613 37071 42671 37077
rect 42886 37068 42892 37120
rect 42944 37108 42950 37120
rect 43349 37111 43407 37117
rect 43349 37108 43361 37111
rect 42944 37080 43361 37108
rect 42944 37068 42950 37080
rect 43349 37077 43361 37080
rect 43395 37077 43407 37111
rect 43349 37071 43407 37077
rect 44085 37111 44143 37117
rect 44085 37077 44097 37111
rect 44131 37108 44143 37111
rect 44174 37108 44180 37120
rect 44131 37080 44180 37108
rect 44131 37077 44143 37080
rect 44085 37071 44143 37077
rect 44174 37068 44180 37080
rect 44232 37068 44238 37120
rect 1104 37018 44896 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 44896 37018
rect 1104 36944 44896 36966
rect 566 36864 572 36916
rect 624 36904 630 36916
rect 1489 36907 1547 36913
rect 1489 36904 1501 36907
rect 624 36876 1501 36904
rect 624 36864 630 36876
rect 1489 36873 1501 36876
rect 1535 36873 1547 36907
rect 1489 36867 1547 36873
rect 1762 36864 1768 36916
rect 1820 36904 1826 36916
rect 2225 36907 2283 36913
rect 2225 36904 2237 36907
rect 1820 36876 2237 36904
rect 1820 36864 1826 36876
rect 2225 36873 2237 36876
rect 2271 36873 2283 36907
rect 2225 36867 2283 36873
rect 2958 36864 2964 36916
rect 3016 36904 3022 36916
rect 3145 36907 3203 36913
rect 3145 36904 3157 36907
rect 3016 36876 3157 36904
rect 3016 36864 3022 36876
rect 3145 36873 3157 36876
rect 3191 36873 3203 36907
rect 3145 36867 3203 36873
rect 4154 36864 4160 36916
rect 4212 36904 4218 36916
rect 4433 36907 4491 36913
rect 4433 36904 4445 36907
rect 4212 36876 4445 36904
rect 4212 36864 4218 36876
rect 4433 36873 4445 36876
rect 4479 36873 4491 36907
rect 4433 36867 4491 36873
rect 4798 36864 4804 36916
rect 4856 36904 4862 36916
rect 4985 36907 5043 36913
rect 4985 36904 4997 36907
rect 4856 36876 4997 36904
rect 4856 36864 4862 36876
rect 4985 36873 4997 36876
rect 5031 36873 5043 36907
rect 4985 36867 5043 36873
rect 5534 36864 5540 36916
rect 5592 36904 5598 36916
rect 5629 36907 5687 36913
rect 5629 36904 5641 36907
rect 5592 36876 5641 36904
rect 5592 36864 5598 36876
rect 5629 36873 5641 36876
rect 5675 36873 5687 36907
rect 5629 36867 5687 36873
rect 6638 36864 6644 36916
rect 6696 36904 6702 36916
rect 6825 36907 6883 36913
rect 6825 36904 6837 36907
rect 6696 36876 6837 36904
rect 6696 36864 6702 36876
rect 6825 36873 6837 36876
rect 6871 36873 6883 36907
rect 6825 36867 6883 36873
rect 7834 36864 7840 36916
rect 7892 36904 7898 36916
rect 8021 36907 8079 36913
rect 8021 36904 8033 36907
rect 7892 36876 8033 36904
rect 7892 36864 7898 36876
rect 8021 36873 8033 36876
rect 8067 36873 8079 36907
rect 8021 36867 8079 36873
rect 9030 36864 9036 36916
rect 9088 36904 9094 36916
rect 9217 36907 9275 36913
rect 9217 36904 9229 36907
rect 9088 36876 9229 36904
rect 9088 36864 9094 36876
rect 9217 36873 9229 36876
rect 9263 36873 9275 36907
rect 9217 36867 9275 36873
rect 9398 36864 9404 36916
rect 9456 36904 9462 36916
rect 9953 36907 10011 36913
rect 9953 36904 9965 36907
rect 9456 36876 9965 36904
rect 9456 36864 9462 36876
rect 9953 36873 9965 36876
rect 9999 36873 10011 36907
rect 9953 36867 10011 36873
rect 10686 36864 10692 36916
rect 10744 36904 10750 36916
rect 10781 36907 10839 36913
rect 10781 36904 10793 36907
rect 10744 36876 10793 36904
rect 10744 36864 10750 36876
rect 10781 36873 10793 36876
rect 10827 36873 10839 36907
rect 10781 36867 10839 36873
rect 11422 36864 11428 36916
rect 11480 36904 11486 36916
rect 12345 36907 12403 36913
rect 12345 36904 12357 36907
rect 11480 36876 12357 36904
rect 11480 36864 11486 36876
rect 12345 36873 12357 36876
rect 12391 36873 12403 36907
rect 12345 36867 12403 36873
rect 13078 36864 13084 36916
rect 13136 36904 13142 36916
rect 13265 36907 13323 36913
rect 13265 36904 13277 36907
rect 13136 36876 13277 36904
rect 13136 36864 13142 36876
rect 13265 36873 13277 36876
rect 13311 36873 13323 36907
rect 13265 36867 13323 36873
rect 13906 36864 13912 36916
rect 13964 36904 13970 36916
rect 14093 36907 14151 36913
rect 14093 36904 14105 36907
rect 13964 36876 14105 36904
rect 13964 36864 13970 36876
rect 14093 36873 14105 36876
rect 14139 36873 14151 36907
rect 16666 36904 16672 36916
rect 16627 36876 16672 36904
rect 14093 36867 14151 36873
rect 16666 36864 16672 36876
rect 16724 36864 16730 36916
rect 18690 36864 18696 36916
rect 18748 36904 18754 36916
rect 18877 36907 18935 36913
rect 18877 36904 18889 36907
rect 18748 36876 18889 36904
rect 18748 36864 18754 36876
rect 18877 36873 18889 36876
rect 18923 36873 18935 36907
rect 18877 36867 18935 36873
rect 20346 36864 20352 36916
rect 20404 36904 20410 36916
rect 21085 36907 21143 36913
rect 21085 36904 21097 36907
rect 20404 36876 21097 36904
rect 20404 36864 20410 36876
rect 21085 36873 21097 36876
rect 21131 36873 21143 36907
rect 21085 36867 21143 36873
rect 21174 36864 21180 36916
rect 21232 36904 21238 36916
rect 21913 36907 21971 36913
rect 21913 36904 21925 36907
rect 21232 36876 21925 36904
rect 21232 36864 21238 36876
rect 21913 36873 21925 36876
rect 21959 36873 21971 36907
rect 21913 36867 21971 36873
rect 22370 36864 22376 36916
rect 22428 36904 22434 36916
rect 22649 36907 22707 36913
rect 22649 36904 22661 36907
rect 22428 36876 22661 36904
rect 22428 36864 22434 36876
rect 22649 36873 22661 36876
rect 22695 36873 22707 36907
rect 22649 36867 22707 36873
rect 23566 36864 23572 36916
rect 23624 36904 23630 36916
rect 23845 36907 23903 36913
rect 23845 36904 23857 36907
rect 23624 36876 23857 36904
rect 23624 36864 23630 36876
rect 23845 36873 23857 36876
rect 23891 36873 23903 36907
rect 23845 36867 23903 36873
rect 24854 36864 24860 36916
rect 24912 36904 24918 36916
rect 24949 36907 25007 36913
rect 24949 36904 24961 36907
rect 24912 36876 24961 36904
rect 24912 36864 24918 36876
rect 24949 36873 24961 36876
rect 24995 36873 25007 36907
rect 24949 36867 25007 36873
rect 25958 36864 25964 36916
rect 26016 36904 26022 36916
rect 26237 36907 26295 36913
rect 26237 36904 26249 36907
rect 26016 36876 26249 36904
rect 26016 36864 26022 36876
rect 26237 36873 26249 36876
rect 26283 36873 26295 36907
rect 26237 36867 26295 36873
rect 27154 36864 27160 36916
rect 27212 36904 27218 36916
rect 27433 36907 27491 36913
rect 27433 36904 27445 36907
rect 27212 36876 27445 36904
rect 27212 36864 27218 36876
rect 27433 36873 27445 36876
rect 27479 36873 27491 36907
rect 27433 36867 27491 36873
rect 27522 36864 27528 36916
rect 27580 36904 27586 36916
rect 27985 36907 28043 36913
rect 27985 36904 27997 36907
rect 27580 36876 27997 36904
rect 27580 36864 27586 36876
rect 27985 36873 27997 36876
rect 28031 36873 28043 36907
rect 27985 36867 28043 36873
rect 28442 36864 28448 36916
rect 28500 36904 28506 36916
rect 28721 36907 28779 36913
rect 28721 36904 28733 36907
rect 28500 36876 28733 36904
rect 28500 36864 28506 36876
rect 28721 36873 28733 36876
rect 28767 36873 28779 36907
rect 28721 36867 28779 36873
rect 29638 36864 29644 36916
rect 29696 36904 29702 36916
rect 29917 36907 29975 36913
rect 29917 36904 29929 36907
rect 29696 36876 29929 36904
rect 29696 36864 29702 36876
rect 29917 36873 29929 36876
rect 29963 36873 29975 36907
rect 29917 36867 29975 36873
rect 30374 36864 30380 36916
rect 30432 36904 30438 36916
rect 30653 36907 30711 36913
rect 30653 36904 30665 36907
rect 30432 36876 30665 36904
rect 30432 36864 30438 36876
rect 30653 36873 30665 36876
rect 30699 36873 30711 36907
rect 30653 36867 30711 36873
rect 30834 36864 30840 36916
rect 30892 36904 30898 36916
rect 31389 36907 31447 36913
rect 31389 36904 31401 36907
rect 30892 36876 31401 36904
rect 30892 36864 30898 36876
rect 31389 36873 31401 36876
rect 31435 36873 31447 36907
rect 31389 36867 31447 36873
rect 32030 36864 32036 36916
rect 32088 36904 32094 36916
rect 32309 36907 32367 36913
rect 32309 36904 32321 36907
rect 32088 36876 32321 36904
rect 32088 36864 32094 36876
rect 32309 36873 32321 36876
rect 32355 36873 32367 36907
rect 32309 36867 32367 36873
rect 32398 36864 32404 36916
rect 32456 36904 32462 36916
rect 33045 36907 33103 36913
rect 33045 36904 33057 36907
rect 32456 36876 33057 36904
rect 32456 36864 32462 36876
rect 33045 36873 33057 36876
rect 33091 36873 33103 36907
rect 33045 36867 33103 36873
rect 33226 36864 33232 36916
rect 33284 36904 33290 36916
rect 33873 36907 33931 36913
rect 33873 36904 33885 36907
rect 33284 36876 33885 36904
rect 33284 36864 33290 36876
rect 33873 36873 33885 36876
rect 33919 36873 33931 36907
rect 33873 36867 33931 36873
rect 34514 36864 34520 36916
rect 34572 36904 34578 36916
rect 34701 36907 34759 36913
rect 34701 36904 34713 36907
rect 34572 36876 34713 36904
rect 34572 36864 34578 36876
rect 34701 36873 34713 36876
rect 34747 36873 34759 36907
rect 34701 36867 34759 36873
rect 35618 36864 35624 36916
rect 35676 36904 35682 36916
rect 35805 36907 35863 36913
rect 35805 36904 35817 36907
rect 35676 36876 35817 36904
rect 35676 36864 35682 36876
rect 35805 36873 35817 36876
rect 35851 36873 35863 36907
rect 35805 36867 35863 36873
rect 36078 36864 36084 36916
rect 36136 36904 36142 36916
rect 36633 36907 36691 36913
rect 36633 36904 36645 36907
rect 36136 36876 36645 36904
rect 36136 36864 36142 36876
rect 36633 36873 36645 36876
rect 36679 36873 36691 36907
rect 36633 36867 36691 36873
rect 37274 36864 37280 36916
rect 37332 36904 37338 36916
rect 38197 36907 38255 36913
rect 38197 36904 38209 36907
rect 37332 36876 38209 36904
rect 37332 36864 37338 36876
rect 38197 36873 38209 36876
rect 38243 36873 38255 36907
rect 38197 36867 38255 36873
rect 38378 36864 38384 36916
rect 38436 36904 38442 36916
rect 38749 36907 38807 36913
rect 38749 36904 38761 36907
rect 38436 36876 38761 36904
rect 38436 36864 38442 36876
rect 38749 36873 38761 36876
rect 38795 36873 38807 36907
rect 38749 36867 38807 36873
rect 39298 36864 39304 36916
rect 39356 36904 39362 36916
rect 39577 36907 39635 36913
rect 39577 36904 39589 36907
rect 39356 36876 39589 36904
rect 39356 36864 39362 36876
rect 39577 36873 39589 36876
rect 39623 36873 39635 36907
rect 39577 36867 39635 36873
rect 40494 36864 40500 36916
rect 40552 36904 40558 36916
rect 40773 36907 40831 36913
rect 40773 36904 40785 36907
rect 40552 36876 40785 36904
rect 40552 36864 40558 36876
rect 40773 36873 40785 36876
rect 40819 36873 40831 36907
rect 40773 36867 40831 36873
rect 42150 36864 42156 36916
rect 42208 36904 42214 36916
rect 42613 36907 42671 36913
rect 42613 36904 42625 36907
rect 42208 36876 42625 36904
rect 42208 36864 42214 36876
rect 42613 36873 42625 36876
rect 42659 36873 42671 36907
rect 43346 36904 43352 36916
rect 43307 36876 43352 36904
rect 42613 36867 42671 36873
rect 43346 36864 43352 36876
rect 43404 36864 43410 36916
rect 44085 36907 44143 36913
rect 44085 36873 44097 36907
rect 44131 36904 44143 36907
rect 45370 36904 45376 36916
rect 44131 36876 45376 36904
rect 44131 36873 44143 36876
rect 44085 36867 44143 36873
rect 45370 36864 45376 36876
rect 45428 36864 45434 36916
rect 1302 36796 1308 36848
rect 1360 36836 1366 36848
rect 1360 36808 2452 36836
rect 1360 36796 1366 36808
rect 2424 36777 2452 36808
rect 1673 36771 1731 36777
rect 1673 36737 1685 36771
rect 1719 36737 1731 36771
rect 1673 36731 1731 36737
rect 2409 36771 2467 36777
rect 2409 36737 2421 36771
rect 2455 36737 2467 36771
rect 2409 36731 2467 36737
rect 3329 36771 3387 36777
rect 3329 36737 3341 36771
rect 3375 36768 3387 36771
rect 3878 36768 3884 36780
rect 3375 36740 3884 36768
rect 3375 36737 3387 36740
rect 3329 36731 3387 36737
rect 1688 36700 1716 36731
rect 3878 36728 3884 36740
rect 3936 36728 3942 36780
rect 4249 36771 4307 36777
rect 4249 36737 4261 36771
rect 4295 36768 4307 36771
rect 4706 36768 4712 36780
rect 4295 36740 4712 36768
rect 4295 36737 4307 36740
rect 4249 36731 4307 36737
rect 4706 36728 4712 36740
rect 4764 36728 4770 36780
rect 5813 36771 5871 36777
rect 5813 36737 5825 36771
rect 5859 36768 5871 36771
rect 6454 36768 6460 36780
rect 5859 36740 6460 36768
rect 5859 36737 5871 36740
rect 5813 36731 5871 36737
rect 6454 36728 6460 36740
rect 6512 36728 6518 36780
rect 7009 36771 7067 36777
rect 7009 36737 7021 36771
rect 7055 36737 7067 36771
rect 7009 36731 7067 36737
rect 8205 36771 8263 36777
rect 8205 36737 8217 36771
rect 8251 36768 8263 36771
rect 8662 36768 8668 36780
rect 8251 36740 8668 36768
rect 8251 36737 8263 36740
rect 8205 36731 8263 36737
rect 2498 36700 2504 36712
rect 1688 36672 2504 36700
rect 2498 36660 2504 36672
rect 2556 36660 2562 36712
rect 7024 36564 7052 36731
rect 8662 36728 8668 36740
rect 8720 36728 8726 36780
rect 9401 36771 9459 36777
rect 9401 36737 9413 36771
rect 9447 36768 9459 36771
rect 9490 36768 9496 36780
rect 9447 36740 9496 36768
rect 9447 36737 9459 36740
rect 9401 36731 9459 36737
rect 9490 36728 9496 36740
rect 9548 36728 9554 36780
rect 10137 36771 10195 36777
rect 10137 36737 10149 36771
rect 10183 36737 10195 36771
rect 10962 36768 10968 36780
rect 10923 36740 10968 36768
rect 10137 36731 10195 36737
rect 10152 36700 10180 36731
rect 10962 36728 10968 36740
rect 11020 36728 11026 36780
rect 11793 36771 11851 36777
rect 11793 36737 11805 36771
rect 11839 36768 11851 36771
rect 11974 36768 11980 36780
rect 11839 36740 11980 36768
rect 11839 36737 11851 36740
rect 11793 36731 11851 36737
rect 11974 36728 11980 36740
rect 12032 36728 12038 36780
rect 12529 36771 12587 36777
rect 12529 36737 12541 36771
rect 12575 36768 12587 36771
rect 12618 36768 12624 36780
rect 12575 36740 12624 36768
rect 12575 36737 12587 36740
rect 12529 36731 12587 36737
rect 12618 36728 12624 36740
rect 12676 36728 12682 36780
rect 13449 36771 13507 36777
rect 13449 36737 13461 36771
rect 13495 36768 13507 36771
rect 13722 36768 13728 36780
rect 13495 36740 13728 36768
rect 13495 36737 13507 36740
rect 13449 36731 13507 36737
rect 13722 36728 13728 36740
rect 13780 36728 13786 36780
rect 14277 36771 14335 36777
rect 14277 36737 14289 36771
rect 14323 36768 14335 36771
rect 14458 36768 14464 36780
rect 14323 36740 14464 36768
rect 14323 36737 14335 36740
rect 14277 36731 14335 36737
rect 14458 36728 14464 36740
rect 14516 36728 14522 36780
rect 15289 36771 15347 36777
rect 15289 36737 15301 36771
rect 15335 36768 15347 36771
rect 15654 36768 15660 36780
rect 15335 36740 15660 36768
rect 15335 36737 15347 36740
rect 15289 36731 15347 36737
rect 15654 36728 15660 36740
rect 15712 36728 15718 36780
rect 17126 36728 17132 36780
rect 17184 36768 17190 36780
rect 17221 36771 17279 36777
rect 17221 36768 17233 36771
rect 17184 36740 17233 36768
rect 17184 36728 17190 36740
rect 17221 36737 17233 36740
rect 17267 36737 17279 36771
rect 17221 36731 17279 36737
rect 18230 36728 18236 36780
rect 18288 36768 18294 36780
rect 19061 36771 19119 36777
rect 19061 36768 19073 36771
rect 18288 36740 19073 36768
rect 18288 36728 18294 36740
rect 19061 36737 19073 36740
rect 19107 36737 19119 36771
rect 19061 36731 19119 36737
rect 19426 36728 19432 36780
rect 19484 36768 19490 36780
rect 19613 36771 19671 36777
rect 19613 36768 19625 36771
rect 19484 36740 19625 36768
rect 19484 36728 19490 36740
rect 19613 36737 19625 36740
rect 19659 36737 19671 36771
rect 19613 36731 19671 36737
rect 20622 36728 20628 36780
rect 20680 36768 20686 36780
rect 20901 36771 20959 36777
rect 20901 36768 20913 36771
rect 20680 36740 20913 36768
rect 20680 36728 20686 36740
rect 20901 36737 20913 36740
rect 20947 36737 20959 36771
rect 20901 36731 20959 36737
rect 22097 36771 22155 36777
rect 22097 36737 22109 36771
rect 22143 36768 22155 36771
rect 22646 36768 22652 36780
rect 22143 36740 22652 36768
rect 22143 36737 22155 36740
rect 22097 36731 22155 36737
rect 22646 36728 22652 36740
rect 22704 36728 22710 36780
rect 22833 36771 22891 36777
rect 22833 36737 22845 36771
rect 22879 36768 22891 36771
rect 23198 36768 23204 36780
rect 22879 36740 23204 36768
rect 22879 36737 22891 36740
rect 22833 36731 22891 36737
rect 23198 36728 23204 36740
rect 23256 36728 23262 36780
rect 23658 36768 23664 36780
rect 23619 36740 23664 36768
rect 23658 36728 23664 36740
rect 23716 36728 23722 36780
rect 25133 36771 25191 36777
rect 25133 36737 25145 36771
rect 25179 36768 25191 36771
rect 25222 36768 25228 36780
rect 25179 36740 25228 36768
rect 25179 36737 25191 36740
rect 25133 36731 25191 36737
rect 25222 36728 25228 36740
rect 25280 36728 25286 36780
rect 26050 36768 26056 36780
rect 26011 36740 26056 36768
rect 26050 36728 26056 36740
rect 26108 36728 26114 36780
rect 27062 36728 27068 36780
rect 27120 36768 27126 36780
rect 27249 36771 27307 36777
rect 27249 36768 27261 36771
rect 27120 36740 27261 36768
rect 27120 36728 27126 36740
rect 27249 36737 27261 36740
rect 27295 36737 27307 36771
rect 28534 36768 28540 36780
rect 28495 36740 28540 36768
rect 27249 36731 27307 36737
rect 28534 36728 28540 36740
rect 28592 36728 28598 36780
rect 29546 36728 29552 36780
rect 29604 36768 29610 36780
rect 29733 36771 29791 36777
rect 29733 36768 29745 36771
rect 29604 36740 29745 36768
rect 29604 36728 29610 36740
rect 29733 36737 29745 36740
rect 29779 36737 29791 36771
rect 29733 36731 29791 36737
rect 30374 36728 30380 36780
rect 30432 36768 30438 36780
rect 30469 36771 30527 36777
rect 30469 36768 30481 36771
rect 30432 36740 30481 36768
rect 30432 36728 30438 36740
rect 30469 36737 30481 36740
rect 30515 36737 30527 36771
rect 30469 36731 30527 36737
rect 31018 36728 31024 36780
rect 31076 36768 31082 36780
rect 31205 36771 31263 36777
rect 31205 36768 31217 36771
rect 31076 36740 31217 36768
rect 31076 36728 31082 36740
rect 31205 36737 31217 36740
rect 31251 36737 31263 36771
rect 32122 36768 32128 36780
rect 32083 36740 32128 36768
rect 31205 36731 31263 36737
rect 32122 36728 32128 36740
rect 32180 36728 32186 36780
rect 32674 36728 32680 36780
rect 32732 36768 32738 36780
rect 32861 36771 32919 36777
rect 32861 36768 32873 36771
rect 32732 36740 32873 36768
rect 32732 36728 32738 36740
rect 32861 36737 32873 36740
rect 32907 36737 32919 36771
rect 32861 36731 32919 36737
rect 33502 36728 33508 36780
rect 33560 36768 33566 36780
rect 33689 36771 33747 36777
rect 33689 36768 33701 36771
rect 33560 36740 33701 36768
rect 33560 36728 33566 36740
rect 33689 36737 33701 36740
rect 33735 36737 33747 36771
rect 33689 36731 33747 36737
rect 34238 36728 34244 36780
rect 34296 36768 34302 36780
rect 34517 36771 34575 36777
rect 34517 36768 34529 36771
rect 34296 36740 34529 36768
rect 34296 36728 34302 36740
rect 34517 36737 34529 36740
rect 34563 36737 34575 36771
rect 35986 36768 35992 36780
rect 35947 36740 35992 36768
rect 34517 36731 34575 36737
rect 35986 36728 35992 36740
rect 36044 36728 36050 36780
rect 36262 36728 36268 36780
rect 36320 36768 36326 36780
rect 36449 36771 36507 36777
rect 36449 36768 36461 36771
rect 36320 36740 36461 36768
rect 36320 36728 36326 36740
rect 36449 36737 36461 36740
rect 36495 36737 36507 36771
rect 36449 36731 36507 36737
rect 36538 36728 36544 36780
rect 36596 36768 36602 36780
rect 37090 36768 37096 36780
rect 36596 36740 37096 36768
rect 36596 36728 36602 36740
rect 37090 36728 37096 36740
rect 37148 36768 37154 36780
rect 37461 36771 37519 36777
rect 37461 36768 37473 36771
rect 37148 36740 37473 36768
rect 37148 36728 37154 36740
rect 37461 36737 37473 36740
rect 37507 36737 37519 36771
rect 37461 36731 37519 36737
rect 37826 36728 37832 36780
rect 37884 36768 37890 36780
rect 38013 36771 38071 36777
rect 38013 36768 38025 36771
rect 37884 36740 38025 36768
rect 37884 36728 37890 36740
rect 38013 36737 38025 36740
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 39206 36728 39212 36780
rect 39264 36768 39270 36780
rect 39393 36771 39451 36777
rect 39393 36768 39405 36771
rect 39264 36740 39405 36768
rect 39264 36728 39270 36740
rect 39393 36737 39405 36740
rect 39439 36737 39451 36771
rect 40586 36768 40592 36780
rect 40547 36740 40592 36768
rect 39393 36731 39451 36737
rect 40586 36728 40592 36740
rect 40644 36728 40650 36780
rect 41414 36728 41420 36780
rect 41472 36768 41478 36780
rect 41601 36771 41659 36777
rect 41601 36768 41613 36771
rect 41472 36740 41613 36768
rect 41472 36728 41478 36740
rect 41601 36737 41613 36740
rect 41647 36737 41659 36771
rect 42426 36768 42432 36780
rect 42387 36740 42432 36768
rect 41601 36731 41659 36737
rect 42426 36728 42432 36740
rect 42484 36728 42490 36780
rect 43162 36768 43168 36780
rect 43123 36740 43168 36768
rect 43162 36728 43168 36740
rect 43220 36728 43226 36780
rect 43530 36728 43536 36780
rect 43588 36768 43594 36780
rect 43901 36771 43959 36777
rect 43901 36768 43913 36771
rect 43588 36740 43913 36768
rect 43588 36728 43594 36740
rect 43901 36737 43913 36740
rect 43947 36737 43959 36771
rect 43901 36731 43959 36737
rect 10870 36700 10876 36712
rect 10152 36672 10876 36700
rect 10870 36660 10876 36672
rect 10928 36660 10934 36712
rect 15194 36660 15200 36712
rect 15252 36700 15258 36712
rect 15565 36703 15623 36709
rect 15565 36700 15577 36703
rect 15252 36672 15577 36700
rect 15252 36660 15258 36672
rect 15565 36669 15577 36672
rect 15611 36700 15623 36703
rect 16025 36703 16083 36709
rect 16025 36700 16037 36703
rect 15611 36672 16037 36700
rect 15611 36669 15623 36672
rect 15565 36663 15623 36669
rect 16025 36669 16037 36672
rect 16071 36669 16083 36703
rect 17494 36700 17500 36712
rect 17455 36672 17500 36700
rect 16025 36663 16083 36669
rect 17494 36660 17500 36672
rect 17552 36660 17558 36712
rect 19886 36700 19892 36712
rect 19847 36672 19892 36700
rect 19886 36660 19892 36672
rect 19944 36660 19950 36712
rect 10226 36592 10232 36644
rect 10284 36632 10290 36644
rect 11609 36635 11667 36641
rect 11609 36632 11621 36635
rect 10284 36604 11621 36632
rect 10284 36592 10290 36604
rect 11609 36601 11621 36604
rect 11655 36601 11667 36635
rect 37274 36632 37280 36644
rect 37235 36604 37280 36632
rect 11609 36595 11667 36601
rect 37274 36592 37280 36604
rect 37332 36592 37338 36644
rect 10778 36564 10784 36576
rect 7024 36536 10784 36564
rect 10778 36524 10784 36536
rect 10836 36524 10842 36576
rect 41509 36567 41567 36573
rect 41509 36533 41521 36567
rect 41555 36564 41567 36567
rect 41598 36564 41604 36576
rect 41555 36536 41604 36564
rect 41555 36533 41567 36536
rect 41509 36527 41567 36533
rect 41598 36524 41604 36536
rect 41656 36524 41662 36576
rect 1104 36474 44896 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 44896 36474
rect 1104 36400 44896 36422
rect 934 36320 940 36372
rect 992 36360 998 36372
rect 1489 36363 1547 36369
rect 1489 36360 1501 36363
rect 992 36332 1501 36360
rect 992 36320 998 36332
rect 1489 36329 1501 36332
rect 1535 36329 1547 36363
rect 1489 36323 1547 36329
rect 2130 36320 2136 36372
rect 2188 36360 2194 36372
rect 2317 36363 2375 36369
rect 2317 36360 2329 36363
rect 2188 36332 2329 36360
rect 2188 36320 2194 36332
rect 2317 36329 2329 36332
rect 2363 36329 2375 36363
rect 2317 36323 2375 36329
rect 3418 36320 3424 36372
rect 3476 36360 3482 36372
rect 3881 36363 3939 36369
rect 3881 36360 3893 36363
rect 3476 36332 3893 36360
rect 3476 36320 3482 36332
rect 3881 36329 3893 36332
rect 3927 36329 3939 36363
rect 3881 36323 3939 36329
rect 4614 36320 4620 36372
rect 4672 36360 4678 36372
rect 4801 36363 4859 36369
rect 4801 36360 4813 36363
rect 4672 36332 4813 36360
rect 4672 36320 4678 36332
rect 4801 36329 4813 36332
rect 4847 36329 4859 36363
rect 4801 36323 4859 36329
rect 5810 36320 5816 36372
rect 5868 36360 5874 36372
rect 5997 36363 6055 36369
rect 5997 36360 6009 36363
rect 5868 36332 6009 36360
rect 5868 36320 5874 36332
rect 5997 36329 6009 36332
rect 6043 36329 6055 36363
rect 5997 36323 6055 36329
rect 7006 36320 7012 36372
rect 7064 36360 7070 36372
rect 7193 36363 7251 36369
rect 7193 36360 7205 36363
rect 7064 36332 7205 36360
rect 7064 36320 7070 36332
rect 7193 36329 7205 36332
rect 7239 36329 7251 36363
rect 7193 36323 7251 36329
rect 7374 36320 7380 36372
rect 7432 36360 7438 36372
rect 7837 36363 7895 36369
rect 7837 36360 7849 36363
rect 7432 36332 7849 36360
rect 7432 36320 7438 36332
rect 7837 36329 7849 36332
rect 7883 36329 7895 36363
rect 7837 36323 7895 36329
rect 8294 36320 8300 36372
rect 8352 36360 8358 36372
rect 9033 36363 9091 36369
rect 9033 36360 9045 36363
rect 8352 36332 9045 36360
rect 8352 36320 8358 36332
rect 9033 36329 9045 36332
rect 9079 36329 9091 36363
rect 9033 36323 9091 36329
rect 9582 36320 9588 36372
rect 9640 36360 9646 36372
rect 9677 36363 9735 36369
rect 9677 36360 9689 36363
rect 9640 36332 9689 36360
rect 9640 36320 9646 36332
rect 9677 36329 9689 36332
rect 9723 36329 9735 36363
rect 9677 36323 9735 36329
rect 9858 36320 9864 36372
rect 9916 36360 9922 36372
rect 10229 36363 10287 36369
rect 10229 36360 10241 36363
rect 9916 36332 10241 36360
rect 9916 36320 9922 36332
rect 10229 36329 10241 36332
rect 10275 36329 10287 36363
rect 10229 36323 10287 36329
rect 11054 36320 11060 36372
rect 11112 36360 11118 36372
rect 11333 36363 11391 36369
rect 11333 36360 11345 36363
rect 11112 36332 11345 36360
rect 11112 36320 11118 36332
rect 11333 36329 11345 36332
rect 11379 36329 11391 36363
rect 11333 36323 11391 36329
rect 11882 36320 11888 36372
rect 11940 36360 11946 36372
rect 12345 36363 12403 36369
rect 12345 36360 12357 36363
rect 11940 36332 12357 36360
rect 11940 36320 11946 36332
rect 12345 36329 12357 36332
rect 12391 36329 12403 36363
rect 13446 36360 13452 36372
rect 13407 36332 13452 36360
rect 12345 36323 12403 36329
rect 13446 36320 13452 36332
rect 13504 36320 13510 36372
rect 14274 36320 14280 36372
rect 14332 36360 14338 36372
rect 14553 36363 14611 36369
rect 14553 36360 14565 36363
rect 14332 36332 14565 36360
rect 14332 36320 14338 36332
rect 14553 36329 14565 36332
rect 14599 36329 14611 36363
rect 14553 36323 14611 36329
rect 15470 36320 15476 36372
rect 15528 36360 15534 36372
rect 15749 36363 15807 36369
rect 15749 36360 15761 36363
rect 15528 36332 15761 36360
rect 15528 36320 15534 36332
rect 15749 36329 15761 36332
rect 15795 36329 15807 36363
rect 15749 36323 15807 36329
rect 16758 36320 16764 36372
rect 16816 36360 16822 36372
rect 16853 36363 16911 36369
rect 16853 36360 16865 36363
rect 16816 36332 16865 36360
rect 16816 36320 16822 36332
rect 16853 36329 16865 36332
rect 16899 36329 16911 36363
rect 16853 36323 16911 36329
rect 17586 36320 17592 36372
rect 17644 36360 17650 36372
rect 17773 36363 17831 36369
rect 17773 36360 17785 36363
rect 17644 36332 17785 36360
rect 17644 36320 17650 36332
rect 17773 36329 17785 36332
rect 17819 36329 17831 36363
rect 17773 36323 17831 36329
rect 17954 36320 17960 36372
rect 18012 36360 18018 36372
rect 18509 36363 18567 36369
rect 18509 36360 18521 36363
rect 18012 36332 18521 36360
rect 18012 36320 18018 36332
rect 18509 36329 18521 36332
rect 18555 36329 18567 36363
rect 18509 36323 18567 36329
rect 19978 36320 19984 36372
rect 20036 36360 20042 36372
rect 20073 36363 20131 36369
rect 20073 36360 20085 36363
rect 20036 36332 20085 36360
rect 20036 36320 20042 36332
rect 20073 36329 20085 36332
rect 20119 36329 20131 36363
rect 20714 36360 20720 36372
rect 20675 36332 20720 36360
rect 20073 36323 20131 36329
rect 20714 36320 20720 36332
rect 20772 36320 20778 36372
rect 21542 36320 21548 36372
rect 21600 36360 21606 36372
rect 21729 36363 21787 36369
rect 21729 36360 21741 36363
rect 21600 36332 21741 36360
rect 21600 36320 21606 36332
rect 21729 36329 21741 36332
rect 21775 36329 21787 36363
rect 21729 36323 21787 36329
rect 22738 36320 22744 36372
rect 22796 36360 22802 36372
rect 22925 36363 22983 36369
rect 22925 36360 22937 36363
rect 22796 36332 22937 36360
rect 22796 36320 22802 36332
rect 22925 36329 22937 36332
rect 22971 36329 22983 36363
rect 22925 36323 22983 36329
rect 23382 36320 23388 36372
rect 23440 36360 23446 36372
rect 23569 36363 23627 36369
rect 23569 36360 23581 36363
rect 23440 36332 23581 36360
rect 23440 36320 23446 36332
rect 23569 36329 23581 36332
rect 23615 36329 23627 36363
rect 23569 36323 23627 36329
rect 23934 36320 23940 36372
rect 23992 36360 23998 36372
rect 24581 36363 24639 36369
rect 24581 36360 24593 36363
rect 23992 36332 24593 36360
rect 23992 36320 23998 36332
rect 24581 36329 24593 36332
rect 24627 36329 24639 36363
rect 24581 36323 24639 36329
rect 25130 36320 25136 36372
rect 25188 36360 25194 36372
rect 25409 36363 25467 36369
rect 25409 36360 25421 36363
rect 25188 36332 25421 36360
rect 25188 36320 25194 36332
rect 25409 36329 25421 36332
rect 25455 36329 25467 36363
rect 25409 36323 25467 36329
rect 25590 36320 25596 36372
rect 25648 36360 25654 36372
rect 25961 36363 26019 36369
rect 25961 36360 25973 36363
rect 25648 36332 25973 36360
rect 25648 36320 25654 36332
rect 25961 36329 25973 36332
rect 26007 36329 26019 36363
rect 25961 36323 26019 36329
rect 26418 36320 26424 36372
rect 26476 36360 26482 36372
rect 26697 36363 26755 36369
rect 26697 36360 26709 36363
rect 26476 36332 26709 36360
rect 26476 36320 26482 36332
rect 26697 36329 26709 36332
rect 26743 36329 26755 36363
rect 26697 36323 26755 36329
rect 27614 36320 27620 36372
rect 27672 36360 27678 36372
rect 27893 36363 27951 36369
rect 27893 36360 27905 36363
rect 27672 36332 27905 36360
rect 27672 36320 27678 36332
rect 27893 36329 27905 36332
rect 27939 36329 27951 36363
rect 28534 36360 28540 36372
rect 28495 36332 28540 36360
rect 27893 36323 27951 36329
rect 28534 36320 28540 36332
rect 28592 36320 28598 36372
rect 30466 36360 30472 36372
rect 30427 36332 30472 36360
rect 30466 36320 30472 36332
rect 30524 36320 30530 36372
rect 31202 36320 31208 36372
rect 31260 36360 31266 36372
rect 31481 36363 31539 36369
rect 31481 36360 31493 36363
rect 31260 36332 31493 36360
rect 31260 36320 31266 36332
rect 31481 36329 31493 36332
rect 31527 36329 31539 36363
rect 33134 36360 33140 36372
rect 33095 36332 33140 36360
rect 31481 36323 31539 36329
rect 33134 36320 33140 36332
rect 33192 36320 33198 36372
rect 33686 36320 33692 36372
rect 33744 36360 33750 36372
rect 33965 36363 34023 36369
rect 33965 36360 33977 36363
rect 33744 36332 33977 36360
rect 33744 36320 33750 36332
rect 33965 36329 33977 36332
rect 34011 36329 34023 36363
rect 33965 36323 34023 36329
rect 34790 36320 34796 36372
rect 34848 36360 34854 36372
rect 35161 36363 35219 36369
rect 35161 36360 35173 36363
rect 34848 36332 35173 36360
rect 34848 36320 34854 36332
rect 35161 36329 35173 36332
rect 35207 36329 35219 36363
rect 35710 36360 35716 36372
rect 35671 36332 35716 36360
rect 35161 36323 35219 36329
rect 35710 36320 35716 36332
rect 35768 36320 35774 36372
rect 35986 36320 35992 36372
rect 36044 36360 36050 36372
rect 36265 36363 36323 36369
rect 36265 36360 36277 36363
rect 36044 36332 36277 36360
rect 36044 36320 36050 36332
rect 36265 36329 36277 36332
rect 36311 36329 36323 36363
rect 37090 36360 37096 36372
rect 37051 36332 37096 36360
rect 36265 36323 36323 36329
rect 37090 36320 37096 36332
rect 37148 36320 37154 36372
rect 37366 36320 37372 36372
rect 37424 36360 37430 36372
rect 38197 36363 38255 36369
rect 38197 36360 38209 36363
rect 37424 36332 38209 36360
rect 37424 36320 37430 36332
rect 38197 36329 38209 36332
rect 38243 36329 38255 36363
rect 40034 36360 40040 36372
rect 39995 36332 40040 36360
rect 38197 36323 38255 36329
rect 40034 36320 40040 36332
rect 40092 36320 40098 36372
rect 40862 36320 40868 36372
rect 40920 36360 40926 36372
rect 41141 36363 41199 36369
rect 41141 36360 41153 36363
rect 40920 36332 41153 36360
rect 40920 36320 40926 36332
rect 41141 36329 41153 36332
rect 41187 36329 41199 36363
rect 41141 36323 41199 36329
rect 41506 36320 41512 36372
rect 41564 36360 41570 36372
rect 41693 36363 41751 36369
rect 41693 36360 41705 36363
rect 41564 36332 41705 36360
rect 41564 36320 41570 36332
rect 41693 36329 41705 36332
rect 41739 36329 41751 36363
rect 42334 36360 42340 36372
rect 42295 36332 42340 36360
rect 41693 36323 41751 36329
rect 42334 36320 42340 36332
rect 42392 36320 42398 36372
rect 43070 36360 43076 36372
rect 43031 36332 43076 36360
rect 43070 36320 43076 36332
rect 43128 36320 43134 36372
rect 44085 36363 44143 36369
rect 44085 36329 44097 36363
rect 44131 36360 44143 36363
rect 44542 36360 44548 36372
rect 44131 36332 44548 36360
rect 44131 36329 44143 36332
rect 44085 36323 44143 36329
rect 44542 36320 44548 36332
rect 44600 36320 44606 36372
rect 4614 36224 4620 36236
rect 2516 36196 4620 36224
rect 2516 36165 2544 36196
rect 4614 36184 4620 36196
rect 4672 36184 4678 36236
rect 1673 36159 1731 36165
rect 1673 36125 1685 36159
rect 1719 36125 1731 36159
rect 1673 36119 1731 36125
rect 2501 36159 2559 36165
rect 2501 36125 2513 36159
rect 2547 36125 2559 36159
rect 3142 36156 3148 36168
rect 3103 36128 3148 36156
rect 2501 36119 2559 36125
rect 1688 36088 1716 36119
rect 3142 36116 3148 36128
rect 3200 36116 3206 36168
rect 4065 36159 4123 36165
rect 4065 36125 4077 36159
rect 4111 36125 4123 36159
rect 4982 36156 4988 36168
rect 4943 36128 4988 36156
rect 4065 36119 4123 36125
rect 3234 36088 3240 36100
rect 1688 36060 3240 36088
rect 3234 36048 3240 36060
rect 3292 36048 3298 36100
rect 4080 36088 4108 36119
rect 4982 36116 4988 36128
rect 5040 36116 5046 36168
rect 6181 36159 6239 36165
rect 6181 36125 6193 36159
rect 6227 36156 6239 36159
rect 6914 36156 6920 36168
rect 6227 36128 6920 36156
rect 6227 36125 6239 36128
rect 6181 36119 6239 36125
rect 6914 36116 6920 36128
rect 6972 36116 6978 36168
rect 7374 36156 7380 36168
rect 7335 36128 7380 36156
rect 7374 36116 7380 36128
rect 7432 36116 7438 36168
rect 9217 36159 9275 36165
rect 9217 36125 9229 36159
rect 9263 36156 9275 36159
rect 10134 36156 10140 36168
rect 9263 36128 10140 36156
rect 9263 36125 9275 36128
rect 9217 36119 9275 36125
rect 10134 36116 10140 36128
rect 10192 36116 10198 36168
rect 12529 36159 12587 36165
rect 12529 36125 12541 36159
rect 12575 36156 12587 36159
rect 13170 36156 13176 36168
rect 12575 36128 13176 36156
rect 12575 36125 12587 36128
rect 12529 36119 12587 36125
rect 13170 36116 13176 36128
rect 13228 36116 13234 36168
rect 14366 36156 14372 36168
rect 14327 36128 14372 36156
rect 14366 36116 14372 36128
rect 14424 36116 14430 36168
rect 15470 36116 15476 36168
rect 15528 36156 15534 36168
rect 15565 36159 15623 36165
rect 15565 36156 15577 36159
rect 15528 36128 15577 36156
rect 15528 36116 15534 36128
rect 15565 36125 15577 36128
rect 15611 36125 15623 36159
rect 15565 36119 15623 36125
rect 16942 36116 16948 36168
rect 17000 36156 17006 36168
rect 17037 36159 17095 36165
rect 17037 36156 17049 36159
rect 17000 36128 17049 36156
rect 17000 36116 17006 36128
rect 17037 36125 17049 36128
rect 17083 36125 17095 36159
rect 17586 36156 17592 36168
rect 17547 36128 17592 36156
rect 17037 36119 17095 36125
rect 17586 36116 17592 36128
rect 17644 36116 17650 36168
rect 18322 36156 18328 36168
rect 18283 36128 18328 36156
rect 18322 36116 18328 36128
rect 18380 36116 18386 36168
rect 19521 36159 19579 36165
rect 19521 36125 19533 36159
rect 19567 36125 19579 36159
rect 19521 36119 19579 36125
rect 20257 36159 20315 36165
rect 20257 36125 20269 36159
rect 20303 36156 20315 36159
rect 20530 36156 20536 36168
rect 20303 36128 20536 36156
rect 20303 36125 20315 36128
rect 20257 36119 20315 36125
rect 5534 36088 5540 36100
rect 4080 36060 5540 36088
rect 5534 36048 5540 36060
rect 5592 36048 5598 36100
rect 19536 36088 19564 36119
rect 20530 36116 20536 36128
rect 20588 36116 20594 36168
rect 21913 36159 21971 36165
rect 21913 36125 21925 36159
rect 21959 36156 21971 36159
rect 22186 36156 22192 36168
rect 21959 36128 22192 36156
rect 21959 36125 21971 36128
rect 21913 36119 21971 36125
rect 22186 36116 22192 36128
rect 22244 36116 22250 36168
rect 23109 36159 23167 36165
rect 23109 36125 23121 36159
rect 23155 36156 23167 36159
rect 23290 36156 23296 36168
rect 23155 36128 23296 36156
rect 23155 36125 23167 36128
rect 23109 36119 23167 36125
rect 23290 36116 23296 36128
rect 23348 36116 23354 36168
rect 23382 36116 23388 36168
rect 23440 36156 23446 36168
rect 24397 36159 24455 36165
rect 24397 36156 24409 36159
rect 23440 36128 24409 36156
rect 23440 36116 23446 36128
rect 24397 36125 24409 36128
rect 24443 36125 24455 36159
rect 24397 36119 24455 36125
rect 25038 36116 25044 36168
rect 25096 36156 25102 36168
rect 25225 36159 25283 36165
rect 25225 36156 25237 36159
rect 25096 36128 25237 36156
rect 25096 36116 25102 36128
rect 25225 36125 25237 36128
rect 25271 36125 25283 36159
rect 26510 36156 26516 36168
rect 26471 36128 26516 36156
rect 25225 36119 25283 36125
rect 26510 36116 26516 36128
rect 26568 36116 26574 36168
rect 27614 36116 27620 36168
rect 27672 36156 27678 36168
rect 27709 36159 27767 36165
rect 27709 36156 27721 36159
rect 27672 36128 27721 36156
rect 27672 36116 27678 36128
rect 27709 36125 27721 36128
rect 27755 36125 27767 36159
rect 27709 36119 27767 36125
rect 29825 36159 29883 36165
rect 29825 36125 29837 36159
rect 29871 36156 29883 36159
rect 30098 36156 30104 36168
rect 29871 36128 30104 36156
rect 29871 36125 29883 36128
rect 29825 36119 29883 36125
rect 30098 36116 30104 36128
rect 30156 36116 30162 36168
rect 31110 36116 31116 36168
rect 31168 36156 31174 36168
rect 31297 36159 31355 36165
rect 31297 36156 31309 36159
rect 31168 36128 31309 36156
rect 31168 36116 31174 36128
rect 31297 36125 31309 36128
rect 31343 36125 31355 36159
rect 31297 36119 31355 36125
rect 33594 36116 33600 36168
rect 33652 36156 33658 36168
rect 33781 36159 33839 36165
rect 33781 36156 33793 36159
rect 33652 36128 33793 36156
rect 33652 36116 33658 36128
rect 33781 36125 33793 36128
rect 33827 36125 33839 36159
rect 33781 36119 33839 36125
rect 34698 36116 34704 36168
rect 34756 36156 34762 36168
rect 34977 36159 35035 36165
rect 34977 36156 34989 36159
rect 34756 36128 34989 36156
rect 34756 36116 34762 36128
rect 34977 36125 34989 36128
rect 35023 36125 35035 36159
rect 38010 36156 38016 36168
rect 37971 36128 38016 36156
rect 34977 36119 35035 36125
rect 38010 36116 38016 36128
rect 38068 36116 38074 36168
rect 38654 36116 38660 36168
rect 38712 36156 38718 36168
rect 38749 36159 38807 36165
rect 38749 36156 38761 36159
rect 38712 36128 38761 36156
rect 38712 36116 38718 36128
rect 38749 36125 38761 36128
rect 38795 36125 38807 36159
rect 39850 36156 39856 36168
rect 39811 36128 39856 36156
rect 38749 36119 38807 36125
rect 39850 36116 39856 36128
rect 39908 36116 39914 36168
rect 40770 36116 40776 36168
rect 40828 36156 40834 36168
rect 40957 36159 41015 36165
rect 40957 36156 40969 36159
rect 40828 36128 40969 36156
rect 40828 36116 40834 36128
rect 40957 36125 40969 36128
rect 41003 36125 41015 36159
rect 40957 36119 41015 36125
rect 43714 36116 43720 36168
rect 43772 36156 43778 36168
rect 43901 36159 43959 36165
rect 43901 36156 43913 36159
rect 43772 36128 43913 36156
rect 43772 36116 43778 36128
rect 43901 36125 43913 36128
rect 43947 36125 43959 36159
rect 43901 36119 43959 36125
rect 20438 36088 20444 36100
rect 19536 36060 20444 36088
rect 20438 36048 20444 36060
rect 20496 36048 20502 36100
rect 2958 36020 2964 36032
rect 2919 35992 2964 36020
rect 2958 35980 2964 35992
rect 3016 35980 3022 36032
rect 4062 35980 4068 36032
rect 4120 36020 4126 36032
rect 8018 36020 8024 36032
rect 4120 35992 8024 36020
rect 4120 35980 4126 35992
rect 8018 35980 8024 35992
rect 8076 35980 8082 36032
rect 10870 36020 10876 36032
rect 10831 35992 10876 36020
rect 10870 35980 10876 35992
rect 10928 35980 10934 36032
rect 19334 36020 19340 36032
rect 19295 35992 19340 36020
rect 19334 35980 19340 35992
rect 19392 35980 19398 36032
rect 29638 36020 29644 36032
rect 29599 35992 29644 36020
rect 29638 35980 29644 35992
rect 29696 35980 29702 36032
rect 30282 35980 30288 36032
rect 30340 36020 30346 36032
rect 32033 36023 32091 36029
rect 32033 36020 32045 36023
rect 30340 35992 32045 36020
rect 30340 35980 30346 35992
rect 32033 35989 32045 35992
rect 32079 36020 32091 36023
rect 32122 36020 32128 36032
rect 32079 35992 32128 36020
rect 32079 35989 32091 35992
rect 32033 35983 32091 35989
rect 32122 35980 32128 35992
rect 32180 35980 32186 36032
rect 38930 36020 38936 36032
rect 38891 35992 38936 36020
rect 38930 35980 38936 35992
rect 38988 35980 38994 36032
rect 1104 35930 44896 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 44896 35930
rect 1104 35856 44896 35878
rect 2406 35776 2412 35828
rect 2464 35816 2470 35828
rect 2961 35819 3019 35825
rect 2961 35816 2973 35819
rect 2464 35788 2973 35816
rect 2464 35776 2470 35788
rect 2961 35785 2973 35788
rect 3007 35785 3019 35819
rect 2961 35779 3019 35785
rect 3142 35776 3148 35828
rect 3200 35816 3206 35828
rect 4157 35819 4215 35825
rect 4157 35816 4169 35819
rect 3200 35788 4169 35816
rect 3200 35776 3206 35788
rect 4157 35785 4169 35788
rect 4203 35785 4215 35819
rect 4890 35816 4896 35828
rect 4851 35788 4896 35816
rect 4157 35779 4215 35785
rect 4890 35776 4896 35788
rect 4948 35776 4954 35828
rect 17126 35816 17132 35828
rect 17087 35788 17132 35816
rect 17126 35776 17132 35788
rect 17184 35776 17190 35828
rect 19058 35816 19064 35828
rect 19019 35788 19064 35816
rect 19058 35776 19064 35788
rect 19116 35776 19122 35828
rect 19426 35776 19432 35828
rect 19484 35816 19490 35828
rect 19613 35819 19671 35825
rect 19613 35816 19625 35819
rect 19484 35788 19625 35816
rect 19484 35776 19490 35788
rect 19613 35785 19625 35788
rect 19659 35785 19671 35819
rect 22094 35816 22100 35828
rect 22055 35788 22100 35816
rect 19613 35779 19671 35785
rect 22094 35776 22100 35788
rect 22152 35776 22158 35828
rect 24394 35776 24400 35828
rect 24452 35816 24458 35828
rect 24581 35819 24639 35825
rect 24581 35816 24593 35819
rect 24452 35788 24593 35816
rect 24452 35776 24458 35788
rect 24581 35785 24593 35788
rect 24627 35785 24639 35819
rect 24581 35779 24639 35785
rect 28810 35776 28816 35828
rect 28868 35816 28874 35828
rect 29638 35816 29644 35828
rect 28868 35788 29644 35816
rect 28868 35776 28874 35788
rect 29638 35776 29644 35788
rect 29696 35776 29702 35828
rect 38102 35776 38108 35828
rect 38160 35816 38166 35828
rect 38838 35816 38844 35828
rect 38160 35788 38844 35816
rect 38160 35776 38166 35788
rect 38838 35776 38844 35788
rect 38896 35776 38902 35828
rect 40126 35816 40132 35828
rect 40087 35788 40132 35816
rect 40126 35776 40132 35788
rect 40184 35776 40190 35828
rect 41325 35819 41383 35825
rect 41325 35785 41337 35819
rect 41371 35816 41383 35819
rect 41414 35816 41420 35828
rect 41371 35788 41420 35816
rect 41371 35785 41383 35788
rect 41325 35779 41383 35785
rect 41414 35776 41420 35788
rect 41472 35776 41478 35828
rect 44085 35819 44143 35825
rect 44085 35785 44097 35819
rect 44131 35816 44143 35819
rect 45738 35816 45744 35828
rect 44131 35788 45744 35816
rect 44131 35785 44143 35788
rect 44085 35779 44143 35785
rect 45738 35776 45744 35788
rect 45796 35776 45802 35828
rect 1397 35751 1455 35757
rect 1397 35717 1409 35751
rect 1443 35748 1455 35751
rect 1443 35720 2452 35748
rect 1443 35717 1455 35720
rect 1397 35711 1455 35717
rect 1673 35683 1731 35689
rect 1673 35649 1685 35683
rect 1719 35680 1731 35683
rect 1719 35652 2360 35680
rect 1719 35649 1731 35652
rect 1673 35643 1731 35649
rect 1581 35615 1639 35621
rect 1581 35581 1593 35615
rect 1627 35612 1639 35615
rect 2038 35612 2044 35624
rect 1627 35584 2044 35612
rect 1627 35581 1639 35584
rect 1581 35575 1639 35581
rect 2038 35572 2044 35584
rect 2096 35572 2102 35624
rect 2332 35553 2360 35652
rect 2424 35612 2452 35720
rect 2682 35708 2688 35760
rect 2740 35748 2746 35760
rect 3513 35751 3571 35757
rect 3513 35748 3525 35751
rect 2740 35720 3525 35748
rect 2740 35708 2746 35720
rect 3513 35717 3525 35720
rect 3559 35717 3571 35751
rect 22646 35748 22652 35760
rect 22559 35720 22652 35748
rect 3513 35711 3571 35717
rect 22646 35708 22652 35720
rect 22704 35748 22710 35760
rect 28718 35748 28724 35760
rect 22704 35720 28724 35748
rect 22704 35708 22710 35720
rect 28718 35708 28724 35720
rect 28776 35708 28782 35760
rect 38470 35708 38476 35760
rect 38528 35748 38534 35760
rect 38930 35748 38936 35760
rect 38528 35720 38936 35748
rect 38528 35708 38534 35720
rect 38930 35708 38936 35720
rect 38988 35708 38994 35760
rect 2501 35683 2559 35689
rect 2501 35649 2513 35683
rect 2547 35680 2559 35683
rect 2774 35680 2780 35692
rect 2547 35652 2780 35680
rect 2547 35649 2559 35652
rect 2501 35643 2559 35649
rect 2774 35640 2780 35652
rect 2832 35640 2838 35692
rect 33502 35680 33508 35692
rect 26206 35652 33508 35680
rect 2958 35612 2964 35624
rect 2424 35584 2964 35612
rect 2958 35572 2964 35584
rect 3016 35572 3022 35624
rect 2317 35547 2375 35553
rect 2317 35513 2329 35547
rect 2363 35513 2375 35547
rect 6454 35544 6460 35556
rect 6367 35516 6460 35544
rect 2317 35507 2375 35513
rect 6454 35504 6460 35516
rect 6512 35544 6518 35556
rect 9398 35544 9404 35556
rect 6512 35516 9404 35544
rect 6512 35504 6518 35516
rect 9398 35504 9404 35516
rect 9456 35504 9462 35556
rect 10134 35544 10140 35556
rect 10047 35516 10140 35544
rect 10134 35504 10140 35516
rect 10192 35544 10198 35556
rect 12250 35544 12256 35556
rect 10192 35516 12256 35544
rect 10192 35504 10198 35516
rect 12250 35504 12256 35516
rect 12308 35504 12314 35556
rect 25590 35504 25596 35556
rect 25648 35544 25654 35556
rect 26206 35544 26234 35652
rect 33502 35640 33508 35652
rect 33560 35640 33566 35692
rect 43622 35640 43628 35692
rect 43680 35680 43686 35692
rect 43901 35683 43959 35689
rect 43901 35680 43913 35683
rect 43680 35652 43913 35680
rect 43680 35640 43686 35652
rect 43901 35649 43913 35652
rect 43947 35649 43959 35683
rect 43901 35643 43959 35649
rect 26326 35572 26332 35624
rect 26384 35612 26390 35624
rect 30098 35612 30104 35624
rect 26384 35584 30104 35612
rect 26384 35572 26390 35584
rect 30098 35572 30104 35584
rect 30156 35572 30162 35624
rect 27614 35544 27620 35556
rect 25648 35516 26234 35544
rect 27575 35516 27620 35544
rect 25648 35504 25654 35516
rect 27614 35504 27620 35516
rect 27672 35504 27678 35556
rect 1578 35476 1584 35488
rect 1539 35448 1584 35476
rect 1578 35436 1584 35448
rect 1636 35436 1642 35488
rect 1857 35479 1915 35485
rect 1857 35445 1869 35479
rect 1903 35476 1915 35479
rect 2406 35476 2412 35488
rect 1903 35448 2412 35476
rect 1903 35445 1915 35448
rect 1857 35439 1915 35445
rect 2406 35436 2412 35448
rect 2464 35436 2470 35488
rect 8389 35479 8447 35485
rect 8389 35445 8401 35479
rect 8435 35476 8447 35479
rect 8662 35476 8668 35488
rect 8435 35448 8668 35476
rect 8435 35445 8447 35448
rect 8389 35439 8447 35445
rect 8662 35436 8668 35448
rect 8720 35436 8726 35488
rect 9490 35476 9496 35488
rect 9451 35448 9496 35476
rect 9490 35436 9496 35448
rect 9548 35436 9554 35488
rect 10962 35476 10968 35488
rect 10923 35448 10968 35476
rect 10962 35436 10968 35448
rect 11020 35436 11026 35488
rect 11974 35476 11980 35488
rect 11935 35448 11980 35476
rect 11974 35436 11980 35448
rect 12032 35436 12038 35488
rect 12618 35476 12624 35488
rect 12579 35448 12624 35476
rect 12618 35436 12624 35448
rect 12676 35436 12682 35488
rect 13170 35476 13176 35488
rect 13131 35448 13176 35476
rect 13170 35436 13176 35448
rect 13228 35436 13234 35488
rect 14458 35476 14464 35488
rect 14419 35448 14464 35476
rect 14458 35436 14464 35448
rect 14516 35436 14522 35488
rect 23198 35476 23204 35488
rect 23159 35448 23204 35476
rect 23198 35436 23204 35448
rect 23256 35436 23262 35488
rect 23658 35476 23664 35488
rect 23619 35448 23664 35476
rect 23658 35436 23664 35448
rect 23716 35436 23722 35488
rect 25222 35476 25228 35488
rect 25183 35448 25228 35476
rect 25222 35436 25228 35448
rect 25280 35436 25286 35488
rect 25961 35479 26019 35485
rect 25961 35445 25973 35479
rect 26007 35476 26019 35479
rect 26050 35476 26056 35488
rect 26007 35448 26056 35476
rect 26007 35445 26019 35448
rect 25961 35439 26019 35445
rect 26050 35436 26056 35448
rect 26108 35436 26114 35488
rect 27062 35476 27068 35488
rect 27023 35448 27068 35476
rect 27062 35436 27068 35448
rect 27120 35436 27126 35488
rect 29546 35476 29552 35488
rect 29507 35448 29552 35476
rect 29546 35436 29552 35448
rect 29604 35436 29610 35488
rect 31018 35476 31024 35488
rect 30979 35448 31024 35476
rect 31018 35436 31024 35448
rect 31076 35436 31082 35488
rect 32674 35476 32680 35488
rect 32635 35448 32680 35476
rect 32674 35436 32680 35448
rect 32732 35436 32738 35488
rect 34238 35436 34244 35488
rect 34296 35476 34302 35488
rect 34333 35479 34391 35485
rect 34333 35476 34345 35479
rect 34296 35448 34345 35476
rect 34296 35436 34302 35448
rect 34333 35445 34345 35448
rect 34379 35445 34391 35479
rect 34333 35439 34391 35445
rect 34698 35436 34704 35488
rect 34756 35476 34762 35488
rect 34885 35479 34943 35485
rect 34885 35476 34897 35479
rect 34756 35448 34897 35476
rect 34756 35436 34762 35448
rect 34885 35445 34897 35448
rect 34931 35445 34943 35479
rect 36262 35476 36268 35488
rect 36223 35448 36268 35476
rect 34885 35439 34943 35445
rect 36262 35436 36268 35448
rect 36320 35436 36326 35488
rect 37826 35476 37832 35488
rect 37787 35448 37832 35476
rect 37826 35436 37832 35448
rect 37884 35436 37890 35488
rect 38562 35476 38568 35488
rect 38523 35448 38568 35476
rect 38562 35436 38568 35448
rect 38620 35436 38626 35488
rect 39206 35476 39212 35488
rect 39167 35448 39212 35476
rect 39206 35436 39212 35448
rect 39264 35436 39270 35488
rect 40586 35476 40592 35488
rect 40547 35448 40592 35476
rect 40586 35436 40592 35448
rect 40644 35436 40650 35488
rect 42426 35476 42432 35488
rect 42387 35448 42432 35476
rect 42426 35436 42432 35448
rect 42484 35436 42490 35488
rect 43346 35476 43352 35488
rect 43307 35448 43352 35476
rect 43346 35436 43352 35448
rect 43404 35436 43410 35488
rect 1104 35386 44896 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 44896 35386
rect 1104 35312 44896 35334
rect 1578 35272 1584 35284
rect 1539 35244 1584 35272
rect 1578 35232 1584 35244
rect 1636 35232 1642 35284
rect 2038 35272 2044 35284
rect 1999 35244 2044 35272
rect 2038 35232 2044 35244
rect 2096 35232 2102 35284
rect 2222 35232 2228 35284
rect 2280 35272 2286 35284
rect 2685 35275 2743 35281
rect 2685 35272 2697 35275
rect 2280 35244 2697 35272
rect 2280 35232 2286 35244
rect 2685 35241 2697 35244
rect 2731 35241 2743 35275
rect 2685 35235 2743 35241
rect 22370 35232 22376 35284
rect 22428 35272 22434 35284
rect 26326 35272 26332 35284
rect 22428 35244 26332 35272
rect 22428 35232 22434 35244
rect 26326 35232 26332 35244
rect 26384 35232 26390 35284
rect 26421 35275 26479 35281
rect 26421 35241 26433 35275
rect 26467 35272 26479 35275
rect 26510 35272 26516 35284
rect 26467 35244 26516 35272
rect 26467 35241 26479 35244
rect 26421 35235 26479 35241
rect 26510 35232 26516 35244
rect 26568 35232 26574 35284
rect 37921 35275 37979 35281
rect 37921 35241 37933 35275
rect 37967 35272 37979 35275
rect 38010 35272 38016 35284
rect 37967 35244 38016 35272
rect 37967 35241 37979 35244
rect 37921 35235 37979 35241
rect 38010 35232 38016 35244
rect 38068 35232 38074 35284
rect 22097 35207 22155 35213
rect 22097 35173 22109 35207
rect 22143 35204 22155 35207
rect 22186 35204 22192 35216
rect 22143 35176 22192 35204
rect 22143 35173 22155 35176
rect 22097 35167 22155 35173
rect 22186 35164 22192 35176
rect 22244 35204 22250 35216
rect 26234 35204 26240 35216
rect 22244 35176 26240 35204
rect 22244 35164 22250 35176
rect 26234 35164 26240 35176
rect 26292 35164 26298 35216
rect 24210 35096 24216 35148
rect 24268 35136 24274 35148
rect 32674 35136 32680 35148
rect 24268 35108 32680 35136
rect 24268 35096 24274 35108
rect 32674 35096 32680 35108
rect 32732 35096 32738 35148
rect 1394 35068 1400 35080
rect 1355 35040 1400 35068
rect 1394 35028 1400 35040
rect 1452 35028 1458 35080
rect 2225 35071 2283 35077
rect 2225 35037 2237 35071
rect 2271 35068 2283 35071
rect 2866 35068 2872 35080
rect 2271 35040 2872 35068
rect 2271 35037 2283 35040
rect 2225 35031 2283 35037
rect 2866 35028 2872 35040
rect 2924 35028 2930 35080
rect 18414 35028 18420 35080
rect 18472 35068 18478 35080
rect 26510 35068 26516 35080
rect 18472 35040 26516 35068
rect 18472 35028 18478 35040
rect 26510 35028 26516 35040
rect 26568 35028 26574 35080
rect 4433 35003 4491 35009
rect 4433 34969 4445 35003
rect 4479 35000 4491 35003
rect 4614 35000 4620 35012
rect 4479 34972 4620 35000
rect 4479 34969 4491 34972
rect 4433 34963 4491 34969
rect 4614 34960 4620 34972
rect 4672 35000 4678 35012
rect 6362 35000 6368 35012
rect 4672 34972 6368 35000
rect 4672 34960 4678 34972
rect 6362 34960 6368 34972
rect 6420 34960 6426 35012
rect 20162 34960 20168 35012
rect 20220 35000 20226 35012
rect 26050 35000 26056 35012
rect 20220 34972 26056 35000
rect 20220 34960 20226 34972
rect 26050 34960 26056 34972
rect 26108 34960 26114 35012
rect 3878 34932 3884 34944
rect 3839 34904 3884 34932
rect 3878 34892 3884 34904
rect 3936 34892 3942 34944
rect 4985 34935 5043 34941
rect 4985 34901 4997 34935
rect 5031 34932 5043 34935
rect 5534 34932 5540 34944
rect 5031 34904 5540 34932
rect 5031 34901 5043 34904
rect 4985 34895 5043 34901
rect 5534 34892 5540 34904
rect 5592 34932 5598 34944
rect 6730 34932 6736 34944
rect 5592 34904 6736 34932
rect 5592 34892 5598 34904
rect 6730 34892 6736 34904
rect 6788 34892 6794 34944
rect 23290 34932 23296 34944
rect 23251 34904 23296 34932
rect 23290 34892 23296 34904
rect 23348 34892 23354 34944
rect 23382 34892 23388 34944
rect 23440 34932 23446 34944
rect 24397 34935 24455 34941
rect 24397 34932 24409 34935
rect 23440 34904 24409 34932
rect 23440 34892 23446 34904
rect 24397 34901 24409 34904
rect 24443 34901 24455 34935
rect 25038 34932 25044 34944
rect 24999 34904 25044 34932
rect 24397 34895 24455 34901
rect 25038 34892 25044 34904
rect 25096 34892 25102 34944
rect 30374 34932 30380 34944
rect 30335 34904 30380 34932
rect 30374 34892 30380 34904
rect 30432 34892 30438 34944
rect 31110 34932 31116 34944
rect 31071 34904 31116 34932
rect 31110 34892 31116 34904
rect 31168 34892 31174 34944
rect 33594 34932 33600 34944
rect 33555 34904 33600 34932
rect 33594 34892 33600 34904
rect 33652 34892 33658 34944
rect 34514 34892 34520 34944
rect 34572 34932 34578 34944
rect 38010 34932 38016 34944
rect 34572 34904 38016 34932
rect 34572 34892 34578 34904
rect 38010 34892 38016 34904
rect 38068 34892 38074 34944
rect 38654 34932 38660 34944
rect 38615 34904 38660 34932
rect 38654 34892 38660 34904
rect 38712 34892 38718 34944
rect 39850 34932 39856 34944
rect 39811 34904 39856 34932
rect 39850 34892 39856 34904
rect 39908 34892 39914 34944
rect 40770 34932 40776 34944
rect 40731 34904 40776 34932
rect 40770 34892 40776 34904
rect 40828 34892 40834 34944
rect 41322 34892 41328 34944
rect 41380 34932 41386 34944
rect 42981 34935 43039 34941
rect 42981 34932 42993 34935
rect 41380 34904 42993 34932
rect 41380 34892 41386 34904
rect 42981 34901 42993 34904
rect 43027 34932 43039 34935
rect 43162 34932 43168 34944
rect 43027 34904 43168 34932
rect 43027 34901 43039 34904
rect 42981 34895 43039 34901
rect 43162 34892 43168 34904
rect 43220 34892 43226 34944
rect 43530 34892 43536 34944
rect 43588 34932 43594 34944
rect 43717 34935 43775 34941
rect 43717 34932 43729 34935
rect 43588 34904 43729 34932
rect 43588 34892 43594 34904
rect 43717 34901 43729 34904
rect 43763 34901 43775 34935
rect 43717 34895 43775 34901
rect 1104 34842 44896 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 44896 34842
rect 1104 34768 44896 34790
rect 2685 34731 2743 34737
rect 2685 34697 2697 34731
rect 2731 34728 2743 34731
rect 2774 34728 2780 34740
rect 2731 34700 2780 34728
rect 2731 34697 2743 34700
rect 2685 34691 2743 34697
rect 2774 34688 2780 34700
rect 2832 34688 2838 34740
rect 25774 34688 25780 34740
rect 25832 34728 25838 34740
rect 33594 34728 33600 34740
rect 25832 34700 33600 34728
rect 25832 34688 25838 34700
rect 33594 34688 33600 34700
rect 33652 34688 33658 34740
rect 20990 34620 20996 34672
rect 21048 34660 21054 34672
rect 23658 34660 23664 34672
rect 21048 34632 23664 34660
rect 21048 34620 21054 34632
rect 23658 34620 23664 34632
rect 23716 34620 23722 34672
rect 1394 34592 1400 34604
rect 1355 34564 1400 34592
rect 1394 34552 1400 34564
rect 1452 34592 1458 34604
rect 2041 34595 2099 34601
rect 2041 34592 2053 34595
rect 1452 34564 2053 34592
rect 1452 34552 1458 34564
rect 2041 34561 2053 34564
rect 2087 34561 2099 34595
rect 3234 34592 3240 34604
rect 3147 34564 3240 34592
rect 2041 34555 2099 34561
rect 3234 34552 3240 34564
rect 3292 34592 3298 34604
rect 5166 34592 5172 34604
rect 3292 34564 5172 34592
rect 3292 34552 3298 34564
rect 5166 34552 5172 34564
rect 5224 34552 5230 34604
rect 10962 34552 10968 34604
rect 11020 34592 11026 34604
rect 12986 34592 12992 34604
rect 11020 34564 12992 34592
rect 11020 34552 11026 34564
rect 12986 34552 12992 34564
rect 13044 34552 13050 34604
rect 22830 34552 22836 34604
rect 22888 34592 22894 34604
rect 25222 34592 25228 34604
rect 22888 34564 25228 34592
rect 22888 34552 22894 34564
rect 25222 34552 25228 34564
rect 25280 34552 25286 34604
rect 3510 34484 3516 34536
rect 3568 34524 3574 34536
rect 6822 34524 6828 34536
rect 3568 34496 6828 34524
rect 3568 34484 3574 34496
rect 6822 34484 6828 34496
rect 6880 34484 6886 34536
rect 11974 34484 11980 34536
rect 12032 34524 12038 34536
rect 13262 34524 13268 34536
rect 12032 34496 13268 34524
rect 12032 34484 12038 34496
rect 13262 34484 13268 34496
rect 13320 34484 13326 34536
rect 14458 34484 14464 34536
rect 14516 34524 14522 34536
rect 15010 34524 15016 34536
rect 14516 34496 15016 34524
rect 14516 34484 14522 34496
rect 15010 34484 15016 34496
rect 15068 34484 15074 34536
rect 22738 34484 22744 34536
rect 22796 34524 22802 34536
rect 23382 34524 23388 34536
rect 22796 34496 23388 34524
rect 22796 34484 22802 34496
rect 23382 34484 23388 34496
rect 23440 34484 23446 34536
rect 26234 34484 26240 34536
rect 26292 34524 26298 34536
rect 27246 34524 27252 34536
rect 26292 34496 27252 34524
rect 26292 34484 26298 34496
rect 27246 34484 27252 34496
rect 27304 34484 27310 34536
rect 43714 34524 43720 34536
rect 43675 34496 43720 34524
rect 43714 34484 43720 34496
rect 43772 34484 43778 34536
rect 1578 34388 1584 34400
rect 1539 34360 1584 34388
rect 1578 34348 1584 34360
rect 1636 34348 1642 34400
rect 1104 34298 44896 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 44896 34298
rect 1104 34224 44896 34246
rect 1486 34184 1492 34196
rect 1447 34156 1492 34184
rect 1486 34144 1492 34156
rect 1544 34144 1550 34196
rect 2041 34187 2099 34193
rect 2041 34153 2053 34187
rect 2087 34184 2099 34187
rect 2866 34184 2872 34196
rect 2087 34156 2872 34184
rect 2087 34153 2099 34156
rect 2041 34147 2099 34153
rect 2866 34144 2872 34156
rect 2924 34144 2930 34196
rect 2498 33844 2504 33856
rect 2459 33816 2504 33844
rect 2498 33804 2504 33816
rect 2556 33804 2562 33856
rect 23198 33804 23204 33856
rect 23256 33844 23262 33856
rect 29454 33844 29460 33856
rect 23256 33816 29460 33844
rect 23256 33804 23262 33816
rect 29454 33804 29460 33816
rect 29512 33804 29518 33856
rect 43622 33804 43628 33856
rect 43680 33844 43686 33856
rect 43717 33847 43775 33853
rect 43717 33844 43729 33847
rect 43680 33816 43729 33844
rect 43680 33804 43686 33816
rect 43717 33813 43729 33816
rect 43763 33813 43775 33847
rect 43717 33807 43775 33813
rect 1104 33754 44896 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 44896 33754
rect 1104 33680 44896 33702
rect 1486 33464 1492 33516
rect 1544 33504 1550 33516
rect 1581 33507 1639 33513
rect 1581 33504 1593 33507
rect 1544 33476 1593 33504
rect 1544 33464 1550 33476
rect 1581 33473 1593 33476
rect 1627 33504 1639 33507
rect 2041 33507 2099 33513
rect 2041 33504 2053 33507
rect 1627 33476 2053 33504
rect 1627 33473 1639 33476
rect 1581 33467 1639 33473
rect 2041 33473 2053 33476
rect 2087 33473 2099 33507
rect 2041 33467 2099 33473
rect 1394 33300 1400 33312
rect 1355 33272 1400 33300
rect 1394 33260 1400 33272
rect 1452 33260 1458 33312
rect 1104 33210 44896 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 44896 33210
rect 1104 33136 44896 33158
rect 21542 33056 21548 33108
rect 21600 33096 21606 33108
rect 28534 33096 28540 33108
rect 21600 33068 28540 33096
rect 21600 33056 21606 33068
rect 28534 33056 28540 33068
rect 28592 33056 28598 33108
rect 1104 32666 44896 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 44896 32666
rect 1104 32592 44896 32614
rect 2590 32444 2596 32496
rect 2648 32484 2654 32496
rect 20070 32484 20076 32496
rect 2648 32456 20076 32484
rect 2648 32444 2654 32456
rect 20070 32444 20076 32456
rect 20128 32444 20134 32496
rect 35342 32444 35348 32496
rect 35400 32484 35406 32496
rect 43714 32484 43720 32496
rect 35400 32456 43720 32484
rect 35400 32444 35406 32456
rect 43714 32444 43720 32456
rect 43772 32444 43778 32496
rect 1397 32419 1455 32425
rect 1397 32385 1409 32419
rect 1443 32416 1455 32419
rect 1486 32416 1492 32428
rect 1443 32388 1492 32416
rect 1443 32385 1455 32388
rect 1397 32379 1455 32385
rect 1486 32376 1492 32388
rect 1544 32416 1550 32428
rect 2041 32419 2099 32425
rect 2041 32416 2053 32419
rect 1544 32388 2053 32416
rect 1544 32376 1550 32388
rect 2041 32385 2053 32388
rect 2087 32385 2099 32419
rect 2041 32379 2099 32385
rect 32766 32376 32772 32428
rect 32824 32416 32830 32428
rect 43070 32416 43076 32428
rect 32824 32388 43076 32416
rect 32824 32376 32830 32388
rect 43070 32376 43076 32388
rect 43128 32376 43134 32428
rect 1581 32215 1639 32221
rect 1581 32181 1593 32215
rect 1627 32212 1639 32215
rect 1670 32212 1676 32224
rect 1627 32184 1676 32212
rect 1627 32181 1639 32184
rect 1581 32175 1639 32181
rect 1670 32172 1676 32184
rect 1728 32172 1734 32224
rect 1104 32122 44896 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 44896 32122
rect 1104 32048 44896 32070
rect 1673 32011 1731 32017
rect 1673 31977 1685 32011
rect 1719 32008 1731 32011
rect 1762 32008 1768 32020
rect 1719 31980 1768 32008
rect 1719 31977 1731 31980
rect 1673 31971 1731 31977
rect 1762 31968 1768 31980
rect 1820 31968 1826 32020
rect 1578 31872 1584 31884
rect 1539 31844 1584 31872
rect 1578 31832 1584 31844
rect 1636 31832 1642 31884
rect 1394 31804 1400 31816
rect 1355 31776 1400 31804
rect 1394 31764 1400 31776
rect 1452 31764 1458 31816
rect 1670 31804 1676 31816
rect 1631 31776 1676 31804
rect 1670 31764 1676 31776
rect 1728 31764 1734 31816
rect 1854 31668 1860 31680
rect 1815 31640 1860 31668
rect 1854 31628 1860 31640
rect 1912 31628 1918 31680
rect 1104 31578 44896 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 44896 31578
rect 1104 31504 44896 31526
rect 1581 31467 1639 31473
rect 1581 31433 1593 31467
rect 1627 31464 1639 31467
rect 1762 31464 1768 31476
rect 1627 31436 1768 31464
rect 1627 31433 1639 31436
rect 1581 31427 1639 31433
rect 1762 31424 1768 31436
rect 1820 31424 1826 31476
rect 1394 31328 1400 31340
rect 1355 31300 1400 31328
rect 1394 31288 1400 31300
rect 1452 31328 1458 31340
rect 2041 31331 2099 31337
rect 2041 31328 2053 31331
rect 1452 31300 2053 31328
rect 1452 31288 1458 31300
rect 2041 31297 2053 31300
rect 2087 31297 2099 31331
rect 2041 31291 2099 31297
rect 1104 31034 44896 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 44896 31034
rect 1104 30960 44896 30982
rect 1104 30490 44896 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 44896 30490
rect 1104 30416 44896 30438
rect 1394 30240 1400 30252
rect 1355 30212 1400 30240
rect 1394 30200 1400 30212
rect 1452 30240 1458 30252
rect 2041 30243 2099 30249
rect 2041 30240 2053 30243
rect 1452 30212 2053 30240
rect 1452 30200 1458 30212
rect 2041 30209 2053 30212
rect 2087 30209 2099 30243
rect 2041 30203 2099 30209
rect 28994 30200 29000 30252
rect 29052 30240 29058 30252
rect 43349 30243 43407 30249
rect 43349 30240 43361 30243
rect 29052 30212 43361 30240
rect 29052 30200 29058 30212
rect 43349 30209 43361 30212
rect 43395 30240 43407 30243
rect 43901 30243 43959 30249
rect 43901 30240 43913 30243
rect 43395 30212 43913 30240
rect 43395 30209 43407 30212
rect 43349 30203 43407 30209
rect 43901 30209 43913 30212
rect 43947 30209 43959 30243
rect 43901 30203 43959 30209
rect 1578 30036 1584 30048
rect 1539 30008 1584 30036
rect 1578 29996 1584 30008
rect 1636 29996 1642 30048
rect 44082 30036 44088 30048
rect 44043 30008 44088 30036
rect 44082 29996 44088 30008
rect 44140 29996 44146 30048
rect 1104 29946 44896 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 44896 29946
rect 1104 29872 44896 29894
rect 33134 29656 33140 29708
rect 33192 29696 33198 29708
rect 41322 29696 41328 29708
rect 33192 29668 41328 29696
rect 33192 29656 33198 29668
rect 41322 29656 41328 29668
rect 41380 29656 41386 29708
rect 28074 29588 28080 29640
rect 28132 29628 28138 29640
rect 41598 29628 41604 29640
rect 28132 29600 41604 29628
rect 28132 29588 28138 29600
rect 41598 29588 41604 29600
rect 41656 29588 41662 29640
rect 1104 29402 44896 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 44896 29402
rect 1104 29328 44896 29350
rect 3510 28976 3516 29028
rect 3568 29016 3574 29028
rect 4890 29016 4896 29028
rect 3568 28988 4896 29016
rect 3568 28976 3574 28988
rect 4890 28976 4896 28988
rect 4948 28976 4954 29028
rect 1104 28858 44896 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 44896 28858
rect 1104 28784 44896 28806
rect 1486 28500 1492 28552
rect 1544 28540 1550 28552
rect 1581 28543 1639 28549
rect 1581 28540 1593 28543
rect 1544 28512 1593 28540
rect 1544 28500 1550 28512
rect 1581 28509 1593 28512
rect 1627 28540 1639 28543
rect 2041 28543 2099 28549
rect 2041 28540 2053 28543
rect 1627 28512 2053 28540
rect 1627 28509 1639 28512
rect 1581 28503 1639 28509
rect 2041 28509 2053 28512
rect 2087 28509 2099 28543
rect 2041 28503 2099 28509
rect 1394 28404 1400 28416
rect 1355 28376 1400 28404
rect 1394 28364 1400 28376
rect 1452 28364 1458 28416
rect 29270 28364 29276 28416
rect 29328 28404 29334 28416
rect 39850 28404 39856 28416
rect 29328 28376 39856 28404
rect 29328 28364 29334 28376
rect 39850 28364 39856 28376
rect 39908 28364 39914 28416
rect 1104 28314 44896 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 44896 28314
rect 1104 28240 44896 28262
rect 1394 28132 1400 28144
rect 1355 28104 1400 28132
rect 1394 28092 1400 28104
rect 1452 28092 1458 28144
rect 1670 28064 1676 28076
rect 1631 28036 1676 28064
rect 1670 28024 1676 28036
rect 1728 28024 1734 28076
rect 1578 27996 1584 28008
rect 1539 27968 1584 27996
rect 1578 27956 1584 27968
rect 1636 27956 1642 28008
rect 10870 27888 10876 27940
rect 10928 27928 10934 27940
rect 10928 27900 12434 27928
rect 10928 27888 10934 27900
rect 1578 27860 1584 27872
rect 1539 27832 1584 27860
rect 1578 27820 1584 27832
rect 1636 27820 1642 27872
rect 1857 27863 1915 27869
rect 1857 27829 1869 27863
rect 1903 27860 1915 27863
rect 2774 27860 2780 27872
rect 1903 27832 2780 27860
rect 1903 27829 1915 27832
rect 1857 27823 1915 27829
rect 2774 27820 2780 27832
rect 2832 27820 2838 27872
rect 8849 27863 8907 27869
rect 8849 27829 8861 27863
rect 8895 27860 8907 27863
rect 11054 27860 11060 27872
rect 8895 27832 11060 27860
rect 8895 27829 8907 27832
rect 8849 27823 8907 27829
rect 11054 27820 11060 27832
rect 11112 27820 11118 27872
rect 12406 27860 12434 27900
rect 31110 27860 31116 27872
rect 12406 27832 31116 27860
rect 31110 27820 31116 27832
rect 31168 27820 31174 27872
rect 1104 27770 44896 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 44896 27770
rect 1104 27696 44896 27718
rect 1581 27659 1639 27665
rect 1581 27625 1593 27659
rect 1627 27656 1639 27659
rect 1670 27656 1676 27668
rect 1627 27628 1676 27656
rect 1627 27625 1639 27628
rect 1581 27619 1639 27625
rect 1670 27616 1676 27628
rect 1728 27616 1734 27668
rect 7466 27616 7472 27668
rect 7524 27656 7530 27668
rect 29362 27656 29368 27668
rect 7524 27628 29368 27656
rect 7524 27616 7530 27628
rect 29362 27616 29368 27628
rect 29420 27616 29426 27668
rect 1854 27548 1860 27600
rect 1912 27588 1918 27600
rect 2547 27591 2605 27597
rect 2547 27588 2559 27591
rect 1912 27560 2559 27588
rect 1912 27548 1918 27560
rect 2547 27557 2559 27560
rect 2593 27557 2605 27591
rect 2682 27588 2688 27600
rect 2643 27560 2688 27588
rect 2547 27551 2605 27557
rect 2682 27548 2688 27560
rect 2740 27548 2746 27600
rect 2774 27480 2780 27532
rect 2832 27520 2838 27532
rect 2832 27492 2877 27520
rect 2832 27480 2838 27492
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27412 1458 27464
rect 2406 27452 2412 27464
rect 2367 27424 2412 27452
rect 2406 27412 2412 27424
rect 2464 27412 2470 27464
rect 3050 27316 3056 27328
rect 3011 27288 3056 27316
rect 3050 27276 3056 27288
rect 3108 27276 3114 27328
rect 8389 27319 8447 27325
rect 8389 27285 8401 27319
rect 8435 27316 8447 27319
rect 8478 27316 8484 27328
rect 8435 27288 8484 27316
rect 8435 27285 8447 27288
rect 8389 27279 8447 27285
rect 8478 27276 8484 27288
rect 8536 27276 8542 27328
rect 9030 27316 9036 27328
rect 8991 27288 9036 27316
rect 9030 27276 9036 27288
rect 9088 27276 9094 27328
rect 9582 27316 9588 27328
rect 9543 27288 9588 27316
rect 9582 27276 9588 27288
rect 9640 27276 9646 27328
rect 10962 27276 10968 27328
rect 11020 27316 11026 27328
rect 11149 27319 11207 27325
rect 11149 27316 11161 27319
rect 11020 27288 11161 27316
rect 11020 27276 11026 27288
rect 11149 27285 11161 27288
rect 11195 27316 11207 27319
rect 26602 27316 26608 27328
rect 11195 27288 26608 27316
rect 11195 27285 11207 27288
rect 11149 27279 11207 27285
rect 26602 27276 26608 27288
rect 26660 27276 26666 27328
rect 1104 27226 44896 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 44896 27226
rect 1104 27152 44896 27174
rect 1394 27112 1400 27124
rect 1355 27084 1400 27112
rect 1394 27072 1400 27084
rect 1452 27072 1458 27124
rect 8018 27112 8024 27124
rect 7979 27084 8024 27112
rect 8018 27072 8024 27084
rect 8076 27072 8082 27124
rect 9309 27115 9367 27121
rect 9309 27081 9321 27115
rect 9355 27112 9367 27115
rect 9582 27112 9588 27124
rect 9355 27084 9588 27112
rect 9355 27081 9367 27084
rect 9309 27075 9367 27081
rect 9582 27072 9588 27084
rect 9640 27072 9646 27124
rect 9030 27004 9036 27056
rect 9088 27044 9094 27056
rect 17402 27044 17408 27056
rect 9088 27016 17408 27044
rect 9088 27004 9094 27016
rect 17402 27004 17408 27016
rect 17460 27004 17466 27056
rect 4062 26936 4068 26988
rect 4120 26976 4126 26988
rect 11330 26976 11336 26988
rect 4120 26948 11336 26976
rect 4120 26936 4126 26948
rect 11330 26936 11336 26948
rect 11388 26936 11394 26988
rect 10502 26868 10508 26920
rect 10560 26908 10566 26920
rect 25222 26908 25228 26920
rect 10560 26880 25228 26908
rect 10560 26868 10566 26880
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 6638 26800 6644 26852
rect 6696 26840 6702 26852
rect 11514 26840 11520 26852
rect 6696 26812 11520 26840
rect 6696 26800 6702 26812
rect 11514 26800 11520 26812
rect 11572 26800 11578 26852
rect 11698 26800 11704 26852
rect 11756 26840 11762 26852
rect 12621 26843 12679 26849
rect 12621 26840 12633 26843
rect 11756 26812 12633 26840
rect 11756 26800 11762 26812
rect 12621 26809 12633 26812
rect 12667 26809 12679 26843
rect 12621 26803 12679 26809
rect 1854 26732 1860 26784
rect 1912 26772 1918 26784
rect 1949 26775 2007 26781
rect 1949 26772 1961 26775
rect 1912 26744 1961 26772
rect 1912 26732 1918 26744
rect 1949 26741 1961 26744
rect 1995 26741 2007 26775
rect 1949 26735 2007 26741
rect 2222 26732 2228 26784
rect 2280 26772 2286 26784
rect 2501 26775 2559 26781
rect 2501 26772 2513 26775
rect 2280 26744 2513 26772
rect 2280 26732 2286 26744
rect 2501 26741 2513 26744
rect 2547 26741 2559 26775
rect 8570 26772 8576 26784
rect 8531 26744 8576 26772
rect 2501 26735 2559 26741
rect 8570 26732 8576 26744
rect 8628 26732 8634 26784
rect 9861 26775 9919 26781
rect 9861 26741 9873 26775
rect 9907 26772 9919 26775
rect 10042 26772 10048 26784
rect 9907 26744 10048 26772
rect 9907 26741 9919 26744
rect 9861 26735 9919 26741
rect 10042 26732 10048 26744
rect 10100 26732 10106 26784
rect 10226 26732 10232 26784
rect 10284 26772 10290 26784
rect 10321 26775 10379 26781
rect 10321 26772 10333 26775
rect 10284 26744 10333 26772
rect 10284 26732 10290 26744
rect 10321 26741 10333 26744
rect 10367 26772 10379 26775
rect 10870 26772 10876 26784
rect 10367 26744 10876 26772
rect 10367 26741 10379 26744
rect 10321 26735 10379 26741
rect 10870 26732 10876 26744
rect 10928 26732 10934 26784
rect 12161 26775 12219 26781
rect 12161 26741 12173 26775
rect 12207 26772 12219 26775
rect 16298 26772 16304 26784
rect 12207 26744 16304 26772
rect 12207 26741 12219 26744
rect 12161 26735 12219 26741
rect 16298 26732 16304 26744
rect 16356 26732 16362 26784
rect 1104 26682 44896 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 44896 26682
rect 1104 26608 44896 26630
rect 1578 26568 1584 26580
rect 1539 26540 1584 26568
rect 1578 26528 1584 26540
rect 1636 26528 1642 26580
rect 2406 26528 2412 26580
rect 2464 26568 2470 26580
rect 6638 26568 6644 26580
rect 2464 26540 6644 26568
rect 2464 26528 2470 26540
rect 6638 26528 6644 26540
rect 6696 26528 6702 26580
rect 6822 26528 6828 26580
rect 6880 26568 6886 26580
rect 7009 26571 7067 26577
rect 7009 26568 7021 26571
rect 6880 26540 7021 26568
rect 6880 26528 6886 26540
rect 7009 26537 7021 26540
rect 7055 26537 7067 26571
rect 10410 26568 10416 26580
rect 7009 26531 7067 26537
rect 7116 26540 9628 26568
rect 10371 26540 10416 26568
rect 6086 26460 6092 26512
rect 6144 26500 6150 26512
rect 7116 26500 7144 26540
rect 9490 26500 9496 26512
rect 6144 26472 7144 26500
rect 9451 26472 9496 26500
rect 6144 26460 6150 26472
rect 9490 26460 9496 26472
rect 9548 26460 9554 26512
rect 9600 26500 9628 26540
rect 10410 26528 10416 26540
rect 10468 26528 10474 26580
rect 16482 26568 16488 26580
rect 12452 26540 16488 26568
rect 9600 26472 10916 26500
rect 10888 26432 10916 26472
rect 11514 26460 11520 26512
rect 11572 26500 11578 26512
rect 12452 26500 12480 26540
rect 16482 26528 16488 26540
rect 16540 26528 16546 26580
rect 12618 26500 12624 26512
rect 11572 26472 12480 26500
rect 12579 26472 12624 26500
rect 11572 26460 11578 26472
rect 12618 26460 12624 26472
rect 12676 26460 12682 26512
rect 13354 26460 13360 26512
rect 13412 26500 13418 26512
rect 31570 26500 31576 26512
rect 13412 26472 31576 26500
rect 13412 26460 13418 26472
rect 31570 26460 31576 26472
rect 31628 26460 31634 26512
rect 30190 26432 30196 26444
rect 10888 26404 30196 26432
rect 30190 26392 30196 26404
rect 30248 26392 30254 26444
rect 1394 26364 1400 26376
rect 1355 26336 1400 26364
rect 1394 26324 1400 26336
rect 1452 26364 1458 26376
rect 2041 26367 2099 26373
rect 2041 26364 2053 26367
rect 1452 26336 2053 26364
rect 1452 26324 1458 26336
rect 2041 26333 2053 26336
rect 2087 26333 2099 26367
rect 2041 26327 2099 26333
rect 2130 26324 2136 26376
rect 2188 26364 2194 26376
rect 3145 26367 3203 26373
rect 3145 26364 3157 26367
rect 2188 26336 3157 26364
rect 2188 26324 2194 26336
rect 3145 26333 3157 26336
rect 3191 26333 3203 26367
rect 3145 26327 3203 26333
rect 9582 26324 9588 26376
rect 9640 26364 9646 26376
rect 11977 26367 12035 26373
rect 11977 26364 11989 26367
rect 9640 26336 11989 26364
rect 9640 26324 9646 26336
rect 11977 26333 11989 26336
rect 12023 26364 12035 26367
rect 12066 26364 12072 26376
rect 12023 26336 12072 26364
rect 12023 26333 12035 26336
rect 11977 26327 12035 26333
rect 12066 26324 12072 26336
rect 12124 26324 12130 26376
rect 19334 26364 19340 26376
rect 12406 26336 19340 26364
rect 3786 26296 3792 26308
rect 3747 26268 3792 26296
rect 3786 26256 3792 26268
rect 3844 26256 3850 26308
rect 7653 26299 7711 26305
rect 7653 26265 7665 26299
rect 7699 26296 7711 26299
rect 7699 26268 8340 26296
rect 7699 26265 7711 26268
rect 7653 26259 7711 26265
rect 8312 26240 8340 26268
rect 8754 26256 8760 26308
rect 8812 26296 8818 26308
rect 9033 26299 9091 26305
rect 9033 26296 9045 26299
rect 8812 26268 9045 26296
rect 8812 26256 8818 26268
rect 9033 26265 9045 26268
rect 9079 26296 9091 26299
rect 10502 26296 10508 26308
rect 9079 26268 10508 26296
rect 9079 26265 9091 26268
rect 9033 26259 9091 26265
rect 10502 26256 10508 26268
rect 10560 26256 10566 26308
rect 10594 26256 10600 26308
rect 10652 26296 10658 26308
rect 10873 26299 10931 26305
rect 10873 26296 10885 26299
rect 10652 26268 10885 26296
rect 10652 26256 10658 26268
rect 10873 26265 10885 26268
rect 10919 26265 10931 26299
rect 11517 26299 11575 26305
rect 11517 26296 11529 26299
rect 10873 26259 10931 26265
rect 10980 26268 11529 26296
rect 2498 26188 2504 26240
rect 2556 26228 2562 26240
rect 2593 26231 2651 26237
rect 2593 26228 2605 26231
rect 2556 26200 2605 26228
rect 2556 26188 2562 26200
rect 2593 26197 2605 26200
rect 2639 26197 2651 26231
rect 8294 26228 8300 26240
rect 8255 26200 8300 26228
rect 2593 26191 2651 26197
rect 8294 26188 8300 26200
rect 8352 26188 8358 26240
rect 9858 26188 9864 26240
rect 9916 26228 9922 26240
rect 10980 26228 11008 26268
rect 11517 26265 11529 26268
rect 11563 26296 11575 26299
rect 12406 26296 12434 26336
rect 19334 26324 19340 26336
rect 19392 26324 19398 26376
rect 33226 26364 33232 26376
rect 22066 26336 33232 26364
rect 13078 26296 13084 26308
rect 11563 26268 12434 26296
rect 13039 26268 13084 26296
rect 11563 26265 11575 26268
rect 11517 26259 11575 26265
rect 13078 26256 13084 26268
rect 13136 26256 13142 26308
rect 16482 26256 16488 26308
rect 16540 26296 16546 26308
rect 22066 26296 22094 26336
rect 33226 26324 33232 26336
rect 33284 26324 33290 26376
rect 16540 26268 22094 26296
rect 16540 26256 16546 26268
rect 9916 26200 11008 26228
rect 9916 26188 9922 26200
rect 1104 26138 44896 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 44896 26138
rect 1104 26064 44896 26086
rect 6914 26024 6920 26036
rect 6875 25996 6920 26024
rect 6914 25984 6920 25996
rect 6972 25984 6978 26036
rect 10318 25984 10324 26036
rect 10376 26024 10382 26036
rect 10413 26027 10471 26033
rect 10413 26024 10425 26027
rect 10376 25996 10425 26024
rect 10376 25984 10382 25996
rect 10413 25993 10425 25996
rect 10459 25993 10471 26027
rect 12066 26024 12072 26036
rect 12027 25996 12072 26024
rect 10413 25987 10471 25993
rect 12066 25984 12072 25996
rect 12124 25984 12130 26036
rect 7650 25848 7656 25900
rect 7708 25888 7714 25900
rect 10042 25888 10048 25900
rect 7708 25860 10048 25888
rect 7708 25848 7714 25860
rect 10042 25848 10048 25860
rect 10100 25848 10106 25900
rect 1394 25780 1400 25832
rect 1452 25820 1458 25832
rect 1949 25823 2007 25829
rect 1949 25820 1961 25823
rect 1452 25792 1961 25820
rect 1452 25780 1458 25792
rect 1949 25789 1961 25792
rect 1995 25789 2007 25823
rect 1949 25783 2007 25789
rect 8297 25823 8355 25829
rect 8297 25789 8309 25823
rect 8343 25820 8355 25823
rect 8570 25820 8576 25832
rect 8343 25792 8576 25820
rect 8343 25789 8355 25792
rect 8297 25783 8355 25789
rect 8570 25780 8576 25792
rect 8628 25780 8634 25832
rect 10134 25820 10140 25832
rect 9646 25792 10140 25820
rect 5813 25755 5871 25761
rect 5813 25721 5825 25755
rect 5859 25752 5871 25755
rect 9646 25752 9674 25792
rect 10134 25780 10140 25792
rect 10192 25820 10198 25832
rect 13449 25823 13507 25829
rect 13449 25820 13461 25823
rect 10192 25792 13461 25820
rect 10192 25780 10198 25792
rect 13449 25789 13461 25792
rect 13495 25789 13507 25823
rect 13449 25783 13507 25789
rect 5859 25724 9674 25752
rect 5859 25721 5871 25724
rect 5813 25715 5871 25721
rect 12066 25712 12072 25764
rect 12124 25752 12130 25764
rect 25130 25752 25136 25764
rect 12124 25724 25136 25752
rect 12124 25712 12130 25724
rect 25130 25712 25136 25724
rect 25188 25712 25194 25764
rect 1486 25684 1492 25696
rect 1447 25656 1492 25684
rect 1486 25644 1492 25656
rect 1544 25644 1550 25696
rect 2314 25644 2320 25696
rect 2372 25684 2378 25696
rect 2866 25684 2872 25696
rect 2372 25656 2872 25684
rect 2372 25644 2378 25656
rect 2866 25644 2872 25656
rect 2924 25644 2930 25696
rect 2958 25644 2964 25696
rect 3016 25684 3022 25696
rect 3234 25684 3240 25696
rect 3016 25656 3240 25684
rect 3016 25644 3022 25656
rect 3234 25644 3240 25656
rect 3292 25684 3298 25696
rect 3421 25687 3479 25693
rect 3421 25684 3433 25687
rect 3292 25656 3433 25684
rect 3292 25644 3298 25656
rect 3421 25653 3433 25656
rect 3467 25653 3479 25687
rect 3421 25647 3479 25653
rect 3510 25644 3516 25696
rect 3568 25684 3574 25696
rect 3973 25687 4031 25693
rect 3973 25684 3985 25687
rect 3568 25656 3985 25684
rect 3568 25644 3574 25656
rect 3973 25653 3985 25656
rect 4019 25653 4031 25687
rect 3973 25647 4031 25653
rect 5718 25644 5724 25696
rect 5776 25684 5782 25696
rect 7650 25684 7656 25696
rect 5776 25656 7656 25684
rect 5776 25644 5782 25656
rect 7650 25644 7656 25656
rect 7708 25644 7714 25696
rect 8386 25644 8392 25696
rect 8444 25684 8450 25696
rect 8757 25687 8815 25693
rect 8757 25684 8769 25687
rect 8444 25656 8769 25684
rect 8444 25644 8450 25656
rect 8757 25653 8769 25656
rect 8803 25653 8815 25687
rect 8757 25647 8815 25653
rect 9214 25644 9220 25696
rect 9272 25684 9278 25696
rect 9309 25687 9367 25693
rect 9309 25684 9321 25687
rect 9272 25656 9321 25684
rect 9272 25644 9278 25656
rect 9309 25653 9321 25656
rect 9355 25653 9367 25687
rect 9309 25647 9367 25653
rect 9766 25644 9772 25696
rect 9824 25684 9830 25696
rect 9861 25687 9919 25693
rect 9861 25684 9873 25687
rect 9824 25656 9873 25684
rect 9824 25644 9830 25656
rect 9861 25653 9873 25656
rect 9907 25653 9919 25687
rect 11514 25684 11520 25696
rect 11475 25656 11520 25684
rect 9861 25647 9919 25653
rect 11514 25644 11520 25656
rect 11572 25644 11578 25696
rect 12989 25687 13047 25693
rect 12989 25653 13001 25687
rect 13035 25684 13047 25687
rect 13078 25684 13084 25696
rect 13035 25656 13084 25684
rect 13035 25653 13047 25656
rect 12989 25647 13047 25653
rect 13078 25644 13084 25656
rect 13136 25644 13142 25696
rect 14090 25684 14096 25696
rect 14051 25656 14096 25684
rect 14090 25644 14096 25656
rect 14148 25644 14154 25696
rect 1104 25594 44896 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 44896 25594
rect 1104 25520 44896 25542
rect 4433 25483 4491 25489
rect 4433 25449 4445 25483
rect 4479 25480 4491 25483
rect 4982 25480 4988 25492
rect 4479 25452 4988 25480
rect 4479 25449 4491 25452
rect 4433 25443 4491 25449
rect 4982 25440 4988 25452
rect 5040 25440 5046 25492
rect 5074 25440 5080 25492
rect 5132 25480 5138 25492
rect 5442 25480 5448 25492
rect 5132 25452 5448 25480
rect 5132 25440 5138 25452
rect 5442 25440 5448 25452
rect 5500 25480 5506 25492
rect 5537 25483 5595 25489
rect 5537 25480 5549 25483
rect 5500 25452 5549 25480
rect 5500 25440 5506 25452
rect 5537 25449 5549 25452
rect 5583 25449 5595 25483
rect 7558 25480 7564 25492
rect 5537 25443 5595 25449
rect 6104 25452 7564 25480
rect 750 25372 756 25424
rect 808 25412 814 25424
rect 3142 25412 3148 25424
rect 808 25384 3148 25412
rect 808 25372 814 25384
rect 3142 25372 3148 25384
rect 3200 25372 3206 25424
rect 3602 25372 3608 25424
rect 3660 25412 3666 25424
rect 6104 25421 6132 25452
rect 7558 25440 7564 25452
rect 7616 25440 7622 25492
rect 9030 25440 9036 25492
rect 9088 25480 9094 25492
rect 9125 25483 9183 25489
rect 9125 25480 9137 25483
rect 9088 25452 9137 25480
rect 9088 25440 9094 25452
rect 9125 25449 9137 25452
rect 9171 25480 9183 25483
rect 9582 25480 9588 25492
rect 9171 25452 9588 25480
rect 9171 25449 9183 25452
rect 9125 25443 9183 25449
rect 9582 25440 9588 25452
rect 9640 25440 9646 25492
rect 10321 25483 10379 25489
rect 10321 25449 10333 25483
rect 10367 25480 10379 25483
rect 10502 25480 10508 25492
rect 10367 25452 10508 25480
rect 10367 25449 10379 25452
rect 10321 25443 10379 25449
rect 10502 25440 10508 25452
rect 10560 25440 10566 25492
rect 11146 25480 11152 25492
rect 11107 25452 11152 25480
rect 11146 25440 11152 25452
rect 11204 25440 11210 25492
rect 11422 25440 11428 25492
rect 11480 25480 11486 25492
rect 11701 25483 11759 25489
rect 11701 25480 11713 25483
rect 11480 25452 11713 25480
rect 11480 25440 11486 25452
rect 11701 25449 11713 25452
rect 11747 25480 11759 25483
rect 12526 25480 12532 25492
rect 11747 25452 12532 25480
rect 11747 25449 11759 25452
rect 11701 25443 11759 25449
rect 12526 25440 12532 25452
rect 12584 25440 12590 25492
rect 6089 25415 6147 25421
rect 6089 25412 6101 25415
rect 3660 25384 6101 25412
rect 3660 25372 3666 25384
rect 6089 25381 6101 25384
rect 6135 25381 6147 25415
rect 6089 25375 6147 25381
rect 9769 25415 9827 25421
rect 9769 25381 9781 25415
rect 9815 25412 9827 25415
rect 11238 25412 11244 25424
rect 9815 25384 11244 25412
rect 9815 25381 9827 25384
rect 9769 25375 9827 25381
rect 11238 25372 11244 25384
rect 11296 25372 11302 25424
rect 12618 25372 12624 25424
rect 12676 25412 12682 25424
rect 18874 25412 18880 25424
rect 12676 25384 18880 25412
rect 12676 25372 12682 25384
rect 18874 25372 18880 25384
rect 18932 25372 18938 25424
rect 1210 25304 1216 25356
rect 1268 25344 1274 25356
rect 1268 25316 9628 25344
rect 1268 25304 1274 25316
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 1946 25236 1952 25288
rect 2004 25276 2010 25288
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 2004 25248 3801 25276
rect 2004 25236 2010 25248
rect 3789 25245 3801 25248
rect 3835 25276 3847 25279
rect 5718 25276 5724 25288
rect 3835 25248 5724 25276
rect 3835 25245 3847 25248
rect 3789 25239 3847 25245
rect 5718 25236 5724 25248
rect 5776 25236 5782 25288
rect 5902 25236 5908 25288
rect 5960 25276 5966 25288
rect 7929 25279 7987 25285
rect 7929 25276 7941 25279
rect 5960 25248 7941 25276
rect 5960 25236 5966 25248
rect 7929 25245 7941 25248
rect 7975 25245 7987 25279
rect 7929 25239 7987 25245
rect 8294 25236 8300 25288
rect 8352 25276 8358 25288
rect 9600 25285 9628 25316
rect 12434 25304 12440 25356
rect 12492 25344 12498 25356
rect 12805 25347 12863 25353
rect 12805 25344 12817 25347
rect 12492 25316 12817 25344
rect 12492 25304 12498 25316
rect 12805 25313 12817 25316
rect 12851 25344 12863 25347
rect 13357 25347 13415 25353
rect 13357 25344 13369 25347
rect 12851 25316 13369 25344
rect 12851 25313 12863 25316
rect 12805 25307 12863 25313
rect 13357 25313 13369 25316
rect 13403 25344 13415 25347
rect 31754 25344 31760 25356
rect 13403 25316 31760 25344
rect 13403 25313 13415 25316
rect 13357 25307 13415 25313
rect 31754 25304 31760 25316
rect 31812 25304 31818 25356
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8352 25248 8953 25276
rect 8352 25236 8358 25248
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 9585 25279 9643 25285
rect 9585 25245 9597 25279
rect 9631 25245 9643 25279
rect 9585 25239 9643 25245
rect 11330 25236 11336 25288
rect 11388 25276 11394 25288
rect 11882 25276 11888 25288
rect 11388 25248 11888 25276
rect 11388 25236 11394 25248
rect 11882 25236 11888 25248
rect 11940 25276 11946 25288
rect 14093 25279 14151 25285
rect 14093 25276 14105 25279
rect 11940 25248 14105 25276
rect 11940 25236 11946 25248
rect 14093 25245 14105 25248
rect 14139 25245 14151 25279
rect 14093 25239 14151 25245
rect 14458 25236 14464 25288
rect 14516 25276 14522 25288
rect 23842 25276 23848 25288
rect 14516 25248 23848 25276
rect 14516 25236 14522 25248
rect 23842 25236 23848 25248
rect 23900 25236 23906 25288
rect 2501 25211 2559 25217
rect 2501 25177 2513 25211
rect 2547 25208 2559 25211
rect 8478 25208 8484 25220
rect 2547 25180 8484 25208
rect 2547 25177 2559 25180
rect 2501 25171 2559 25177
rect 8478 25168 8484 25180
rect 8536 25168 8542 25220
rect 18874 25168 18880 25220
rect 18932 25208 18938 25220
rect 23014 25208 23020 25220
rect 18932 25180 23020 25208
rect 18932 25168 18938 25180
rect 23014 25168 23020 25180
rect 23072 25168 23078 25220
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 3053 25143 3111 25149
rect 3053 25109 3065 25143
rect 3099 25140 3111 25143
rect 3142 25140 3148 25152
rect 3099 25112 3148 25140
rect 3099 25109 3111 25112
rect 3053 25103 3111 25109
rect 3142 25100 3148 25112
rect 3200 25100 3206 25152
rect 3878 25100 3884 25152
rect 3936 25140 3942 25152
rect 4893 25143 4951 25149
rect 4893 25140 4905 25143
rect 3936 25112 4905 25140
rect 3936 25100 3942 25112
rect 4893 25109 4905 25112
rect 4939 25109 4951 25143
rect 6638 25140 6644 25152
rect 6599 25112 6644 25140
rect 4893 25103 4951 25109
rect 6638 25100 6644 25112
rect 6696 25100 6702 25152
rect 7190 25140 7196 25152
rect 7151 25112 7196 25140
rect 7190 25100 7196 25112
rect 7248 25100 7254 25152
rect 7282 25100 7288 25152
rect 7340 25140 7346 25152
rect 7745 25143 7803 25149
rect 7745 25140 7757 25143
rect 7340 25112 7757 25140
rect 7340 25100 7346 25112
rect 7745 25109 7757 25112
rect 7791 25109 7803 25143
rect 7745 25103 7803 25109
rect 12253 25143 12311 25149
rect 12253 25109 12265 25143
rect 12299 25140 12311 25143
rect 12342 25140 12348 25152
rect 12299 25112 12348 25140
rect 12299 25109 12311 25112
rect 12253 25103 12311 25109
rect 12342 25100 12348 25112
rect 12400 25100 12406 25152
rect 14737 25143 14795 25149
rect 14737 25109 14749 25143
rect 14783 25140 14795 25143
rect 16758 25140 16764 25152
rect 14783 25112 16764 25140
rect 14783 25109 14795 25112
rect 14737 25103 14795 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 1104 25050 44896 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 44896 25050
rect 1104 24976 44896 24998
rect 3142 24896 3148 24948
rect 3200 24936 3206 24948
rect 9858 24936 9864 24948
rect 3200 24908 9864 24936
rect 3200 24896 3206 24908
rect 9858 24896 9864 24908
rect 9916 24896 9922 24948
rect 11054 24896 11060 24948
rect 11112 24936 11118 24948
rect 15746 24936 15752 24948
rect 11112 24908 15752 24936
rect 11112 24896 11118 24908
rect 15746 24896 15752 24908
rect 15804 24936 15810 24948
rect 18690 24936 18696 24948
rect 15804 24908 18696 24936
rect 15804 24896 15810 24908
rect 18690 24896 18696 24908
rect 18748 24896 18754 24948
rect 18782 24896 18788 24948
rect 18840 24936 18846 24948
rect 26326 24936 26332 24948
rect 18840 24908 26332 24936
rect 18840 24896 18846 24908
rect 26326 24896 26332 24908
rect 26384 24896 26390 24948
rect 9217 24871 9275 24877
rect 9217 24837 9229 24871
rect 9263 24868 9275 24871
rect 10042 24868 10048 24880
rect 9263 24840 10048 24868
rect 9263 24837 9275 24840
rect 9217 24831 9275 24837
rect 10042 24828 10048 24840
rect 10100 24828 10106 24880
rect 12342 24828 12348 24880
rect 12400 24868 12406 24880
rect 12713 24871 12771 24877
rect 12713 24868 12725 24871
rect 12400 24840 12725 24868
rect 12400 24828 12406 24840
rect 12713 24837 12725 24840
rect 12759 24868 12771 24871
rect 17678 24868 17684 24880
rect 12759 24840 17684 24868
rect 12759 24837 12771 24840
rect 12713 24831 12771 24837
rect 17678 24828 17684 24840
rect 17736 24828 17742 24880
rect 18046 24828 18052 24880
rect 18104 24868 18110 24880
rect 33502 24868 33508 24880
rect 18104 24840 33508 24868
rect 18104 24828 18110 24840
rect 33502 24828 33508 24840
rect 33560 24828 33566 24880
rect 3142 24760 3148 24812
rect 3200 24800 3206 24812
rect 3418 24800 3424 24812
rect 3200 24772 3424 24800
rect 3200 24760 3206 24772
rect 3418 24760 3424 24772
rect 3476 24800 3482 24812
rect 3513 24803 3571 24809
rect 3513 24800 3525 24803
rect 3476 24772 3525 24800
rect 3476 24760 3482 24772
rect 3513 24769 3525 24772
rect 3559 24769 3571 24803
rect 3513 24763 3571 24769
rect 5258 24760 5264 24812
rect 5316 24800 5322 24812
rect 7285 24803 7343 24809
rect 7285 24800 7297 24803
rect 5316 24772 7297 24800
rect 5316 24760 5322 24772
rect 7285 24769 7297 24772
rect 7331 24769 7343 24803
rect 7285 24763 7343 24769
rect 7929 24803 7987 24809
rect 7929 24769 7941 24803
rect 7975 24800 7987 24803
rect 8294 24800 8300 24812
rect 7975 24772 8300 24800
rect 7975 24769 7987 24772
rect 7929 24763 7987 24769
rect 1857 24735 1915 24741
rect 1857 24701 1869 24735
rect 1903 24732 1915 24735
rect 2774 24732 2780 24744
rect 1903 24704 2780 24732
rect 1903 24701 1915 24704
rect 1857 24695 1915 24701
rect 2774 24692 2780 24704
rect 2832 24732 2838 24744
rect 3050 24732 3056 24744
rect 2832 24704 3056 24732
rect 2832 24692 2838 24704
rect 3050 24692 3056 24704
rect 3108 24692 3114 24744
rect 7944 24732 7972 24763
rect 8294 24760 8300 24772
rect 8352 24760 8358 24812
rect 8570 24800 8576 24812
rect 8531 24772 8576 24800
rect 8570 24760 8576 24772
rect 8628 24760 8634 24812
rect 9766 24800 9772 24812
rect 9727 24772 9772 24800
rect 9766 24760 9772 24772
rect 9824 24760 9830 24812
rect 10594 24800 10600 24812
rect 10555 24772 10600 24800
rect 10594 24760 10600 24772
rect 10652 24760 10658 24812
rect 14090 24760 14096 24812
rect 14148 24800 14154 24812
rect 15838 24800 15844 24812
rect 14148 24772 15844 24800
rect 14148 24760 14154 24772
rect 15838 24760 15844 24772
rect 15896 24800 15902 24812
rect 22922 24800 22928 24812
rect 15896 24772 22928 24800
rect 15896 24760 15902 24772
rect 22922 24760 22928 24772
rect 22980 24760 22986 24812
rect 5184 24704 7972 24732
rect 2038 24624 2044 24676
rect 2096 24664 2102 24676
rect 2961 24667 3019 24673
rect 2961 24664 2973 24667
rect 2096 24636 2973 24664
rect 2096 24624 2102 24636
rect 2961 24633 2973 24636
rect 3007 24633 3019 24667
rect 4154 24664 4160 24676
rect 4115 24636 4160 24664
rect 2961 24627 3019 24633
rect 4154 24624 4160 24636
rect 4212 24624 4218 24676
rect 2406 24596 2412 24608
rect 2367 24568 2412 24596
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 4706 24596 4712 24608
rect 4667 24568 4712 24596
rect 4706 24556 4712 24568
rect 4764 24556 4770 24608
rect 5074 24556 5080 24608
rect 5132 24596 5138 24608
rect 5184 24605 5212 24704
rect 8386 24692 8392 24744
rect 8444 24732 8450 24744
rect 14921 24735 14979 24741
rect 8444 24704 10548 24732
rect 8444 24692 8450 24704
rect 7466 24624 7472 24676
rect 7524 24664 7530 24676
rect 10413 24667 10471 24673
rect 10413 24664 10425 24667
rect 7524 24636 10425 24664
rect 7524 24624 7530 24636
rect 10413 24633 10425 24636
rect 10459 24633 10471 24667
rect 10520 24664 10548 24704
rect 14921 24701 14933 24735
rect 14967 24732 14979 24735
rect 15473 24735 15531 24741
rect 15473 24732 15485 24735
rect 14967 24704 15485 24732
rect 14967 24701 14979 24704
rect 14921 24695 14979 24701
rect 15473 24701 15485 24704
rect 15519 24732 15531 24735
rect 16390 24732 16396 24744
rect 15519 24704 16396 24732
rect 15519 24701 15531 24704
rect 15473 24695 15531 24701
rect 16390 24692 16396 24704
rect 16448 24732 16454 24744
rect 26970 24732 26976 24744
rect 16448 24704 26976 24732
rect 16448 24692 16454 24704
rect 26970 24692 26976 24704
rect 27028 24692 27034 24744
rect 11517 24667 11575 24673
rect 11517 24664 11529 24667
rect 10520 24636 11529 24664
rect 10413 24627 10471 24633
rect 11517 24633 11529 24636
rect 11563 24664 11575 24667
rect 11606 24664 11612 24676
rect 11563 24636 11612 24664
rect 11563 24633 11575 24636
rect 11517 24627 11575 24633
rect 11606 24624 11612 24636
rect 11664 24624 11670 24676
rect 16761 24667 16819 24673
rect 16761 24633 16773 24667
rect 16807 24664 16819 24667
rect 17310 24664 17316 24676
rect 16807 24636 17316 24664
rect 16807 24633 16819 24636
rect 16761 24627 16819 24633
rect 17310 24624 17316 24636
rect 17368 24624 17374 24676
rect 5169 24599 5227 24605
rect 5169 24596 5181 24599
rect 5132 24568 5181 24596
rect 5132 24556 5138 24568
rect 5169 24565 5181 24568
rect 5215 24565 5227 24599
rect 5810 24596 5816 24608
rect 5771 24568 5816 24596
rect 5169 24559 5227 24565
rect 5810 24556 5816 24568
rect 5868 24556 5874 24608
rect 6270 24556 6276 24608
rect 6328 24596 6334 24608
rect 6549 24599 6607 24605
rect 6549 24596 6561 24599
rect 6328 24568 6561 24596
rect 6328 24556 6334 24568
rect 6549 24565 6561 24568
rect 6595 24565 6607 24599
rect 7098 24596 7104 24608
rect 7059 24568 7104 24596
rect 6549 24559 6607 24565
rect 7098 24556 7104 24568
rect 7156 24556 7162 24608
rect 7745 24599 7803 24605
rect 7745 24565 7757 24599
rect 7791 24596 7803 24599
rect 8110 24596 8116 24608
rect 7791 24568 8116 24596
rect 7791 24565 7803 24568
rect 7745 24559 7803 24565
rect 8110 24556 8116 24568
rect 8168 24556 8174 24608
rect 8294 24556 8300 24608
rect 8352 24596 8358 24608
rect 8389 24599 8447 24605
rect 8389 24596 8401 24599
rect 8352 24568 8401 24596
rect 8352 24556 8358 24568
rect 8389 24565 8401 24568
rect 8435 24565 8447 24599
rect 8389 24559 8447 24565
rect 8938 24556 8944 24608
rect 8996 24596 9002 24608
rect 9125 24599 9183 24605
rect 9125 24596 9137 24599
rect 8996 24568 9137 24596
rect 8996 24556 9002 24568
rect 9125 24565 9137 24568
rect 9171 24565 9183 24599
rect 9950 24596 9956 24608
rect 9911 24568 9956 24596
rect 9125 24559 9183 24565
rect 9950 24556 9956 24568
rect 10008 24556 10014 24608
rect 12158 24596 12164 24608
rect 12119 24568 12164 24596
rect 12158 24556 12164 24568
rect 12216 24556 12222 24608
rect 12802 24556 12808 24608
rect 12860 24596 12866 24608
rect 13265 24599 13323 24605
rect 13265 24596 13277 24599
rect 12860 24568 13277 24596
rect 12860 24556 12866 24568
rect 13265 24565 13277 24568
rect 13311 24596 13323 24599
rect 13725 24599 13783 24605
rect 13725 24596 13737 24599
rect 13311 24568 13737 24596
rect 13311 24565 13323 24568
rect 13265 24559 13323 24565
rect 13725 24565 13737 24568
rect 13771 24565 13783 24599
rect 14366 24596 14372 24608
rect 14327 24568 14372 24596
rect 13725 24559 13783 24565
rect 14366 24556 14372 24568
rect 14424 24556 14430 24608
rect 15930 24596 15936 24608
rect 15891 24568 15936 24596
rect 15930 24556 15936 24568
rect 15988 24556 15994 24608
rect 17034 24556 17040 24608
rect 17092 24596 17098 24608
rect 17221 24599 17279 24605
rect 17221 24596 17233 24599
rect 17092 24568 17233 24596
rect 17092 24556 17098 24568
rect 17221 24565 17233 24568
rect 17267 24565 17279 24599
rect 17221 24559 17279 24565
rect 1104 24506 44896 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 44896 24506
rect 1104 24432 44896 24454
rect 1673 24395 1731 24401
rect 1673 24361 1685 24395
rect 1719 24392 1731 24395
rect 1762 24392 1768 24404
rect 1719 24364 1768 24392
rect 1719 24361 1731 24364
rect 1673 24355 1731 24361
rect 1762 24352 1768 24364
rect 1820 24352 1826 24404
rect 1857 24395 1915 24401
rect 1857 24361 1869 24395
rect 1903 24392 1915 24395
rect 2682 24392 2688 24404
rect 1903 24364 2688 24392
rect 1903 24361 1915 24364
rect 1857 24355 1915 24361
rect 2682 24352 2688 24364
rect 2740 24352 2746 24404
rect 11514 24392 11520 24404
rect 11475 24364 11520 24392
rect 11514 24352 11520 24364
rect 11572 24352 11578 24404
rect 12066 24352 12072 24404
rect 12124 24392 12130 24404
rect 12529 24395 12587 24401
rect 12529 24392 12541 24395
rect 12124 24364 12541 24392
rect 12124 24352 12130 24364
rect 12529 24361 12541 24364
rect 12575 24361 12587 24395
rect 12529 24355 12587 24361
rect 13170 24352 13176 24404
rect 13228 24392 13234 24404
rect 14737 24395 14795 24401
rect 14737 24392 14749 24395
rect 13228 24364 14749 24392
rect 13228 24352 13234 24364
rect 14737 24361 14749 24364
rect 14783 24392 14795 24395
rect 15194 24392 15200 24404
rect 14783 24364 15200 24392
rect 14783 24361 14795 24364
rect 14737 24355 14795 24361
rect 15194 24352 15200 24364
rect 15252 24352 15258 24404
rect 16298 24392 16304 24404
rect 16259 24364 16304 24392
rect 16298 24352 16304 24364
rect 16356 24352 16362 24404
rect 17218 24352 17224 24404
rect 17276 24392 17282 24404
rect 17402 24392 17408 24404
rect 17276 24364 17408 24392
rect 17276 24352 17282 24364
rect 17402 24352 17408 24364
rect 17460 24352 17466 24404
rect 17770 24352 17776 24404
rect 17828 24392 17834 24404
rect 18782 24392 18788 24404
rect 17828 24364 18788 24392
rect 17828 24352 17834 24364
rect 18782 24352 18788 24364
rect 18840 24352 18846 24404
rect 19150 24352 19156 24404
rect 19208 24392 19214 24404
rect 19337 24395 19395 24401
rect 19337 24392 19349 24395
rect 19208 24364 19349 24392
rect 19208 24352 19214 24364
rect 19337 24361 19349 24364
rect 19383 24392 19395 24395
rect 19978 24392 19984 24404
rect 19383 24364 19984 24392
rect 19383 24361 19395 24364
rect 19337 24355 19395 24361
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 22094 24352 22100 24404
rect 22152 24392 22158 24404
rect 22152 24364 22197 24392
rect 22152 24352 22158 24364
rect 7742 24324 7748 24336
rect 7703 24296 7748 24324
rect 7742 24284 7748 24296
rect 7800 24284 7806 24336
rect 9401 24327 9459 24333
rect 9401 24293 9413 24327
rect 9447 24324 9459 24327
rect 9582 24324 9588 24336
rect 9447 24296 9588 24324
rect 9447 24293 9459 24296
rect 9401 24287 9459 24293
rect 9582 24284 9588 24296
rect 9640 24284 9646 24336
rect 9858 24284 9864 24336
rect 9916 24324 9922 24336
rect 13081 24327 13139 24333
rect 13081 24324 13093 24327
rect 9916 24296 13093 24324
rect 9916 24284 9922 24296
rect 13081 24293 13093 24296
rect 13127 24293 13139 24327
rect 13081 24287 13139 24293
rect 13630 24284 13636 24336
rect 13688 24324 13694 24336
rect 13688 24296 20024 24324
rect 13688 24284 13694 24296
rect 19996 24268 20024 24296
rect 1578 24256 1584 24268
rect 1539 24228 1584 24256
rect 1578 24216 1584 24228
rect 1636 24216 1642 24268
rect 9030 24256 9036 24268
rect 8991 24228 9036 24256
rect 9030 24216 9036 24228
rect 9088 24216 9094 24268
rect 9493 24259 9551 24265
rect 9493 24225 9505 24259
rect 9539 24256 9551 24259
rect 14182 24256 14188 24268
rect 9539 24228 12572 24256
rect 14095 24228 14188 24256
rect 9539 24225 9551 24228
rect 9493 24219 9551 24225
rect 1670 24188 1676 24200
rect 1631 24160 1676 24188
rect 1670 24148 1676 24160
rect 1728 24148 1734 24200
rect 5718 24148 5724 24200
rect 5776 24188 5782 24200
rect 7193 24191 7251 24197
rect 7193 24188 7205 24191
rect 5776 24160 7205 24188
rect 5776 24148 5782 24160
rect 7193 24157 7205 24160
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 9674 24148 9680 24200
rect 9732 24188 9738 24200
rect 10689 24191 10747 24197
rect 10689 24188 10701 24191
rect 9732 24160 10701 24188
rect 9732 24148 9738 24160
rect 10689 24157 10701 24160
rect 10735 24157 10747 24191
rect 11330 24188 11336 24200
rect 11291 24160 11336 24188
rect 10689 24151 10747 24157
rect 11330 24148 11336 24160
rect 11388 24148 11394 24200
rect 11977 24191 12035 24197
rect 11977 24188 11989 24191
rect 11440 24160 11989 24188
rect 1394 24120 1400 24132
rect 1355 24092 1400 24120
rect 1394 24080 1400 24092
rect 1452 24080 1458 24132
rect 5074 24120 5080 24132
rect 3804 24092 5080 24120
rect 2406 24052 2412 24064
rect 2367 24024 2412 24052
rect 2406 24012 2412 24024
rect 2464 24012 2470 24064
rect 2866 24052 2872 24064
rect 2827 24024 2872 24052
rect 2866 24012 2872 24024
rect 2924 24012 2930 24064
rect 3694 24012 3700 24064
rect 3752 24052 3758 24064
rect 3804 24061 3832 24092
rect 5074 24080 5080 24092
rect 5132 24080 5138 24132
rect 6270 24080 6276 24132
rect 6328 24120 6334 24132
rect 7926 24120 7932 24132
rect 6328 24092 7932 24120
rect 6328 24080 6334 24092
rect 7926 24080 7932 24092
rect 7984 24080 7990 24132
rect 8110 24120 8116 24132
rect 8071 24092 8116 24120
rect 8110 24080 8116 24092
rect 8168 24080 8174 24132
rect 10042 24120 10048 24132
rect 10003 24092 10048 24120
rect 10042 24080 10048 24092
rect 10100 24080 10106 24132
rect 10134 24080 10140 24132
rect 10192 24120 10198 24132
rect 10229 24123 10287 24129
rect 10229 24120 10241 24123
rect 10192 24092 10241 24120
rect 10192 24080 10198 24092
rect 10229 24089 10241 24092
rect 10275 24089 10287 24123
rect 11440 24120 11468 24160
rect 11977 24157 11989 24160
rect 12023 24188 12035 24191
rect 12066 24188 12072 24200
rect 12023 24160 12072 24188
rect 12023 24157 12035 24160
rect 11977 24151 12035 24157
rect 12066 24148 12072 24160
rect 12124 24148 12130 24200
rect 10229 24083 10287 24089
rect 10428 24092 11468 24120
rect 3789 24055 3847 24061
rect 3789 24052 3801 24055
rect 3752 24024 3801 24052
rect 3752 24012 3758 24024
rect 3789 24021 3801 24024
rect 3835 24021 3847 24055
rect 3789 24015 3847 24021
rect 3970 24012 3976 24064
rect 4028 24052 4034 24064
rect 4341 24055 4399 24061
rect 4341 24052 4353 24055
rect 4028 24024 4353 24052
rect 4028 24012 4034 24024
rect 4341 24021 4353 24024
rect 4387 24021 4399 24055
rect 4341 24015 4399 24021
rect 4798 24012 4804 24064
rect 4856 24052 4862 24064
rect 4893 24055 4951 24061
rect 4893 24052 4905 24055
rect 4856 24024 4905 24052
rect 4856 24012 4862 24024
rect 4893 24021 4905 24024
rect 4939 24021 4951 24055
rect 4893 24015 4951 24021
rect 5537 24055 5595 24061
rect 5537 24021 5549 24055
rect 5583 24052 5595 24055
rect 5994 24052 6000 24064
rect 5583 24024 6000 24052
rect 5583 24021 5595 24024
rect 5537 24015 5595 24021
rect 5994 24012 6000 24024
rect 6052 24012 6058 24064
rect 6454 24052 6460 24064
rect 6415 24024 6460 24052
rect 6454 24012 6460 24024
rect 6512 24012 6518 24064
rect 7006 24052 7012 24064
rect 6967 24024 7012 24052
rect 7006 24012 7012 24024
rect 7064 24012 7070 24064
rect 7650 24052 7656 24064
rect 7611 24024 7656 24052
rect 7650 24012 7656 24024
rect 7708 24012 7714 24064
rect 8570 24012 8576 24064
rect 8628 24052 8634 24064
rect 10428 24052 10456 24092
rect 11790 24080 11796 24132
rect 11848 24120 11854 24132
rect 12544 24120 12572 24228
rect 14182 24216 14188 24228
rect 14240 24256 14246 24268
rect 14240 24228 18920 24256
rect 14240 24216 14246 24228
rect 13630 24148 13636 24200
rect 13688 24188 13694 24200
rect 15289 24191 15347 24197
rect 15289 24188 15301 24191
rect 13688 24160 15301 24188
rect 13688 24148 13694 24160
rect 15289 24157 15301 24160
rect 15335 24188 15347 24191
rect 18782 24188 18788 24200
rect 15335 24160 18788 24188
rect 15335 24157 15347 24160
rect 15289 24151 15347 24157
rect 18782 24148 18788 24160
rect 18840 24148 18846 24200
rect 18892 24188 18920 24228
rect 19978 24216 19984 24268
rect 20036 24216 20042 24268
rect 21726 24188 21732 24200
rect 18892 24160 21732 24188
rect 21726 24148 21732 24160
rect 21784 24148 21790 24200
rect 28994 24148 29000 24200
rect 29052 24188 29058 24200
rect 38654 24188 38660 24200
rect 29052 24160 38660 24188
rect 29052 24148 29058 24160
rect 38654 24148 38660 24160
rect 38712 24148 38718 24200
rect 14090 24120 14096 24132
rect 11848 24092 12434 24120
rect 12544 24092 14096 24120
rect 11848 24080 11854 24092
rect 8628 24024 10456 24052
rect 10873 24055 10931 24061
rect 8628 24012 8634 24024
rect 10873 24021 10885 24055
rect 10919 24052 10931 24055
rect 11422 24052 11428 24064
rect 10919 24024 11428 24052
rect 10919 24021 10931 24024
rect 10873 24015 10931 24021
rect 11422 24012 11428 24024
rect 11480 24012 11486 24064
rect 12406 24052 12434 24092
rect 14090 24080 14096 24092
rect 14148 24080 14154 24132
rect 17957 24123 18015 24129
rect 17957 24120 17969 24123
rect 16868 24092 17969 24120
rect 16868 24064 16896 24092
rect 17957 24089 17969 24092
rect 18003 24089 18015 24123
rect 17957 24083 18015 24089
rect 18601 24123 18659 24129
rect 18601 24089 18613 24123
rect 18647 24120 18659 24123
rect 19334 24120 19340 24132
rect 18647 24092 19340 24120
rect 18647 24089 18659 24092
rect 18601 24083 18659 24089
rect 19334 24080 19340 24092
rect 19392 24120 19398 24132
rect 20254 24120 20260 24132
rect 19392 24092 20260 24120
rect 19392 24080 19398 24092
rect 20254 24080 20260 24092
rect 20312 24080 20318 24132
rect 27154 24080 27160 24132
rect 27212 24120 27218 24132
rect 35986 24120 35992 24132
rect 27212 24092 35992 24120
rect 27212 24080 27218 24092
rect 35986 24080 35992 24092
rect 36044 24080 36050 24132
rect 14182 24052 14188 24064
rect 12406 24024 14188 24052
rect 14182 24012 14188 24024
rect 14240 24012 14246 24064
rect 15746 24052 15752 24064
rect 15707 24024 15752 24052
rect 15746 24012 15752 24024
rect 15804 24012 15810 24064
rect 16850 24052 16856 24064
rect 16811 24024 16856 24052
rect 16850 24012 16856 24024
rect 16908 24012 16914 24064
rect 17218 24012 17224 24064
rect 17276 24052 17282 24064
rect 29914 24052 29920 24064
rect 17276 24024 29920 24052
rect 17276 24012 17282 24024
rect 29914 24012 29920 24024
rect 29972 24012 29978 24064
rect 1104 23962 44896 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 44896 23962
rect 1104 23888 44896 23910
rect 1394 23848 1400 23860
rect 1355 23820 1400 23848
rect 1394 23808 1400 23820
rect 1452 23808 1458 23860
rect 2866 23808 2872 23860
rect 2924 23848 2930 23860
rect 2924 23820 4016 23848
rect 2924 23808 2930 23820
rect 1026 23740 1032 23792
rect 1084 23780 1090 23792
rect 3329 23783 3387 23789
rect 3329 23780 3341 23783
rect 1084 23752 3341 23780
rect 1084 23740 1090 23752
rect 1486 23672 1492 23724
rect 1544 23712 1550 23724
rect 1581 23715 1639 23721
rect 1581 23712 1593 23715
rect 1544 23684 1593 23712
rect 1544 23672 1550 23684
rect 1581 23681 1593 23684
rect 1627 23681 1639 23715
rect 1581 23675 1639 23681
rect 2317 23579 2375 23585
rect 2317 23545 2329 23579
rect 2363 23576 2375 23579
rect 2958 23576 2964 23588
rect 2363 23548 2964 23576
rect 2363 23545 2375 23548
rect 2317 23539 2375 23545
rect 2958 23536 2964 23548
rect 3016 23536 3022 23588
rect 2866 23508 2872 23520
rect 2827 23480 2872 23508
rect 2866 23468 2872 23480
rect 2924 23468 2930 23520
rect 3068 23508 3096 23752
rect 3329 23749 3341 23752
rect 3375 23749 3387 23783
rect 3988 23780 4016 23820
rect 4062 23808 4068 23860
rect 4120 23848 4126 23860
rect 9861 23851 9919 23857
rect 4120 23820 9536 23848
rect 4120 23808 4126 23820
rect 4157 23783 4215 23789
rect 4157 23780 4169 23783
rect 3988 23752 4169 23780
rect 3329 23743 3387 23749
rect 4157 23749 4169 23752
rect 4203 23780 4215 23783
rect 4982 23780 4988 23792
rect 4203 23752 4988 23780
rect 4203 23749 4215 23752
rect 4157 23743 4215 23749
rect 4982 23740 4988 23752
rect 5040 23740 5046 23792
rect 5074 23740 5080 23792
rect 5132 23780 5138 23792
rect 7745 23783 7803 23789
rect 7745 23780 7757 23783
rect 5132 23752 7757 23780
rect 5132 23740 5138 23752
rect 7745 23749 7757 23752
rect 7791 23749 7803 23783
rect 7745 23743 7803 23749
rect 7926 23740 7932 23792
rect 7984 23780 7990 23792
rect 8205 23783 8263 23789
rect 8205 23780 8217 23783
rect 7984 23752 8217 23780
rect 7984 23740 7990 23752
rect 8205 23749 8217 23752
rect 8251 23780 8263 23783
rect 8846 23780 8852 23792
rect 8251 23752 8852 23780
rect 8251 23749 8263 23752
rect 8205 23743 8263 23749
rect 8846 23740 8852 23752
rect 8904 23740 8910 23792
rect 9030 23740 9036 23792
rect 9088 23780 9094 23792
rect 9401 23783 9459 23789
rect 9401 23780 9413 23783
rect 9088 23752 9413 23780
rect 9088 23740 9094 23752
rect 9401 23749 9413 23752
rect 9447 23749 9459 23783
rect 9401 23743 9459 23749
rect 3418 23672 3424 23724
rect 3476 23712 3482 23724
rect 5813 23715 5871 23721
rect 5813 23712 5825 23715
rect 3476 23684 5825 23712
rect 3476 23672 3482 23684
rect 5813 23681 5825 23684
rect 5859 23681 5871 23715
rect 5813 23675 5871 23681
rect 6454 23672 6460 23724
rect 6512 23712 6518 23724
rect 6825 23715 6883 23721
rect 6825 23712 6837 23715
rect 6512 23684 6837 23712
rect 6512 23672 6518 23684
rect 6825 23681 6837 23684
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 8481 23715 8539 23721
rect 8481 23681 8493 23715
rect 8527 23712 8539 23715
rect 8754 23712 8760 23724
rect 8527 23684 8760 23712
rect 8527 23681 8539 23684
rect 8481 23675 8539 23681
rect 8754 23672 8760 23684
rect 8812 23672 8818 23724
rect 8297 23647 8355 23653
rect 8297 23644 8309 23647
rect 7392 23616 8309 23644
rect 3234 23536 3240 23588
rect 3292 23576 3298 23588
rect 3602 23576 3608 23588
rect 3292 23548 3608 23576
rect 3292 23536 3298 23548
rect 3602 23536 3608 23548
rect 3660 23576 3666 23588
rect 4709 23579 4767 23585
rect 4709 23576 4721 23579
rect 3660 23548 4721 23576
rect 3660 23536 3666 23548
rect 4709 23545 4721 23548
rect 4755 23545 4767 23579
rect 5626 23576 5632 23588
rect 5587 23548 5632 23576
rect 4709 23539 4767 23545
rect 5626 23536 5632 23548
rect 5684 23536 5690 23588
rect 6178 23536 6184 23588
rect 6236 23576 6242 23588
rect 7285 23579 7343 23585
rect 7285 23576 7297 23579
rect 6236 23548 7297 23576
rect 6236 23536 6242 23548
rect 7285 23545 7297 23548
rect 7331 23545 7343 23579
rect 7285 23539 7343 23545
rect 6641 23511 6699 23517
rect 6641 23508 6653 23511
rect 3068 23480 6653 23508
rect 6641 23477 6653 23480
rect 6687 23508 6699 23511
rect 7190 23508 7196 23520
rect 6687 23480 7196 23508
rect 6687 23477 6699 23480
rect 6641 23471 6699 23477
rect 7190 23468 7196 23480
rect 7248 23508 7254 23520
rect 7392 23508 7420 23616
rect 8297 23613 8309 23616
rect 8343 23644 8355 23647
rect 9214 23644 9220 23656
rect 8343 23616 9220 23644
rect 8343 23613 8355 23616
rect 8297 23607 8355 23613
rect 9214 23604 9220 23616
rect 9272 23604 9278 23656
rect 9508 23644 9536 23820
rect 9861 23817 9873 23851
rect 9907 23848 9919 23851
rect 11330 23848 11336 23860
rect 9907 23820 11336 23848
rect 9907 23817 9919 23820
rect 9861 23811 9919 23817
rect 11330 23808 11336 23820
rect 11388 23808 11394 23860
rect 11606 23808 11612 23860
rect 11664 23848 11670 23860
rect 14274 23848 14280 23860
rect 11664 23820 14136 23848
rect 14235 23820 14280 23848
rect 11664 23808 11670 23820
rect 10410 23740 10416 23792
rect 10468 23780 10474 23792
rect 10689 23783 10747 23789
rect 10689 23780 10701 23783
rect 10468 23752 10701 23780
rect 10468 23740 10474 23752
rect 10689 23749 10701 23752
rect 10735 23749 10747 23783
rect 11698 23780 11704 23792
rect 11659 23752 11704 23780
rect 10689 23743 10747 23749
rect 11698 23740 11704 23752
rect 11756 23740 11762 23792
rect 12342 23780 12348 23792
rect 11992 23752 12348 23780
rect 9950 23672 9956 23724
rect 10008 23712 10014 23724
rect 10505 23715 10563 23721
rect 10505 23712 10517 23715
rect 10008 23684 10517 23712
rect 10008 23672 10014 23684
rect 10505 23681 10517 23684
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 10781 23715 10839 23721
rect 10781 23681 10793 23715
rect 10827 23712 10839 23715
rect 10870 23712 10876 23724
rect 10827 23684 10876 23712
rect 10827 23681 10839 23684
rect 10781 23675 10839 23681
rect 10870 23672 10876 23684
rect 10928 23712 10934 23724
rect 11992 23712 12020 23752
rect 12342 23740 12348 23752
rect 12400 23740 12406 23792
rect 10928 23684 12020 23712
rect 10928 23672 10934 23684
rect 12066 23672 12072 23724
rect 12124 23712 12130 23724
rect 12253 23715 12311 23721
rect 12253 23712 12265 23715
rect 12124 23684 12265 23712
rect 12124 23672 12130 23684
rect 12253 23681 12265 23684
rect 12299 23681 12311 23715
rect 13078 23712 13084 23724
rect 13039 23684 13084 23712
rect 12253 23675 12311 23681
rect 13078 23672 13084 23684
rect 13136 23672 13142 23724
rect 13541 23715 13599 23721
rect 13541 23681 13553 23715
rect 13587 23681 13599 23715
rect 14108 23712 14136 23820
rect 14274 23808 14280 23820
rect 14332 23808 14338 23860
rect 15286 23848 15292 23860
rect 15199 23820 15292 23848
rect 15286 23808 15292 23820
rect 15344 23848 15350 23860
rect 15746 23848 15752 23860
rect 15344 23820 15752 23848
rect 15344 23808 15350 23820
rect 15746 23808 15752 23820
rect 15804 23808 15810 23860
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 17037 23851 17095 23857
rect 17037 23848 17049 23851
rect 16816 23820 17049 23848
rect 16816 23808 16822 23820
rect 17037 23817 17049 23820
rect 17083 23848 17095 23851
rect 17126 23848 17132 23860
rect 17083 23820 17132 23848
rect 17083 23817 17095 23820
rect 17037 23811 17095 23817
rect 17126 23808 17132 23820
rect 17184 23808 17190 23860
rect 18690 23848 18696 23860
rect 18651 23820 18696 23848
rect 18690 23808 18696 23820
rect 18748 23848 18754 23860
rect 18874 23848 18880 23860
rect 18748 23820 18880 23848
rect 18748 23808 18754 23820
rect 18874 23808 18880 23820
rect 18932 23808 18938 23860
rect 19889 23851 19947 23857
rect 19889 23817 19901 23851
rect 19935 23848 19947 23851
rect 20070 23848 20076 23860
rect 19935 23820 20076 23848
rect 19935 23817 19947 23820
rect 19889 23811 19947 23817
rect 20070 23808 20076 23820
rect 20128 23808 20134 23860
rect 28534 23848 28540 23860
rect 20180 23820 28540 23848
rect 16298 23740 16304 23792
rect 16356 23780 16362 23792
rect 17402 23780 17408 23792
rect 16356 23752 17408 23780
rect 16356 23740 16362 23752
rect 17402 23740 17408 23752
rect 17460 23780 17466 23792
rect 17589 23783 17647 23789
rect 17589 23780 17601 23783
rect 17460 23752 17601 23780
rect 17460 23740 17466 23752
rect 17589 23749 17601 23752
rect 17635 23749 17647 23783
rect 17589 23743 17647 23749
rect 19058 23712 19064 23724
rect 14108 23684 19064 23712
rect 13541 23675 13599 23681
rect 9508 23616 10456 23644
rect 10428 23588 10456 23616
rect 11974 23604 11980 23656
rect 12032 23644 12038 23656
rect 13556 23644 13584 23675
rect 19058 23672 19064 23684
rect 19116 23712 19122 23724
rect 19334 23712 19340 23724
rect 19116 23684 19340 23712
rect 19116 23672 19122 23684
rect 19334 23672 19340 23684
rect 19392 23672 19398 23724
rect 12032 23616 13584 23644
rect 12032 23604 12038 23616
rect 17678 23604 17684 23656
rect 17736 23644 17742 23656
rect 20180 23644 20208 23820
rect 28534 23808 28540 23820
rect 28592 23808 28598 23860
rect 22094 23740 22100 23792
rect 22152 23780 22158 23792
rect 22281 23783 22339 23789
rect 22281 23780 22293 23783
rect 22152 23752 22293 23780
rect 22152 23740 22158 23752
rect 22281 23749 22293 23752
rect 22327 23749 22339 23783
rect 22281 23743 22339 23749
rect 22465 23783 22523 23789
rect 22465 23749 22477 23783
rect 22511 23780 22523 23783
rect 30374 23780 30380 23792
rect 22511 23752 30380 23780
rect 22511 23749 22523 23752
rect 22465 23743 22523 23749
rect 30374 23740 30380 23752
rect 30432 23740 30438 23792
rect 32306 23672 32312 23724
rect 32364 23712 32370 23724
rect 32585 23715 32643 23721
rect 32585 23712 32597 23715
rect 32364 23684 32597 23712
rect 32364 23672 32370 23684
rect 32585 23681 32597 23684
rect 32631 23681 32643 23715
rect 32585 23675 32643 23681
rect 17736 23616 20208 23644
rect 17736 23604 17742 23616
rect 7469 23579 7527 23585
rect 7469 23545 7481 23579
rect 7515 23576 7527 23579
rect 8570 23576 8576 23588
rect 7515 23548 8576 23576
rect 7515 23545 7527 23548
rect 7469 23539 7527 23545
rect 8570 23536 8576 23548
rect 8628 23536 8634 23588
rect 8846 23536 8852 23588
rect 8904 23576 8910 23588
rect 9769 23579 9827 23585
rect 8904 23548 9720 23576
rect 8904 23536 8910 23548
rect 8294 23508 8300 23520
rect 7248 23480 7420 23508
rect 8255 23480 8300 23508
rect 7248 23468 7254 23480
rect 8294 23468 8300 23480
rect 8352 23468 8358 23520
rect 8665 23511 8723 23517
rect 8665 23477 8677 23511
rect 8711 23508 8723 23511
rect 9490 23508 9496 23520
rect 8711 23480 9496 23508
rect 8711 23477 8723 23480
rect 8665 23471 8723 23477
rect 9490 23468 9496 23480
rect 9548 23468 9554 23520
rect 9692 23508 9720 23548
rect 9769 23545 9781 23579
rect 9815 23576 9827 23579
rect 10042 23576 10048 23588
rect 9815 23548 10048 23576
rect 9815 23545 9827 23548
rect 9769 23539 9827 23545
rect 10042 23536 10048 23548
rect 10100 23536 10106 23588
rect 10410 23536 10416 23588
rect 10468 23536 10474 23588
rect 10502 23536 10508 23588
rect 10560 23576 10566 23588
rect 11514 23576 11520 23588
rect 10560 23548 10605 23576
rect 11475 23548 11520 23576
rect 10560 23536 10566 23548
rect 11514 23536 11520 23548
rect 11572 23536 11578 23588
rect 12710 23576 12716 23588
rect 11624 23548 12716 23576
rect 11624 23508 11652 23548
rect 12710 23536 12716 23548
rect 12768 23536 12774 23588
rect 12894 23576 12900 23588
rect 12855 23548 12900 23576
rect 12894 23536 12900 23548
rect 12952 23536 12958 23588
rect 13906 23536 13912 23588
rect 13964 23576 13970 23588
rect 30466 23576 30472 23588
rect 13964 23548 30472 23576
rect 13964 23536 13970 23548
rect 30466 23536 30472 23548
rect 30524 23536 30530 23588
rect 9692 23480 11652 23508
rect 12342 23468 12348 23520
rect 12400 23508 12406 23520
rect 12437 23511 12495 23517
rect 12437 23508 12449 23511
rect 12400 23480 12449 23508
rect 12400 23468 12406 23480
rect 12437 23477 12449 23480
rect 12483 23508 12495 23511
rect 13354 23508 13360 23520
rect 12483 23480 13360 23508
rect 12483 23477 12495 23480
rect 12437 23471 12495 23477
rect 13354 23468 13360 23480
rect 13412 23468 13418 23520
rect 13725 23511 13783 23517
rect 13725 23477 13737 23511
rect 13771 23508 13783 23511
rect 13998 23508 14004 23520
rect 13771 23480 14004 23508
rect 13771 23477 13783 23480
rect 13725 23471 13783 23477
rect 13998 23468 14004 23480
rect 14056 23468 14062 23520
rect 14366 23468 14372 23520
rect 14424 23508 14430 23520
rect 15841 23511 15899 23517
rect 15841 23508 15853 23511
rect 14424 23480 15853 23508
rect 14424 23468 14430 23480
rect 15841 23477 15853 23480
rect 15887 23508 15899 23511
rect 17770 23508 17776 23520
rect 15887 23480 17776 23508
rect 15887 23477 15899 23480
rect 15841 23471 15899 23477
rect 17770 23468 17776 23480
rect 17828 23468 17834 23520
rect 18233 23511 18291 23517
rect 18233 23477 18245 23511
rect 18279 23508 18291 23511
rect 18322 23508 18328 23520
rect 18279 23480 18328 23508
rect 18279 23477 18291 23480
rect 18233 23471 18291 23477
rect 18322 23468 18328 23480
rect 18380 23468 18386 23520
rect 19337 23511 19395 23517
rect 19337 23477 19349 23511
rect 19383 23508 19395 23511
rect 20254 23508 20260 23520
rect 19383 23480 20260 23508
rect 19383 23477 19395 23480
rect 19337 23471 19395 23477
rect 20254 23468 20260 23480
rect 20312 23508 20318 23520
rect 20714 23508 20720 23520
rect 20312 23480 20720 23508
rect 20312 23468 20318 23480
rect 20714 23468 20720 23480
rect 20772 23468 20778 23520
rect 32677 23511 32735 23517
rect 32677 23477 32689 23511
rect 32723 23508 32735 23511
rect 42242 23508 42248 23520
rect 32723 23480 42248 23508
rect 32723 23477 32735 23480
rect 32677 23471 32735 23477
rect 42242 23468 42248 23480
rect 42300 23468 42306 23520
rect 1104 23418 44896 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 44896 23418
rect 1104 23344 44896 23366
rect 1581 23307 1639 23313
rect 1581 23273 1593 23307
rect 1627 23304 1639 23307
rect 1670 23304 1676 23316
rect 1627 23276 1676 23304
rect 1627 23273 1639 23276
rect 1581 23267 1639 23273
rect 1670 23264 1676 23276
rect 1728 23264 1734 23316
rect 3234 23304 3240 23316
rect 3195 23276 3240 23304
rect 3234 23264 3240 23276
rect 3292 23264 3298 23316
rect 4890 23304 4896 23316
rect 4540 23276 4896 23304
rect 4540 23248 4568 23276
rect 4890 23264 4896 23276
rect 4948 23264 4954 23316
rect 4982 23264 4988 23316
rect 5040 23304 5046 23316
rect 5629 23307 5687 23313
rect 5629 23304 5641 23307
rect 5040 23276 5641 23304
rect 5040 23264 5046 23276
rect 5629 23273 5641 23276
rect 5675 23304 5687 23307
rect 6270 23304 6276 23316
rect 5675 23276 6276 23304
rect 5675 23273 5687 23276
rect 5629 23267 5687 23273
rect 6270 23264 6276 23276
rect 6328 23264 6334 23316
rect 6638 23264 6644 23316
rect 6696 23304 6702 23316
rect 6696 23276 7788 23304
rect 6696 23264 6702 23276
rect 4522 23196 4528 23248
rect 4580 23196 4586 23248
rect 5534 23236 5540 23248
rect 5092 23208 5540 23236
rect 1578 23128 1584 23180
rect 1636 23168 1642 23180
rect 2130 23168 2136 23180
rect 1636 23140 2136 23168
rect 1636 23128 1642 23140
rect 2130 23128 2136 23140
rect 2188 23128 2194 23180
rect 3881 23171 3939 23177
rect 3881 23137 3893 23171
rect 3927 23168 3939 23171
rect 5092 23168 5120 23208
rect 5534 23196 5540 23208
rect 5592 23196 5598 23248
rect 6457 23239 6515 23245
rect 6457 23205 6469 23239
rect 6503 23236 6515 23239
rect 6914 23236 6920 23248
rect 6503 23208 6920 23236
rect 6503 23205 6515 23208
rect 6457 23199 6515 23205
rect 6914 23196 6920 23208
rect 6972 23196 6978 23248
rect 7650 23168 7656 23180
rect 3927 23140 5120 23168
rect 5184 23140 7656 23168
rect 3927 23137 3939 23140
rect 3881 23131 3939 23137
rect 1394 23100 1400 23112
rect 1355 23072 1400 23100
rect 1394 23060 1400 23072
rect 1452 23100 1458 23112
rect 3786 23100 3792 23112
rect 1452 23072 3792 23100
rect 1452 23060 1458 23072
rect 3786 23060 3792 23072
rect 3844 23060 3850 23112
rect 1118 22992 1124 23044
rect 1176 23032 1182 23044
rect 3896 23032 3924 23131
rect 5184 23109 5212 23140
rect 7650 23128 7656 23140
rect 7708 23128 7714 23180
rect 7760 23177 7788 23276
rect 8294 23264 8300 23316
rect 8352 23304 8358 23316
rect 9125 23307 9183 23313
rect 9125 23304 9137 23307
rect 8352 23276 9137 23304
rect 8352 23264 8358 23276
rect 9125 23273 9137 23276
rect 9171 23273 9183 23307
rect 9125 23267 9183 23273
rect 11241 23307 11299 23313
rect 11241 23273 11253 23307
rect 11287 23304 11299 23307
rect 13078 23304 13084 23316
rect 11287 23276 13084 23304
rect 11287 23273 11299 23276
rect 11241 23267 11299 23273
rect 13078 23264 13084 23276
rect 13136 23264 13142 23316
rect 15565 23307 15623 23313
rect 15565 23273 15577 23307
rect 15611 23304 15623 23307
rect 16114 23304 16120 23316
rect 15611 23276 16120 23304
rect 15611 23273 15623 23276
rect 15565 23267 15623 23273
rect 16114 23264 16120 23276
rect 16172 23264 16178 23316
rect 16482 23264 16488 23316
rect 16540 23304 16546 23316
rect 16761 23307 16819 23313
rect 16761 23304 16773 23307
rect 16540 23276 16773 23304
rect 16540 23264 16546 23276
rect 16761 23273 16773 23276
rect 16807 23273 16819 23307
rect 17586 23304 17592 23316
rect 17547 23276 17592 23304
rect 16761 23267 16819 23273
rect 17586 23264 17592 23276
rect 17644 23264 17650 23316
rect 17770 23264 17776 23316
rect 17828 23304 17834 23316
rect 18598 23304 18604 23316
rect 17828 23276 18604 23304
rect 17828 23264 17834 23276
rect 18598 23264 18604 23276
rect 18656 23264 18662 23316
rect 20717 23307 20775 23313
rect 20717 23273 20729 23307
rect 20763 23304 20775 23307
rect 27062 23304 27068 23316
rect 20763 23276 27068 23304
rect 20763 23273 20775 23276
rect 20717 23267 20775 23273
rect 27062 23264 27068 23276
rect 27120 23264 27126 23316
rect 28442 23264 28448 23316
rect 28500 23304 28506 23316
rect 29822 23304 29828 23316
rect 28500 23276 29828 23304
rect 28500 23264 28506 23276
rect 29822 23264 29828 23276
rect 29880 23264 29886 23316
rect 7834 23196 7840 23248
rect 7892 23236 7898 23248
rect 8941 23239 8999 23245
rect 8941 23236 8953 23239
rect 7892 23208 8953 23236
rect 7892 23196 7898 23208
rect 8941 23205 8953 23208
rect 8987 23205 8999 23239
rect 8941 23199 8999 23205
rect 9030 23196 9036 23248
rect 9088 23236 9094 23248
rect 10229 23239 10287 23245
rect 9088 23208 10180 23236
rect 9088 23196 9094 23208
rect 7745 23171 7803 23177
rect 7745 23137 7757 23171
rect 7791 23137 7803 23171
rect 9214 23168 9220 23180
rect 9175 23140 9220 23168
rect 7745 23131 7803 23137
rect 9214 23128 9220 23140
rect 9272 23128 9278 23180
rect 9858 23168 9864 23180
rect 9819 23140 9864 23168
rect 9858 23128 9864 23140
rect 9916 23128 9922 23180
rect 10152 23168 10180 23208
rect 10229 23205 10241 23239
rect 10275 23236 10287 23239
rect 10318 23236 10324 23248
rect 10275 23208 10324 23236
rect 10275 23205 10287 23208
rect 10229 23199 10287 23205
rect 10318 23196 10324 23208
rect 10376 23196 10382 23248
rect 10962 23196 10968 23248
rect 11020 23236 11026 23248
rect 11057 23239 11115 23245
rect 11057 23236 11069 23239
rect 11020 23208 11069 23236
rect 11020 23196 11026 23208
rect 11057 23205 11069 23208
rect 11103 23205 11115 23239
rect 11057 23199 11115 23205
rect 11330 23196 11336 23248
rect 11388 23236 11394 23248
rect 11701 23239 11759 23245
rect 11701 23236 11713 23239
rect 11388 23208 11713 23236
rect 11388 23196 11394 23208
rect 11701 23205 11713 23208
rect 11747 23205 11759 23239
rect 11701 23199 11759 23205
rect 12158 23196 12164 23248
rect 12216 23236 12222 23248
rect 12216 23208 12848 23236
rect 12216 23196 12222 23208
rect 10778 23168 10784 23180
rect 10152 23140 10784 23168
rect 10778 23128 10784 23140
rect 10836 23128 10842 23180
rect 11514 23128 11520 23180
rect 11572 23168 11578 23180
rect 11572 23140 12664 23168
rect 11572 23128 11578 23140
rect 5169 23103 5227 23109
rect 5169 23069 5181 23103
rect 5215 23069 5227 23103
rect 5169 23063 5227 23069
rect 5813 23103 5871 23109
rect 5813 23069 5825 23103
rect 5859 23100 5871 23103
rect 5994 23100 6000 23112
rect 5859 23072 6000 23100
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 5994 23060 6000 23072
rect 6052 23060 6058 23112
rect 7561 23103 7619 23109
rect 7561 23069 7573 23103
rect 7607 23100 7619 23103
rect 8018 23100 8024 23112
rect 7607 23072 8024 23100
rect 7607 23069 7619 23072
rect 7561 23063 7619 23069
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 8754 23060 8760 23112
rect 8812 23100 8818 23112
rect 9125 23103 9183 23109
rect 9125 23100 9137 23103
rect 8812 23072 9137 23100
rect 8812 23060 8818 23072
rect 9125 23069 9137 23072
rect 9171 23069 9183 23103
rect 9125 23063 9183 23069
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 11977 23103 12035 23109
rect 9364 23072 11836 23100
rect 9364 23060 9370 23072
rect 1176 23004 3924 23032
rect 1176 22992 1182 23004
rect 4062 22992 4068 23044
rect 4120 23032 4126 23044
rect 4433 23035 4491 23041
rect 4433 23032 4445 23035
rect 4120 23004 4445 23032
rect 4120 22992 4126 23004
rect 4433 23001 4445 23004
rect 4479 23032 4491 23035
rect 4479 23004 5212 23032
rect 4479 23001 4491 23004
rect 4433 22995 4491 23001
rect 5184 22976 5212 23004
rect 5350 22992 5356 23044
rect 5408 23032 5414 23044
rect 6733 23035 6791 23041
rect 6733 23032 6745 23035
rect 5408 23004 6745 23032
rect 5408 22992 5414 23004
rect 6733 23001 6745 23004
rect 6779 23032 6791 23035
rect 8110 23032 8116 23044
rect 6779 23004 8116 23032
rect 6779 23001 6791 23004
rect 6733 22995 6791 23001
rect 8110 22992 8116 23004
rect 8168 22992 8174 23044
rect 8846 22992 8852 23044
rect 8904 23032 8910 23044
rect 9401 23035 9459 23041
rect 9401 23032 9413 23035
rect 8904 23004 9413 23032
rect 8904 22992 8910 23004
rect 9401 23001 9413 23004
rect 9447 23001 9459 23035
rect 9401 22995 9459 23001
rect 10042 22992 10048 23044
rect 10100 23032 10106 23044
rect 10226 23032 10232 23044
rect 10100 23004 10232 23032
rect 10100 22992 10106 23004
rect 10226 22992 10232 23004
rect 10284 22992 10290 23044
rect 11701 23035 11759 23041
rect 11701 23001 11713 23035
rect 11747 23001 11759 23035
rect 11808 23032 11836 23072
rect 11977 23069 11989 23103
rect 12023 23100 12035 23103
rect 12342 23100 12348 23112
rect 12023 23072 12348 23100
rect 12023 23069 12035 23072
rect 11977 23063 12035 23069
rect 12342 23060 12348 23072
rect 12400 23060 12406 23112
rect 12636 23109 12664 23140
rect 12621 23103 12679 23109
rect 12621 23069 12633 23103
rect 12667 23069 12679 23103
rect 12820 23100 12848 23208
rect 12894 23196 12900 23248
rect 12952 23236 12958 23248
rect 14366 23236 14372 23248
rect 12952 23208 14372 23236
rect 12952 23196 12958 23208
rect 14366 23196 14372 23208
rect 14424 23196 14430 23248
rect 18046 23236 18052 23248
rect 18007 23208 18052 23236
rect 18046 23196 18052 23208
rect 18104 23196 18110 23248
rect 21358 23236 21364 23248
rect 18156 23208 21364 23236
rect 14826 23128 14832 23180
rect 14884 23168 14890 23180
rect 18156 23168 18184 23208
rect 21358 23196 21364 23208
rect 21416 23196 21422 23248
rect 21542 23236 21548 23248
rect 21503 23208 21548 23236
rect 21542 23196 21548 23208
rect 21600 23196 21606 23248
rect 21634 23196 21640 23248
rect 21692 23236 21698 23248
rect 28721 23239 28779 23245
rect 21692 23208 22094 23236
rect 21692 23196 21698 23208
rect 19242 23168 19248 23180
rect 14884 23140 18184 23168
rect 19203 23140 19248 23168
rect 14884 23128 14890 23140
rect 19242 23128 19248 23140
rect 19300 23128 19306 23180
rect 19521 23171 19579 23177
rect 19521 23137 19533 23171
rect 19567 23168 19579 23171
rect 20438 23168 20444 23180
rect 19567 23140 20444 23168
rect 19567 23137 19579 23140
rect 19521 23131 19579 23137
rect 20438 23128 20444 23140
rect 20496 23128 20502 23180
rect 22066 23168 22094 23208
rect 28721 23205 28733 23239
rect 28767 23236 28779 23239
rect 38470 23236 38476 23248
rect 28767 23208 38476 23236
rect 28767 23205 28779 23208
rect 28721 23199 28779 23205
rect 38470 23196 38476 23208
rect 38528 23196 38534 23248
rect 30098 23168 30104 23180
rect 22066 23140 30104 23168
rect 30098 23128 30104 23140
rect 30156 23128 30162 23180
rect 30193 23171 30251 23177
rect 30193 23137 30205 23171
rect 30239 23168 30251 23171
rect 39206 23168 39212 23180
rect 30239 23140 39212 23168
rect 30239 23137 30251 23140
rect 30193 23131 30251 23137
rect 39206 23128 39212 23140
rect 39264 23128 39270 23180
rect 13173 23103 13231 23109
rect 13173 23100 13185 23103
rect 12820 23072 13185 23100
rect 12621 23063 12679 23069
rect 13173 23069 13185 23072
rect 13219 23069 13231 23103
rect 14090 23100 14096 23112
rect 14051 23072 14096 23100
rect 13173 23063 13231 23069
rect 12437 23035 12495 23041
rect 12437 23032 12449 23035
rect 11808 23004 12449 23032
rect 11701 22995 11759 23001
rect 12437 23001 12449 23004
rect 12483 23001 12495 23035
rect 13188 23032 13216 23063
rect 14090 23060 14096 23072
rect 14148 23060 14154 23112
rect 14366 23060 14372 23112
rect 14424 23100 14430 23112
rect 15930 23100 15936 23112
rect 14424 23072 15936 23100
rect 14424 23060 14430 23072
rect 15930 23060 15936 23072
rect 15988 23060 15994 23112
rect 17405 23103 17463 23109
rect 17405 23069 17417 23103
rect 17451 23100 17463 23103
rect 21266 23100 21272 23112
rect 17451 23072 21272 23100
rect 17451 23069 17463 23072
rect 17405 23063 17463 23069
rect 21266 23060 21272 23072
rect 21324 23060 21330 23112
rect 29546 23100 29552 23112
rect 25884 23072 29552 23100
rect 14734 23032 14740 23044
rect 13188 23004 14740 23032
rect 12437 22995 12495 23001
rect 2130 22964 2136 22976
rect 2091 22936 2136 22964
rect 2130 22924 2136 22936
rect 2188 22924 2194 22976
rect 2685 22967 2743 22973
rect 2685 22933 2697 22967
rect 2731 22964 2743 22967
rect 3786 22964 3792 22976
rect 2731 22936 3792 22964
rect 2731 22933 2743 22936
rect 2685 22927 2743 22933
rect 3786 22924 3792 22936
rect 3844 22924 3850 22976
rect 4982 22964 4988 22976
rect 4943 22936 4988 22964
rect 4982 22924 4988 22936
rect 5040 22924 5046 22976
rect 5166 22924 5172 22976
rect 5224 22924 5230 22976
rect 6270 22964 6276 22976
rect 6231 22936 6276 22964
rect 6270 22924 6276 22936
rect 6328 22924 6334 22976
rect 7190 22964 7196 22976
rect 7151 22936 7196 22964
rect 7190 22924 7196 22936
rect 7248 22924 7254 22976
rect 7653 22967 7711 22973
rect 7653 22933 7665 22967
rect 7699 22964 7711 22967
rect 8386 22964 8392 22976
rect 7699 22936 8392 22964
rect 7699 22933 7711 22936
rect 7653 22927 7711 22933
rect 8386 22924 8392 22936
rect 8444 22924 8450 22976
rect 10318 22964 10324 22976
rect 10279 22936 10324 22964
rect 10318 22924 10324 22936
rect 10376 22924 10382 22976
rect 10594 22924 10600 22976
rect 10652 22964 10658 22976
rect 10870 22964 10876 22976
rect 10652 22936 10876 22964
rect 10652 22924 10658 22936
rect 10870 22924 10876 22936
rect 10928 22924 10934 22976
rect 11716 22964 11744 22995
rect 14734 22992 14740 23004
rect 14792 22992 14798 23044
rect 17310 22992 17316 23044
rect 17368 23032 17374 23044
rect 17678 23032 17684 23044
rect 17368 23004 17684 23032
rect 17368 22992 17374 23004
rect 17678 22992 17684 23004
rect 17736 22992 17742 23044
rect 19334 22992 19340 23044
rect 19392 23032 19398 23044
rect 20625 23035 20683 23041
rect 20625 23032 20637 23035
rect 19392 23004 20637 23032
rect 19392 22992 19398 23004
rect 20625 23001 20637 23004
rect 20671 23001 20683 23035
rect 20625 22995 20683 23001
rect 21361 23035 21419 23041
rect 21361 23001 21373 23035
rect 21407 23001 21419 23035
rect 21361 22995 21419 23001
rect 22097 23035 22155 23041
rect 22097 23001 22109 23035
rect 22143 23032 22155 23035
rect 22278 23032 22284 23044
rect 22143 23004 22284 23032
rect 22143 23001 22155 23004
rect 22097 22995 22155 23001
rect 11790 22964 11796 22976
rect 11716 22936 11796 22964
rect 11790 22924 11796 22936
rect 11848 22924 11854 22976
rect 11885 22967 11943 22973
rect 11885 22933 11897 22967
rect 11931 22964 11943 22967
rect 12802 22964 12808 22976
rect 11931 22936 12808 22964
rect 11931 22933 11943 22936
rect 11885 22927 11943 22933
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 13357 22967 13415 22973
rect 13357 22933 13369 22967
rect 13403 22964 13415 22967
rect 13446 22964 13452 22976
rect 13403 22936 13452 22964
rect 13403 22933 13415 22936
rect 13357 22927 13415 22933
rect 13446 22924 13452 22936
rect 13504 22924 13510 22976
rect 14182 22924 14188 22976
rect 14240 22964 14246 22976
rect 14277 22967 14335 22973
rect 14277 22964 14289 22967
rect 14240 22936 14289 22964
rect 14240 22924 14246 22936
rect 14277 22933 14289 22936
rect 14323 22933 14335 22967
rect 16298 22964 16304 22976
rect 16259 22936 16304 22964
rect 14277 22927 14335 22933
rect 16298 22924 16304 22936
rect 16356 22924 16362 22976
rect 19242 22924 19248 22976
rect 19300 22964 19306 22976
rect 21376 22964 21404 22995
rect 22278 22992 22284 23004
rect 22336 22992 22342 23044
rect 19300 22936 21404 22964
rect 22189 22967 22247 22973
rect 19300 22924 19306 22936
rect 22189 22933 22201 22967
rect 22235 22964 22247 22967
rect 25884 22964 25912 23072
rect 29546 23060 29552 23072
rect 29604 23060 29610 23112
rect 30929 23103 30987 23109
rect 30929 23069 30941 23103
rect 30975 23100 30987 23103
rect 40586 23100 40592 23112
rect 30975 23072 40592 23100
rect 30975 23069 30987 23072
rect 30929 23063 30987 23069
rect 40586 23060 40592 23072
rect 40644 23060 40650 23112
rect 28537 23035 28595 23041
rect 28537 23001 28549 23035
rect 28583 23001 28595 23035
rect 30006 23032 30012 23044
rect 29967 23004 30012 23032
rect 28537 22995 28595 23001
rect 22235 22936 25912 22964
rect 27985 22967 28043 22973
rect 22235 22933 22247 22936
rect 22189 22927 22247 22933
rect 27985 22933 27997 22967
rect 28031 22964 28043 22967
rect 28552 22964 28580 22995
rect 30006 22992 30012 23004
rect 30064 22992 30070 23044
rect 30558 22992 30564 23044
rect 30616 23032 30622 23044
rect 30745 23035 30803 23041
rect 30745 23032 30757 23035
rect 30616 23004 30757 23032
rect 30616 22992 30622 23004
rect 30745 23001 30757 23004
rect 30791 23001 30803 23035
rect 30745 22995 30803 23001
rect 31294 22992 31300 23044
rect 31352 23032 31358 23044
rect 31481 23035 31539 23041
rect 31481 23032 31493 23035
rect 31352 23004 31493 23032
rect 31352 22992 31358 23004
rect 31481 23001 31493 23004
rect 31527 23001 31539 23035
rect 31481 22995 31539 23001
rect 31665 23035 31723 23041
rect 31665 23001 31677 23035
rect 31711 23032 31723 23035
rect 42426 23032 42432 23044
rect 31711 23004 42432 23032
rect 31711 23001 31723 23004
rect 31665 22995 31723 23001
rect 42426 22992 42432 23004
rect 42484 22992 42490 23044
rect 30926 22964 30932 22976
rect 28031 22936 30932 22964
rect 28031 22933 28043 22936
rect 27985 22927 28043 22933
rect 30926 22924 30932 22936
rect 30984 22924 30990 22976
rect 32306 22964 32312 22976
rect 32267 22936 32312 22964
rect 32306 22924 32312 22936
rect 32364 22924 32370 22976
rect 1104 22874 44896 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 44896 22874
rect 1104 22800 44896 22822
rect 1762 22720 1768 22772
rect 1820 22760 1826 22772
rect 2685 22763 2743 22769
rect 2685 22760 2697 22763
rect 1820 22732 2697 22760
rect 1820 22720 1826 22732
rect 2685 22729 2697 22732
rect 2731 22729 2743 22763
rect 2685 22723 2743 22729
rect 2866 22720 2872 22772
rect 2924 22760 2930 22772
rect 3513 22763 3571 22769
rect 3513 22760 3525 22763
rect 2924 22732 3525 22760
rect 2924 22720 2930 22732
rect 3513 22729 3525 22732
rect 3559 22729 3571 22763
rect 4706 22760 4712 22772
rect 4619 22732 4712 22760
rect 3513 22723 3571 22729
rect 4706 22720 4712 22732
rect 4764 22760 4770 22772
rect 5074 22760 5080 22772
rect 4764 22732 5080 22760
rect 4764 22720 4770 22732
rect 5074 22720 5080 22732
rect 5132 22720 5138 22772
rect 5813 22763 5871 22769
rect 5813 22729 5825 22763
rect 5859 22760 5871 22763
rect 5902 22760 5908 22772
rect 5859 22732 5908 22760
rect 5859 22729 5871 22732
rect 5813 22723 5871 22729
rect 5902 22720 5908 22732
rect 5960 22720 5966 22772
rect 7561 22763 7619 22769
rect 7561 22729 7573 22763
rect 7607 22760 7619 22763
rect 7742 22760 7748 22772
rect 7607 22732 7748 22760
rect 7607 22729 7619 22732
rect 7561 22723 7619 22729
rect 7742 22720 7748 22732
rect 7800 22720 7806 22772
rect 10428 22732 10824 22760
rect 10428 22704 10456 22732
rect 474 22652 480 22704
rect 532 22692 538 22704
rect 3694 22692 3700 22704
rect 532 22664 3700 22692
rect 532 22652 538 22664
rect 3694 22652 3700 22664
rect 3752 22692 3758 22704
rect 6270 22692 6276 22704
rect 3752 22664 4200 22692
rect 3752 22652 3758 22664
rect 1578 22624 1584 22636
rect 1539 22596 1584 22624
rect 1578 22584 1584 22596
rect 1636 22584 1642 22636
rect 2038 22624 2044 22636
rect 1951 22596 2044 22624
rect 2038 22584 2044 22596
rect 2096 22624 2102 22636
rect 2682 22624 2688 22636
rect 2096 22596 2688 22624
rect 2096 22584 2102 22596
rect 2682 22584 2688 22596
rect 2740 22584 2746 22636
rect 2866 22584 2872 22636
rect 2924 22624 2930 22636
rect 3878 22624 3884 22636
rect 2924 22596 3884 22624
rect 2924 22584 2930 22596
rect 3878 22584 3884 22596
rect 3936 22584 3942 22636
rect 2130 22516 2136 22568
rect 2188 22556 2194 22568
rect 2314 22556 2320 22568
rect 2188 22528 2320 22556
rect 2188 22516 2194 22528
rect 2314 22516 2320 22528
rect 2372 22556 2378 22568
rect 4172 22556 4200 22664
rect 4264 22664 6276 22692
rect 4264 22633 4292 22664
rect 6270 22652 6276 22664
rect 6328 22652 6334 22704
rect 7101 22695 7159 22701
rect 7101 22661 7113 22695
rect 7147 22692 7159 22695
rect 8754 22692 8760 22704
rect 7147 22664 8760 22692
rect 7147 22661 7159 22664
rect 7101 22655 7159 22661
rect 8754 22652 8760 22664
rect 8812 22652 8818 22704
rect 10226 22692 10232 22704
rect 10152 22664 10232 22692
rect 4249 22627 4307 22633
rect 4249 22593 4261 22627
rect 4295 22593 4307 22627
rect 4249 22587 4307 22593
rect 4893 22627 4951 22633
rect 4893 22593 4905 22627
rect 4939 22593 4951 22627
rect 4893 22587 4951 22593
rect 4908 22556 4936 22587
rect 5534 22584 5540 22636
rect 5592 22624 5598 22636
rect 6454 22624 6460 22636
rect 5592 22596 6460 22624
rect 5592 22584 5598 22596
rect 6454 22584 6460 22596
rect 6512 22624 6518 22636
rect 7193 22627 7251 22633
rect 6512 22596 7052 22624
rect 6512 22584 6518 22596
rect 2372 22528 2774 22556
rect 4172 22528 4936 22556
rect 2372 22516 2378 22528
rect 2746 22488 2774 22528
rect 5074 22516 5080 22568
rect 5132 22556 5138 22568
rect 5350 22556 5356 22568
rect 5132 22528 5356 22556
rect 5132 22516 5138 22528
rect 5350 22516 5356 22528
rect 5408 22516 5414 22568
rect 6178 22516 6184 22568
rect 6236 22556 6242 22568
rect 6638 22556 6644 22568
rect 6236 22528 6644 22556
rect 6236 22516 6242 22528
rect 6638 22516 6644 22528
rect 6696 22556 6702 22568
rect 6917 22559 6975 22565
rect 6917 22556 6929 22559
rect 6696 22528 6929 22556
rect 6696 22516 6702 22528
rect 6917 22525 6929 22528
rect 6963 22525 6975 22559
rect 7024 22556 7052 22596
rect 7193 22593 7205 22627
rect 7239 22624 7251 22627
rect 7558 22624 7564 22636
rect 7239 22596 7564 22624
rect 7239 22593 7251 22596
rect 7193 22587 7251 22593
rect 7558 22584 7564 22596
rect 7616 22584 7622 22636
rect 7926 22584 7932 22636
rect 7984 22624 7990 22636
rect 8573 22627 8631 22633
rect 8573 22624 8585 22627
rect 7984 22596 8585 22624
rect 7984 22584 7990 22596
rect 8573 22593 8585 22596
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 8849 22627 8907 22633
rect 8849 22593 8861 22627
rect 8895 22624 8907 22627
rect 9030 22624 9036 22636
rect 8895 22596 9036 22624
rect 8895 22593 8907 22596
rect 8849 22587 8907 22593
rect 9030 22584 9036 22596
rect 9088 22584 9094 22636
rect 10152 22633 10180 22664
rect 10226 22652 10232 22664
rect 10284 22652 10290 22704
rect 10410 22652 10416 22704
rect 10468 22652 10474 22704
rect 10796 22692 10824 22732
rect 10870 22720 10876 22772
rect 10928 22760 10934 22772
rect 11974 22760 11980 22772
rect 10928 22732 11560 22760
rect 11935 22732 11980 22760
rect 10928 22720 10934 22732
rect 11532 22701 11560 22732
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 12158 22720 12164 22772
rect 12216 22720 12222 22772
rect 12526 22760 12532 22772
rect 12439 22732 12532 22760
rect 12526 22720 12532 22732
rect 12584 22760 12590 22772
rect 12802 22760 12808 22772
rect 12584 22732 12808 22760
rect 12584 22720 12590 22732
rect 12802 22720 12808 22732
rect 12860 22720 12866 22772
rect 14826 22760 14832 22772
rect 14787 22732 14832 22760
rect 14826 22720 14832 22732
rect 14884 22720 14890 22772
rect 15838 22760 15844 22772
rect 15799 22732 15844 22760
rect 15838 22720 15844 22732
rect 15896 22720 15902 22772
rect 16022 22720 16028 22772
rect 16080 22760 16086 22772
rect 22370 22760 22376 22772
rect 16080 22732 22094 22760
rect 22331 22732 22376 22760
rect 16080 22720 16086 22732
rect 10965 22695 11023 22701
rect 10965 22692 10977 22695
rect 10796 22664 10977 22692
rect 10965 22661 10977 22664
rect 11011 22661 11023 22695
rect 10965 22655 11023 22661
rect 11517 22695 11575 22701
rect 11517 22661 11529 22695
rect 11563 22661 11575 22695
rect 11517 22655 11575 22661
rect 10137 22627 10195 22633
rect 10137 22593 10149 22627
rect 10183 22593 10195 22627
rect 10594 22624 10600 22636
rect 10555 22596 10600 22624
rect 10137 22587 10195 22593
rect 10594 22584 10600 22596
rect 10652 22584 10658 22636
rect 10778 22584 10784 22636
rect 10836 22624 10842 22636
rect 10836 22596 10881 22624
rect 10836 22584 10842 22596
rect 12176 22556 12204 22720
rect 12713 22695 12771 22701
rect 12713 22661 12725 22695
rect 12759 22692 12771 22695
rect 13170 22692 13176 22704
rect 12759 22664 13176 22692
rect 12759 22661 12771 22664
rect 12713 22655 12771 22661
rect 13170 22652 13176 22664
rect 13228 22652 13234 22704
rect 13722 22692 13728 22704
rect 13464 22664 13728 22692
rect 12434 22584 12440 22636
rect 12492 22624 12498 22636
rect 12894 22624 12900 22636
rect 12492 22596 12537 22624
rect 12636 22596 12900 22624
rect 12492 22584 12498 22596
rect 7024 22528 12204 22556
rect 6917 22519 6975 22525
rect 12636 22500 12664 22596
rect 12894 22584 12900 22596
rect 12952 22624 12958 22636
rect 13464 22633 13492 22664
rect 13722 22652 13728 22664
rect 13780 22652 13786 22704
rect 13814 22652 13820 22704
rect 13872 22692 13878 22704
rect 14001 22695 14059 22701
rect 14001 22692 14013 22695
rect 13872 22664 14013 22692
rect 13872 22652 13878 22664
rect 14001 22661 14013 22664
rect 14047 22692 14059 22695
rect 14366 22692 14372 22704
rect 14047 22664 14372 22692
rect 14047 22661 14059 22664
rect 14001 22655 14059 22661
rect 14366 22652 14372 22664
rect 14424 22652 14430 22704
rect 16761 22695 16819 22701
rect 16761 22661 16773 22695
rect 16807 22692 16819 22695
rect 17218 22692 17224 22704
rect 16807 22664 17224 22692
rect 16807 22661 16819 22664
rect 16761 22655 16819 22661
rect 17218 22652 17224 22664
rect 17276 22652 17282 22704
rect 21174 22692 21180 22704
rect 21135 22664 21180 22692
rect 21174 22652 21180 22664
rect 21232 22652 21238 22704
rect 13449 22627 13507 22633
rect 12952 22596 13216 22624
rect 12952 22584 12958 22596
rect 13188 22565 13216 22596
rect 13449 22593 13461 22627
rect 13495 22593 13507 22627
rect 13630 22622 13636 22636
rect 13449 22587 13507 22593
rect 13556 22594 13636 22622
rect 13173 22559 13231 22565
rect 13173 22525 13185 22559
rect 13219 22525 13231 22559
rect 13173 22519 13231 22525
rect 13357 22559 13415 22565
rect 13357 22525 13369 22559
rect 13403 22556 13415 22559
rect 13556 22556 13584 22594
rect 13630 22584 13636 22594
rect 13688 22584 13694 22636
rect 14642 22624 14648 22636
rect 14603 22596 14648 22624
rect 14642 22584 14648 22596
rect 14700 22624 14706 22636
rect 15289 22627 15347 22633
rect 15289 22624 15301 22627
rect 14700 22596 15301 22624
rect 14700 22584 14706 22596
rect 15289 22593 15301 22596
rect 15335 22593 15347 22627
rect 17862 22624 17868 22636
rect 17823 22596 17868 22624
rect 15289 22587 15347 22593
rect 17862 22584 17868 22596
rect 17920 22584 17926 22636
rect 18230 22584 18236 22636
rect 18288 22624 18294 22636
rect 19153 22627 19211 22633
rect 19153 22624 19165 22627
rect 18288 22596 19165 22624
rect 18288 22584 18294 22596
rect 19153 22593 19165 22596
rect 19199 22593 19211 22627
rect 19153 22587 19211 22593
rect 19429 22627 19487 22633
rect 19429 22593 19441 22627
rect 19475 22624 19487 22627
rect 20162 22624 20168 22636
rect 19475 22596 20024 22624
rect 20123 22596 20168 22624
rect 19475 22593 19487 22596
rect 19429 22587 19487 22593
rect 18138 22556 18144 22568
rect 13403 22528 13584 22556
rect 18099 22528 18144 22556
rect 13403 22525 13415 22528
rect 13357 22519 13415 22525
rect 18138 22516 18144 22528
rect 18196 22516 18202 22568
rect 19886 22556 19892 22568
rect 19847 22528 19892 22556
rect 19886 22516 19892 22528
rect 19944 22516 19950 22568
rect 19996 22556 20024 22596
rect 20162 22584 20168 22596
rect 20220 22584 20226 22636
rect 22066 22624 22094 22732
rect 22370 22720 22376 22732
rect 22428 22720 22434 22772
rect 29822 22760 29828 22772
rect 29735 22732 29828 22760
rect 29822 22720 29828 22732
rect 29880 22760 29886 22772
rect 30006 22760 30012 22772
rect 29880 22732 30012 22760
rect 29880 22720 29886 22732
rect 30006 22720 30012 22732
rect 30064 22720 30070 22772
rect 30098 22720 30104 22772
rect 30156 22760 30162 22772
rect 34698 22760 34704 22772
rect 30156 22732 34704 22760
rect 30156 22720 30162 22732
rect 34698 22720 34704 22732
rect 34756 22720 34762 22772
rect 22186 22652 22192 22704
rect 22244 22692 22250 22704
rect 22281 22695 22339 22701
rect 22281 22692 22293 22695
rect 22244 22664 22293 22692
rect 22244 22652 22250 22664
rect 22281 22661 22293 22664
rect 22327 22661 22339 22695
rect 22281 22655 22339 22661
rect 22554 22624 22560 22636
rect 22066 22596 22560 22624
rect 22554 22584 22560 22596
rect 22612 22584 22618 22636
rect 29178 22556 29184 22568
rect 19996 22528 29184 22556
rect 29178 22516 29184 22528
rect 29236 22516 29242 22568
rect 5721 22491 5779 22497
rect 2746 22460 4200 22488
rect 1394 22420 1400 22432
rect 1355 22392 1400 22420
rect 1394 22380 1400 22392
rect 1452 22380 1458 22432
rect 4062 22420 4068 22432
rect 4023 22392 4068 22420
rect 4062 22380 4068 22392
rect 4120 22380 4126 22432
rect 4172 22420 4200 22460
rect 5721 22457 5733 22491
rect 5767 22488 5779 22491
rect 7190 22488 7196 22500
rect 5767 22460 7196 22488
rect 5767 22457 5779 22460
rect 5721 22451 5779 22457
rect 7190 22448 7196 22460
rect 7248 22448 7254 22500
rect 9907 22491 9965 22497
rect 9907 22457 9919 22491
rect 9953 22488 9965 22491
rect 10410 22488 10416 22500
rect 9953 22460 10416 22488
rect 9953 22457 9965 22460
rect 9907 22451 9965 22457
rect 10410 22448 10416 22460
rect 10468 22448 10474 22500
rect 10870 22448 10876 22500
rect 10928 22488 10934 22500
rect 11054 22488 11060 22500
rect 10928 22460 11060 22488
rect 10928 22448 10934 22460
rect 11054 22448 11060 22460
rect 11112 22448 11118 22500
rect 11882 22488 11888 22500
rect 11843 22460 11888 22488
rect 11882 22448 11888 22460
rect 11940 22448 11946 22500
rect 12618 22448 12624 22500
rect 12676 22448 12682 22500
rect 14185 22491 14243 22497
rect 14185 22457 14197 22491
rect 14231 22488 14243 22491
rect 21082 22488 21088 22500
rect 14231 22460 21088 22488
rect 14231 22457 14243 22460
rect 14185 22451 14243 22457
rect 21082 22448 21088 22460
rect 21140 22448 21146 22500
rect 21266 22448 21272 22500
rect 21324 22488 21330 22500
rect 26234 22488 26240 22500
rect 21324 22460 26240 22488
rect 21324 22448 21330 22460
rect 26234 22448 26240 22460
rect 26292 22448 26298 22500
rect 5994 22420 6000 22432
rect 4172 22392 6000 22420
rect 5994 22380 6000 22392
rect 6052 22380 6058 22432
rect 6086 22380 6092 22432
rect 6144 22420 6150 22432
rect 6454 22420 6460 22432
rect 6144 22392 6460 22420
rect 6144 22380 6150 22392
rect 6454 22380 6460 22392
rect 6512 22380 6518 22432
rect 8662 22380 8668 22432
rect 8720 22420 8726 22432
rect 10778 22420 10784 22432
rect 8720 22392 10784 22420
rect 8720 22380 8726 22392
rect 10778 22380 10784 22392
rect 10836 22380 10842 22432
rect 12710 22420 12716 22432
rect 12671 22392 12716 22420
rect 12710 22380 12716 22392
rect 12768 22380 12774 22432
rect 13449 22423 13507 22429
rect 13449 22389 13461 22423
rect 13495 22420 13507 22423
rect 13906 22420 13912 22432
rect 13495 22392 13912 22420
rect 13495 22389 13507 22392
rect 13449 22383 13507 22389
rect 13906 22380 13912 22392
rect 13964 22380 13970 22432
rect 15562 22380 15568 22432
rect 15620 22420 15626 22432
rect 16022 22420 16028 22432
rect 15620 22392 16028 22420
rect 15620 22380 15626 22392
rect 16022 22380 16028 22392
rect 16080 22380 16086 22432
rect 30558 22420 30564 22432
rect 30519 22392 30564 22420
rect 30558 22380 30564 22392
rect 30616 22380 30622 22432
rect 31294 22420 31300 22432
rect 31255 22392 31300 22420
rect 31294 22380 31300 22392
rect 31352 22380 31358 22432
rect 1104 22330 44896 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 44896 22330
rect 1104 22256 44896 22278
rect 3418 22176 3424 22228
rect 3476 22216 3482 22228
rect 5534 22216 5540 22228
rect 3476 22188 5540 22216
rect 3476 22176 3482 22188
rect 5534 22176 5540 22188
rect 5592 22176 5598 22228
rect 5994 22176 6000 22228
rect 6052 22176 6058 22228
rect 6914 22216 6920 22228
rect 6875 22188 6920 22216
rect 6914 22176 6920 22188
rect 6972 22176 6978 22228
rect 7558 22176 7564 22228
rect 7616 22216 7622 22228
rect 10778 22216 10784 22228
rect 7616 22188 10784 22216
rect 7616 22176 7622 22188
rect 10778 22176 10784 22188
rect 10836 22176 10842 22228
rect 10962 22216 10968 22228
rect 10923 22188 10968 22216
rect 10962 22176 10968 22188
rect 11020 22176 11026 22228
rect 14642 22216 14648 22228
rect 11072 22188 14648 22216
rect 1946 22108 1952 22160
rect 2004 22148 2010 22160
rect 2590 22148 2596 22160
rect 2004 22120 2596 22148
rect 2004 22108 2010 22120
rect 2590 22108 2596 22120
rect 2648 22108 2654 22160
rect 3234 22108 3240 22160
rect 3292 22148 3298 22160
rect 4617 22151 4675 22157
rect 4617 22148 4629 22151
rect 3292 22120 4629 22148
rect 3292 22108 3298 22120
rect 4617 22117 4629 22120
rect 4663 22117 4675 22151
rect 5626 22148 5632 22160
rect 4617 22111 4675 22117
rect 4724 22120 5488 22148
rect 5587 22120 5632 22148
rect 2958 22080 2964 22092
rect 2700 22052 2964 22080
rect 1397 22015 1455 22021
rect 1397 21981 1409 22015
rect 1443 21981 1455 22015
rect 2222 22012 2228 22024
rect 2183 21984 2228 22012
rect 1397 21975 1455 21981
rect 1412 21944 1440 21975
rect 2222 21972 2228 21984
rect 2280 22012 2286 22024
rect 2700 22012 2728 22052
rect 2958 22040 2964 22052
rect 3016 22040 3022 22092
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 3694 22080 3700 22092
rect 3200 22052 3700 22080
rect 3200 22040 3206 22052
rect 3694 22040 3700 22052
rect 3752 22040 3758 22092
rect 3786 22040 3792 22092
rect 3844 22080 3850 22092
rect 4724 22080 4752 22120
rect 3844 22052 4752 22080
rect 4801 22083 4859 22089
rect 3844 22040 3850 22052
rect 4801 22049 4813 22083
rect 4847 22080 4859 22083
rect 5258 22080 5264 22092
rect 4847 22052 5264 22080
rect 4847 22049 4859 22052
rect 4801 22043 4859 22049
rect 5258 22040 5264 22052
rect 5316 22040 5322 22092
rect 2280 21984 2728 22012
rect 2280 21972 2286 21984
rect 2774 21972 2780 22024
rect 2832 22012 2838 22024
rect 2869 22015 2927 22021
rect 2869 22012 2881 22015
rect 2832 21984 2881 22012
rect 2832 21972 2838 21984
rect 2869 21981 2881 21984
rect 2915 22012 2927 22015
rect 3510 22012 3516 22024
rect 2915 21984 3516 22012
rect 2915 21981 2927 21984
rect 2869 21975 2927 21981
rect 3510 21972 3516 21984
rect 3568 21972 3574 22024
rect 4706 21972 4712 22024
rect 4764 22012 4770 22024
rect 5460 22012 5488 22120
rect 5626 22108 5632 22120
rect 5684 22108 5690 22160
rect 6012 22148 6040 22176
rect 11072 22148 11100 22188
rect 14642 22176 14648 22188
rect 14700 22176 14706 22228
rect 22097 22219 22155 22225
rect 14752 22188 19334 22216
rect 6012 22120 11100 22148
rect 11146 22108 11152 22160
rect 11204 22148 11210 22160
rect 11701 22151 11759 22157
rect 11701 22148 11713 22151
rect 11204 22120 11713 22148
rect 11204 22108 11210 22120
rect 11701 22117 11713 22120
rect 11747 22117 11759 22151
rect 11701 22111 11759 22117
rect 12713 22151 12771 22157
rect 12713 22117 12725 22151
rect 12759 22148 12771 22151
rect 12894 22148 12900 22160
rect 12759 22120 12900 22148
rect 12759 22117 12771 22120
rect 12713 22111 12771 22117
rect 12894 22108 12900 22120
rect 12952 22108 12958 22160
rect 13446 22108 13452 22160
rect 13504 22148 13510 22160
rect 14752 22148 14780 22188
rect 13504 22120 14780 22148
rect 13504 22108 13510 22120
rect 15194 22108 15200 22160
rect 15252 22148 15258 22160
rect 19306 22148 19334 22188
rect 22097 22185 22109 22219
rect 22143 22216 22155 22219
rect 22186 22216 22192 22228
rect 22143 22188 22192 22216
rect 22143 22185 22155 22188
rect 22097 22179 22155 22185
rect 22186 22176 22192 22188
rect 22244 22176 22250 22228
rect 26142 22148 26148 22160
rect 15252 22120 18276 22148
rect 19306 22120 26148 22148
rect 15252 22108 15258 22120
rect 5718 22080 5724 22092
rect 5679 22052 5724 22080
rect 5718 22040 5724 22052
rect 5776 22040 5782 22092
rect 6178 22040 6184 22092
rect 6236 22080 6242 22092
rect 6273 22083 6331 22089
rect 6273 22080 6285 22083
rect 6236 22052 6285 22080
rect 6236 22040 6242 22052
rect 6273 22049 6285 22052
rect 6319 22049 6331 22083
rect 10318 22080 10324 22092
rect 10279 22052 10324 22080
rect 6273 22043 6331 22049
rect 10318 22040 10324 22052
rect 10376 22040 10382 22092
rect 10410 22040 10416 22092
rect 10468 22080 10474 22092
rect 10686 22080 10692 22092
rect 10468 22052 10692 22080
rect 10468 22040 10474 22052
rect 10686 22040 10692 22052
rect 10744 22040 10750 22092
rect 15378 22080 15384 22092
rect 11072 22052 15240 22080
rect 15339 22052 15384 22080
rect 7558 22012 7564 22024
rect 4764 21984 5212 22012
rect 5460 21984 7564 22012
rect 4764 21972 4770 21984
rect 5184 21956 5212 21984
rect 7558 21972 7564 21984
rect 7616 21972 7622 22024
rect 7926 22012 7932 22024
rect 7887 21984 7932 22012
rect 7926 21972 7932 21984
rect 7984 21972 7990 22024
rect 8110 21972 8116 22024
rect 8168 22012 8174 22024
rect 8205 22015 8263 22021
rect 8205 22012 8217 22015
rect 8168 21984 8217 22012
rect 8168 21972 8174 21984
rect 8205 21981 8217 21984
rect 8251 21981 8263 22015
rect 8205 21975 8263 21981
rect 8478 21972 8484 22024
rect 8536 22012 8542 22024
rect 9493 22015 9551 22021
rect 9493 22012 9505 22015
rect 8536 21984 9505 22012
rect 8536 21972 8542 21984
rect 9493 21981 9505 21984
rect 9539 21981 9551 22015
rect 9493 21975 9551 21981
rect 9769 22015 9827 22021
rect 9769 21981 9781 22015
rect 9815 22012 9827 22015
rect 11072 22012 11100 22052
rect 12066 22012 12072 22024
rect 9815 21984 11100 22012
rect 11164 21984 12072 22012
rect 9815 21981 9827 21984
rect 9769 21975 9827 21981
rect 1854 21944 1860 21956
rect 1412 21916 1860 21944
rect 1854 21904 1860 21916
rect 1912 21944 1918 21956
rect 1912 21916 3096 21944
rect 1912 21904 1918 21916
rect 1578 21876 1584 21888
rect 1539 21848 1584 21876
rect 1578 21836 1584 21848
rect 1636 21836 1642 21888
rect 1670 21836 1676 21888
rect 1728 21876 1734 21888
rect 2041 21879 2099 21885
rect 2041 21876 2053 21879
rect 1728 21848 2053 21876
rect 1728 21836 1734 21848
rect 2041 21845 2053 21848
rect 2087 21845 2099 21879
rect 2041 21839 2099 21845
rect 2222 21836 2228 21888
rect 2280 21876 2286 21888
rect 2685 21879 2743 21885
rect 2685 21876 2697 21879
rect 2280 21848 2697 21876
rect 2280 21836 2286 21848
rect 2685 21845 2697 21848
rect 2731 21845 2743 21879
rect 3068 21876 3096 21916
rect 3142 21904 3148 21956
rect 3200 21944 3206 21956
rect 4341 21947 4399 21953
rect 4341 21944 4353 21947
rect 3200 21916 4353 21944
rect 3200 21904 3206 21916
rect 4341 21913 4353 21916
rect 4387 21944 4399 21947
rect 5074 21944 5080 21956
rect 4387 21916 5080 21944
rect 4387 21913 4399 21916
rect 4341 21907 4399 21913
rect 5074 21904 5080 21916
rect 5132 21904 5138 21956
rect 5166 21904 5172 21956
rect 5224 21944 5230 21956
rect 5261 21947 5319 21953
rect 5261 21944 5273 21947
rect 5224 21916 5273 21944
rect 5224 21904 5230 21916
rect 5261 21913 5273 21916
rect 5307 21913 5319 21947
rect 5261 21907 5319 21913
rect 5534 21904 5540 21956
rect 5592 21944 5598 21956
rect 8938 21944 8944 21956
rect 5592 21916 8944 21944
rect 5592 21904 5598 21916
rect 8938 21904 8944 21916
rect 8996 21944 9002 21956
rect 11164 21944 11192 21984
rect 12066 21972 12072 21984
rect 12124 21972 12130 22024
rect 12342 22012 12348 22024
rect 12303 21984 12348 22012
rect 12342 21972 12348 21984
rect 12400 21972 12406 22024
rect 12710 21972 12716 22024
rect 12768 22012 12774 22024
rect 13265 22015 13323 22021
rect 13265 22012 13277 22015
rect 12768 21984 13277 22012
rect 12768 21972 12774 21984
rect 13265 21981 13277 21984
rect 13311 21981 13323 22015
rect 13265 21975 13323 21981
rect 13357 22015 13415 22021
rect 13357 21981 13369 22015
rect 13403 22012 13415 22015
rect 13403 21984 13768 22012
rect 13403 21981 13415 21984
rect 13357 21975 13415 21981
rect 8996 21916 11192 21944
rect 11425 21947 11483 21953
rect 8996 21904 9002 21916
rect 11425 21913 11437 21947
rect 11471 21944 11483 21947
rect 11606 21944 11612 21956
rect 11471 21916 11612 21944
rect 11471 21913 11483 21916
rect 11425 21907 11483 21913
rect 3510 21876 3516 21888
rect 3068 21848 3516 21876
rect 2685 21839 2743 21845
rect 3510 21836 3516 21848
rect 3568 21836 3574 21888
rect 6270 21836 6276 21888
rect 6328 21876 6334 21888
rect 6457 21879 6515 21885
rect 6457 21876 6469 21879
rect 6328 21848 6469 21876
rect 6328 21836 6334 21848
rect 6457 21845 6469 21848
rect 6503 21845 6515 21879
rect 6457 21839 6515 21845
rect 6549 21879 6607 21885
rect 6549 21845 6561 21879
rect 6595 21876 6607 21879
rect 6914 21876 6920 21888
rect 6595 21848 6920 21876
rect 6595 21845 6607 21848
rect 6549 21839 6607 21845
rect 6914 21836 6920 21848
rect 6972 21836 6978 21888
rect 8294 21836 8300 21888
rect 8352 21876 8358 21888
rect 9122 21876 9128 21888
rect 8352 21848 9128 21876
rect 8352 21836 8358 21848
rect 9122 21836 9128 21848
rect 9180 21836 9186 21888
rect 10042 21836 10048 21888
rect 10100 21876 10106 21888
rect 10502 21876 10508 21888
rect 10100 21848 10508 21876
rect 10100 21836 10106 21848
rect 10502 21836 10508 21848
rect 10560 21836 10566 21888
rect 10594 21836 10600 21888
rect 10652 21876 10658 21888
rect 10652 21848 10697 21876
rect 10652 21836 10658 21848
rect 10962 21836 10968 21888
rect 11020 21876 11026 21888
rect 11440 21876 11468 21907
rect 11606 21904 11612 21916
rect 11664 21904 11670 21956
rect 12618 21904 12624 21956
rect 12676 21944 12682 21956
rect 13541 21947 13599 21953
rect 13541 21944 13553 21947
rect 12676 21916 13553 21944
rect 12676 21904 12682 21916
rect 13541 21913 13553 21916
rect 13587 21913 13599 21947
rect 13740 21944 13768 21984
rect 14090 21972 14096 22024
rect 14148 22012 14154 22024
rect 14277 22015 14335 22021
rect 14148 21984 14193 22012
rect 14148 21972 14154 21984
rect 14277 21981 14289 22015
rect 14323 22012 14335 22015
rect 14826 22012 14832 22024
rect 14323 21984 14832 22012
rect 14323 21981 14335 21984
rect 14277 21975 14335 21981
rect 14826 21972 14832 21984
rect 14884 21972 14890 22024
rect 15212 22012 15240 22052
rect 15378 22040 15384 22052
rect 15436 22040 15442 22092
rect 16298 22080 16304 22092
rect 15580 22052 16304 22080
rect 15580 22012 15608 22052
rect 16298 22040 16304 22052
rect 16356 22040 16362 22092
rect 16758 22040 16764 22092
rect 16816 22080 16822 22092
rect 17402 22080 17408 22092
rect 16816 22052 17408 22080
rect 16816 22040 16822 22052
rect 17402 22040 17408 22052
rect 17460 22040 17466 22092
rect 15212 21984 15608 22012
rect 15657 22015 15715 22021
rect 15657 21981 15669 22015
rect 15703 21981 15715 22015
rect 16850 22012 16856 22024
rect 16811 21984 16856 22012
rect 15657 21975 15715 21981
rect 15194 21944 15200 21956
rect 13740 21916 15200 21944
rect 13541 21907 13599 21913
rect 15194 21904 15200 21916
rect 15252 21904 15258 21956
rect 15672 21944 15700 21975
rect 16850 21972 16856 21984
rect 16908 21972 16914 22024
rect 17129 22015 17187 22021
rect 17129 21981 17141 22015
rect 17175 22012 17187 22015
rect 18138 22012 18144 22024
rect 17175 21984 18144 22012
rect 17175 21981 17187 21984
rect 17129 21975 17187 21981
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 18248 22012 18276 22120
rect 26142 22108 26148 22120
rect 26200 22108 26206 22160
rect 18414 22040 18420 22092
rect 18472 22080 18478 22092
rect 18509 22083 18567 22089
rect 18509 22080 18521 22083
rect 18472 22052 18521 22080
rect 18472 22040 18478 22052
rect 18509 22049 18521 22052
rect 18555 22049 18567 22083
rect 18509 22043 18567 22049
rect 19058 22040 19064 22092
rect 19116 22080 19122 22092
rect 19334 22080 19340 22092
rect 19116 22052 19340 22080
rect 19116 22040 19122 22052
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 19426 22040 19432 22092
rect 19484 22080 19490 22092
rect 19521 22083 19579 22089
rect 19521 22080 19533 22083
rect 19484 22052 19533 22080
rect 19484 22040 19490 22052
rect 19521 22049 19533 22052
rect 19567 22049 19579 22083
rect 20530 22080 20536 22092
rect 20491 22052 20536 22080
rect 19521 22043 19579 22049
rect 20530 22040 20536 22052
rect 20588 22040 20594 22092
rect 20254 22012 20260 22024
rect 18248 21984 20260 22012
rect 20254 21972 20260 21984
rect 20312 21972 20318 22024
rect 20809 22015 20867 22021
rect 20809 21981 20821 22015
rect 20855 22012 20867 22015
rect 31294 22012 31300 22024
rect 20855 21984 31300 22012
rect 20855 21981 20867 21984
rect 20809 21975 20867 21981
rect 31294 21972 31300 21984
rect 31352 21972 31358 22024
rect 17770 21944 17776 21956
rect 15672 21916 17776 21944
rect 17770 21904 17776 21916
rect 17828 21904 17834 21956
rect 18322 21944 18328 21956
rect 18283 21916 18328 21944
rect 18322 21904 18328 21916
rect 18380 21904 18386 21956
rect 19242 21904 19248 21956
rect 19300 21944 19306 21956
rect 19337 21947 19395 21953
rect 19337 21944 19349 21947
rect 19300 21916 19349 21944
rect 19300 21904 19306 21916
rect 19337 21913 19349 21916
rect 19383 21944 19395 21947
rect 21269 21947 21327 21953
rect 21269 21944 21281 21947
rect 19383 21916 21281 21944
rect 19383 21913 19395 21916
rect 19337 21907 19395 21913
rect 21269 21913 21281 21916
rect 21315 21913 21327 21947
rect 21269 21907 21327 21913
rect 11882 21876 11888 21888
rect 11020 21848 11468 21876
rect 11843 21848 11888 21876
rect 11020 21836 11026 21848
rect 11882 21836 11888 21848
rect 11940 21836 11946 21888
rect 12802 21876 12808 21888
rect 12763 21848 12808 21876
rect 12802 21836 12808 21848
rect 12860 21836 12866 21888
rect 12894 21836 12900 21888
rect 12952 21876 12958 21888
rect 13170 21876 13176 21888
rect 12952 21848 13176 21876
rect 12952 21836 12958 21848
rect 13170 21836 13176 21848
rect 13228 21836 13234 21888
rect 13265 21879 13323 21885
rect 13265 21845 13277 21879
rect 13311 21876 13323 21879
rect 15746 21876 15752 21888
rect 13311 21848 15752 21876
rect 13311 21845 13323 21848
rect 13265 21839 13323 21845
rect 15746 21836 15752 21848
rect 15804 21836 15810 21888
rect 17402 21836 17408 21888
rect 17460 21876 17466 21888
rect 17589 21879 17647 21885
rect 17589 21876 17601 21879
rect 17460 21848 17601 21876
rect 17460 21836 17466 21848
rect 17589 21845 17601 21848
rect 17635 21845 17647 21879
rect 17589 21839 17647 21845
rect 1104 21786 44896 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 44896 21786
rect 1104 21712 44896 21734
rect 1673 21675 1731 21681
rect 1673 21641 1685 21675
rect 1719 21672 1731 21675
rect 2590 21672 2596 21684
rect 1719 21644 2596 21672
rect 1719 21641 1731 21644
rect 1673 21635 1731 21641
rect 2590 21632 2596 21644
rect 2648 21632 2654 21684
rect 2961 21675 3019 21681
rect 2961 21641 2973 21675
rect 3007 21672 3019 21675
rect 4062 21672 4068 21684
rect 3007 21644 4068 21672
rect 3007 21641 3019 21644
rect 2961 21635 3019 21641
rect 4062 21632 4068 21644
rect 4120 21632 4126 21684
rect 5902 21672 5908 21684
rect 5276 21644 5908 21672
rect 1486 21536 1492 21548
rect 1447 21508 1492 21536
rect 1486 21496 1492 21508
rect 1544 21496 1550 21548
rect 2317 21539 2375 21545
rect 2317 21505 2329 21539
rect 2363 21536 2375 21539
rect 2498 21536 2504 21548
rect 2363 21508 2504 21536
rect 2363 21505 2375 21508
rect 2317 21499 2375 21505
rect 2498 21496 2504 21508
rect 2556 21496 2562 21548
rect 2777 21539 2835 21545
rect 2777 21505 2789 21539
rect 2823 21505 2835 21539
rect 2777 21499 2835 21505
rect 2792 21468 2820 21499
rect 3050 21496 3056 21548
rect 3108 21536 3114 21548
rect 3513 21539 3571 21545
rect 3513 21536 3525 21539
rect 3108 21508 3525 21536
rect 3108 21496 3114 21508
rect 3513 21505 3525 21508
rect 3559 21505 3571 21539
rect 3513 21499 3571 21505
rect 3697 21539 3755 21545
rect 3697 21505 3709 21539
rect 3743 21536 3755 21539
rect 3786 21536 3792 21548
rect 3743 21508 3792 21536
rect 3743 21505 3755 21508
rect 3697 21499 3755 21505
rect 3786 21496 3792 21508
rect 3844 21536 3850 21548
rect 5276 21536 5304 21644
rect 5902 21632 5908 21644
rect 5960 21632 5966 21684
rect 10318 21672 10324 21684
rect 7668 21644 10324 21672
rect 5350 21564 5356 21616
rect 5408 21604 5414 21616
rect 6457 21607 6515 21613
rect 6457 21604 6469 21607
rect 5408 21576 6469 21604
rect 5408 21564 5414 21576
rect 6457 21573 6469 21576
rect 6503 21573 6515 21607
rect 6638 21604 6644 21616
rect 6599 21576 6644 21604
rect 6457 21567 6515 21573
rect 6638 21564 6644 21576
rect 6696 21564 6702 21616
rect 5442 21536 5448 21548
rect 3844 21508 5304 21536
rect 5403 21508 5448 21536
rect 3844 21496 3850 21508
rect 5442 21496 5448 21508
rect 5500 21496 5506 21548
rect 4157 21471 4215 21477
rect 4157 21468 4169 21471
rect 2792 21440 4169 21468
rect 4157 21437 4169 21440
rect 4203 21437 4215 21471
rect 4617 21471 4675 21477
rect 4157 21431 4215 21437
rect 4264 21440 4568 21468
rect 1486 21360 1492 21412
rect 1544 21400 1550 21412
rect 2133 21403 2191 21409
rect 2133 21400 2145 21403
rect 1544 21372 2145 21400
rect 1544 21360 1550 21372
rect 2133 21369 2145 21372
rect 2179 21369 2191 21403
rect 2133 21363 2191 21369
rect 3878 21292 3884 21344
rect 3936 21332 3942 21344
rect 4264 21332 4292 21440
rect 4341 21403 4399 21409
rect 4341 21369 4353 21403
rect 4387 21369 4399 21403
rect 4540 21400 4568 21440
rect 4617 21437 4629 21471
rect 4663 21468 4675 21471
rect 5166 21468 5172 21480
rect 4663 21440 5172 21468
rect 4663 21437 4675 21440
rect 4617 21431 4675 21437
rect 5166 21428 5172 21440
rect 5224 21428 5230 21480
rect 5258 21428 5264 21480
rect 5316 21468 5322 21480
rect 5537 21471 5595 21477
rect 5537 21468 5549 21471
rect 5316 21440 5549 21468
rect 5316 21428 5322 21440
rect 5537 21437 5549 21440
rect 5583 21437 5595 21471
rect 5537 21431 5595 21437
rect 5629 21471 5687 21477
rect 5629 21437 5641 21471
rect 5675 21468 5687 21471
rect 7668 21468 7696 21644
rect 10318 21632 10324 21644
rect 10376 21672 10382 21684
rect 11330 21672 11336 21684
rect 10376 21644 11336 21672
rect 10376 21632 10382 21644
rect 11330 21632 11336 21644
rect 11388 21632 11394 21684
rect 11606 21632 11612 21684
rect 11664 21672 11670 21684
rect 12618 21672 12624 21684
rect 11664 21644 12624 21672
rect 11664 21632 11670 21644
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 13170 21672 13176 21684
rect 13131 21644 13176 21672
rect 13170 21632 13176 21644
rect 13228 21632 13234 21684
rect 13354 21632 13360 21684
rect 13412 21672 13418 21684
rect 23750 21672 23756 21684
rect 13412 21644 23756 21672
rect 13412 21632 13418 21644
rect 23750 21632 23756 21644
rect 23808 21632 23814 21684
rect 27706 21672 27712 21684
rect 27667 21644 27712 21672
rect 27706 21632 27712 21644
rect 27764 21632 27770 21684
rect 8849 21607 8907 21613
rect 8849 21573 8861 21607
rect 8895 21604 8907 21607
rect 11790 21604 11796 21616
rect 8895 21576 11796 21604
rect 8895 21573 8907 21576
rect 8849 21567 8907 21573
rect 11790 21564 11796 21576
rect 11848 21564 11854 21616
rect 12250 21564 12256 21616
rect 12308 21604 12314 21616
rect 13633 21607 13691 21613
rect 13633 21604 13645 21607
rect 12308 21576 13645 21604
rect 12308 21564 12314 21576
rect 13633 21573 13645 21576
rect 13679 21573 13691 21607
rect 13633 21567 13691 21573
rect 14550 21564 14556 21616
rect 14608 21604 14614 21616
rect 17310 21604 17316 21616
rect 14608 21576 17316 21604
rect 14608 21564 14614 21576
rect 17310 21564 17316 21576
rect 17368 21564 17374 21616
rect 19886 21564 19892 21616
rect 19944 21604 19950 21616
rect 22278 21604 22284 21616
rect 19944 21576 22284 21604
rect 19944 21564 19950 21576
rect 22278 21564 22284 21576
rect 22336 21564 22342 21616
rect 22922 21604 22928 21616
rect 22883 21576 22928 21604
rect 22922 21564 22928 21576
rect 22980 21604 22986 21616
rect 23106 21604 23112 21616
rect 22980 21576 23112 21604
rect 22980 21564 22986 21576
rect 23106 21564 23112 21576
rect 23164 21564 23170 21616
rect 9490 21536 9496 21548
rect 9451 21508 9496 21536
rect 9490 21496 9496 21508
rect 9548 21496 9554 21548
rect 9674 21496 9680 21548
rect 9732 21536 9738 21548
rect 9732 21508 10640 21536
rect 9732 21496 9738 21508
rect 8018 21468 8024 21480
rect 5675 21440 7696 21468
rect 7979 21440 8024 21468
rect 5675 21437 5687 21440
rect 5629 21431 5687 21437
rect 5644 21400 5672 21431
rect 8018 21428 8024 21440
rect 8076 21428 8082 21480
rect 9033 21471 9091 21477
rect 9033 21437 9045 21471
rect 9079 21437 9091 21471
rect 9033 21431 9091 21437
rect 8294 21400 8300 21412
rect 4540 21372 5672 21400
rect 7024 21372 8300 21400
rect 4341 21363 4399 21369
rect 3936 21304 4292 21332
rect 4356 21332 4384 21363
rect 4614 21332 4620 21344
rect 4356 21304 4620 21332
rect 3936 21292 3942 21304
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 4706 21292 4712 21344
rect 4764 21332 4770 21344
rect 5077 21335 5135 21341
rect 5077 21332 5089 21335
rect 4764 21304 5089 21332
rect 4764 21292 4770 21304
rect 5077 21301 5089 21304
rect 5123 21301 5135 21335
rect 5077 21295 5135 21301
rect 5258 21292 5264 21344
rect 5316 21332 5322 21344
rect 7024 21332 7052 21372
rect 8294 21360 8300 21372
rect 8352 21360 8358 21412
rect 8386 21360 8392 21412
rect 8444 21400 8450 21412
rect 9048 21400 9076 21431
rect 8444 21372 9076 21400
rect 8444 21360 8450 21372
rect 9122 21360 9128 21412
rect 9180 21400 9186 21412
rect 10410 21400 10416 21412
rect 9180 21372 10416 21400
rect 9180 21360 9186 21372
rect 10410 21360 10416 21372
rect 10468 21360 10474 21412
rect 10612 21400 10640 21508
rect 10686 21496 10692 21548
rect 10744 21536 10750 21548
rect 10965 21539 11023 21545
rect 10965 21536 10977 21539
rect 10744 21508 10977 21536
rect 10744 21496 10750 21508
rect 10965 21505 10977 21508
rect 11011 21505 11023 21539
rect 10965 21499 11023 21505
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 12158 21536 12164 21548
rect 11931 21508 12164 21536
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 12158 21496 12164 21508
rect 12216 21536 12222 21548
rect 12434 21536 12440 21548
rect 12216 21508 12440 21536
rect 12216 21496 12222 21508
rect 12434 21496 12440 21508
rect 12492 21496 12498 21548
rect 13817 21539 13875 21545
rect 13817 21505 13829 21539
rect 13863 21536 13875 21539
rect 14274 21536 14280 21548
rect 13863 21508 14280 21536
rect 13863 21505 13875 21508
rect 13817 21499 13875 21505
rect 14274 21496 14280 21508
rect 14332 21496 14338 21548
rect 15470 21536 15476 21548
rect 15431 21508 15476 21536
rect 15470 21496 15476 21508
rect 15528 21496 15534 21548
rect 16942 21536 16948 21548
rect 16903 21508 16948 21536
rect 16942 21496 16948 21508
rect 17000 21496 17006 21548
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 19061 21539 19119 21545
rect 19061 21536 19073 21539
rect 18012 21508 19073 21536
rect 18012 21496 18018 21508
rect 19061 21505 19073 21508
rect 19107 21505 19119 21539
rect 20622 21536 20628 21548
rect 20583 21508 20628 21536
rect 19061 21499 19119 21505
rect 20622 21496 20628 21508
rect 20680 21496 20686 21548
rect 31202 21536 31208 21548
rect 20732 21508 31208 21536
rect 11977 21471 12035 21477
rect 11977 21437 11989 21471
rect 12023 21437 12035 21471
rect 11977 21431 12035 21437
rect 11517 21403 11575 21409
rect 11517 21400 11529 21403
rect 10612 21372 11529 21400
rect 11517 21369 11529 21372
rect 11563 21369 11575 21403
rect 11992 21400 12020 21431
rect 12066 21428 12072 21480
rect 12124 21468 12130 21480
rect 12124 21440 12169 21468
rect 12124 21428 12130 21440
rect 12618 21428 12624 21480
rect 12676 21468 12682 21480
rect 12713 21471 12771 21477
rect 12713 21468 12725 21471
rect 12676 21440 12725 21468
rect 12676 21428 12682 21440
rect 12713 21437 12725 21440
rect 12759 21468 12771 21471
rect 14366 21468 14372 21480
rect 12759 21440 14372 21468
rect 12759 21437 12771 21440
rect 12713 21431 12771 21437
rect 14366 21428 14372 21440
rect 14424 21428 14430 21480
rect 15378 21428 15384 21480
rect 15436 21468 15442 21480
rect 15749 21471 15807 21477
rect 15749 21468 15761 21471
rect 15436 21440 15761 21468
rect 15436 21428 15442 21440
rect 15749 21437 15761 21440
rect 15795 21437 15807 21471
rect 16666 21468 16672 21480
rect 16627 21440 16672 21468
rect 15749 21431 15807 21437
rect 16666 21428 16672 21440
rect 16724 21428 16730 21480
rect 16758 21428 16764 21480
rect 16816 21468 16822 21480
rect 20732 21468 20760 21508
rect 31202 21496 31208 21508
rect 31260 21496 31266 21548
rect 16816 21440 20760 21468
rect 20901 21471 20959 21477
rect 16816 21428 16822 21440
rect 20901 21437 20913 21471
rect 20947 21468 20959 21471
rect 23474 21468 23480 21480
rect 20947 21440 23480 21468
rect 20947 21437 20959 21440
rect 20901 21431 20959 21437
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 12158 21400 12164 21412
rect 11992 21372 12164 21400
rect 11517 21363 11575 21369
rect 12158 21360 12164 21372
rect 12216 21360 12222 21412
rect 13081 21403 13139 21409
rect 13081 21369 13093 21403
rect 13127 21400 13139 21403
rect 13170 21400 13176 21412
rect 13127 21372 13176 21400
rect 13127 21369 13139 21372
rect 13081 21363 13139 21369
rect 13170 21360 13176 21372
rect 13228 21360 13234 21412
rect 14292 21372 16160 21400
rect 5316 21304 7052 21332
rect 5316 21292 5322 21304
rect 8202 21292 8208 21344
rect 8260 21332 8266 21344
rect 9723 21335 9781 21341
rect 9723 21332 9735 21335
rect 8260 21304 9735 21332
rect 8260 21292 8266 21304
rect 9723 21301 9735 21304
rect 9769 21301 9781 21335
rect 9723 21295 9781 21301
rect 10226 21292 10232 21344
rect 10284 21332 10290 21344
rect 10781 21335 10839 21341
rect 10781 21332 10793 21335
rect 10284 21304 10793 21332
rect 10284 21292 10290 21304
rect 10781 21301 10793 21304
rect 10827 21301 10839 21335
rect 10781 21295 10839 21301
rect 11974 21292 11980 21344
rect 12032 21332 12038 21344
rect 14292 21332 14320 21372
rect 12032 21304 14320 21332
rect 12032 21292 12038 21304
rect 14366 21292 14372 21344
rect 14424 21332 14430 21344
rect 16132 21332 16160 21372
rect 16206 21360 16212 21412
rect 16264 21400 16270 21412
rect 27798 21400 27804 21412
rect 16264 21372 27804 21400
rect 16264 21360 16270 21372
rect 27798 21360 27804 21372
rect 27856 21360 27862 21412
rect 16942 21332 16948 21344
rect 14424 21304 14469 21332
rect 16132 21304 16948 21332
rect 14424 21292 14430 21304
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 18049 21335 18107 21341
rect 18049 21301 18061 21335
rect 18095 21332 18107 21335
rect 18230 21332 18236 21344
rect 18095 21304 18236 21332
rect 18095 21301 18107 21304
rect 18049 21295 18107 21301
rect 18230 21292 18236 21304
rect 18288 21292 18294 21344
rect 18414 21292 18420 21344
rect 18472 21332 18478 21344
rect 18509 21335 18567 21341
rect 18509 21332 18521 21335
rect 18472 21304 18521 21332
rect 18472 21292 18478 21304
rect 18509 21301 18521 21304
rect 18555 21301 18567 21335
rect 18509 21295 18567 21301
rect 19242 21292 19248 21344
rect 19300 21332 19306 21344
rect 20438 21332 20444 21344
rect 19300 21304 20444 21332
rect 19300 21292 19306 21304
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 21726 21292 21732 21344
rect 21784 21332 21790 21344
rect 21821 21335 21879 21341
rect 21821 21332 21833 21335
rect 21784 21304 21833 21332
rect 21784 21292 21790 21304
rect 21821 21301 21833 21304
rect 21867 21301 21879 21335
rect 21821 21295 21879 21301
rect 22278 21292 22284 21344
rect 22336 21332 22342 21344
rect 22373 21335 22431 21341
rect 22373 21332 22385 21335
rect 22336 21304 22385 21332
rect 22336 21292 22342 21304
rect 22373 21301 22385 21304
rect 22419 21301 22431 21335
rect 23474 21332 23480 21344
rect 23435 21304 23480 21332
rect 22373 21295 22431 21301
rect 23474 21292 23480 21304
rect 23532 21332 23538 21344
rect 23658 21332 23664 21344
rect 23532 21304 23664 21332
rect 23532 21292 23538 21304
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 24118 21332 24124 21344
rect 24079 21304 24124 21332
rect 24118 21292 24124 21304
rect 24176 21292 24182 21344
rect 1104 21242 44896 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 44896 21242
rect 1104 21168 44896 21190
rect 382 21088 388 21140
rect 440 21128 446 21140
rect 2038 21128 2044 21140
rect 440 21100 2044 21128
rect 440 21088 446 21100
rect 2038 21088 2044 21100
rect 2096 21128 2102 21140
rect 3050 21128 3056 21140
rect 2096 21100 3056 21128
rect 2096 21088 2102 21100
rect 3050 21088 3056 21100
rect 3108 21088 3114 21140
rect 3237 21131 3295 21137
rect 3237 21097 3249 21131
rect 3283 21128 3295 21131
rect 3326 21128 3332 21140
rect 3283 21100 3332 21128
rect 3283 21097 3295 21100
rect 3237 21091 3295 21097
rect 3326 21088 3332 21100
rect 3384 21088 3390 21140
rect 4525 21131 4583 21137
rect 4525 21097 4537 21131
rect 4571 21128 4583 21131
rect 4614 21128 4620 21140
rect 4571 21100 4620 21128
rect 4571 21097 4583 21100
rect 4525 21091 4583 21097
rect 4614 21088 4620 21100
rect 4672 21088 4678 21140
rect 5074 21128 5080 21140
rect 4724 21100 5080 21128
rect 1673 21063 1731 21069
rect 1673 21029 1685 21063
rect 1719 21029 1731 21063
rect 1673 21023 1731 21029
rect 2317 21063 2375 21069
rect 2317 21029 2329 21063
rect 2363 21060 2375 21063
rect 3145 21063 3203 21069
rect 2363 21032 3096 21060
rect 2363 21029 2375 21032
rect 2317 21023 2375 21029
rect 1688 20992 1716 21023
rect 3068 20992 3096 21032
rect 3145 21029 3157 21063
rect 3191 21060 3203 21063
rect 4430 21060 4436 21072
rect 3191 21032 4436 21060
rect 3191 21029 3203 21032
rect 3145 21023 3203 21029
rect 4430 21020 4436 21032
rect 4488 21020 4494 21072
rect 4724 20992 4752 21100
rect 5074 21088 5080 21100
rect 5132 21088 5138 21140
rect 8386 21128 8392 21140
rect 8347 21100 8392 21128
rect 8386 21088 8392 21100
rect 8444 21088 8450 21140
rect 8846 21088 8852 21140
rect 8904 21128 8910 21140
rect 10686 21128 10692 21140
rect 8904 21100 10692 21128
rect 8904 21088 8910 21100
rect 10686 21088 10692 21100
rect 10744 21088 10750 21140
rect 11330 21088 11336 21140
rect 11388 21128 11394 21140
rect 12710 21128 12716 21140
rect 11388 21100 12716 21128
rect 11388 21088 11394 21100
rect 12710 21088 12716 21100
rect 12768 21088 12774 21140
rect 13265 21131 13323 21137
rect 13265 21097 13277 21131
rect 13311 21128 13323 21131
rect 13354 21128 13360 21140
rect 13311 21100 13360 21128
rect 13311 21097 13323 21100
rect 13265 21091 13323 21097
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 14366 21088 14372 21140
rect 14424 21128 14430 21140
rect 14424 21100 15792 21128
rect 14424 21088 14430 21100
rect 5718 21060 5724 21072
rect 5000 21032 5724 21060
rect 1688 20964 2774 20992
rect 3068 20964 4752 20992
rect 1489 20927 1547 20933
rect 1489 20893 1501 20927
rect 1535 20924 1547 20927
rect 1946 20924 1952 20936
rect 1535 20896 1952 20924
rect 1535 20893 1547 20896
rect 1489 20887 1547 20893
rect 1946 20884 1952 20896
rect 2004 20884 2010 20936
rect 2130 20924 2136 20936
rect 2091 20896 2136 20924
rect 2130 20884 2136 20896
rect 2188 20884 2194 20936
rect 2746 20924 2774 20964
rect 4798 20952 4804 21004
rect 4856 20992 4862 21004
rect 5000 21001 5028 21032
rect 5718 21020 5724 21032
rect 5776 21020 5782 21072
rect 8018 21020 8024 21072
rect 8076 21060 8082 21072
rect 11606 21060 11612 21072
rect 8076 21032 11612 21060
rect 8076 21020 8082 21032
rect 11606 21020 11612 21032
rect 11664 21020 11670 21072
rect 15654 21060 15660 21072
rect 15615 21032 15660 21060
rect 15654 21020 15660 21032
rect 15712 21020 15718 21072
rect 15764 21060 15792 21100
rect 15838 21088 15844 21140
rect 15896 21128 15902 21140
rect 21358 21128 21364 21140
rect 15896 21100 15941 21128
rect 16408 21100 16712 21128
rect 15896 21088 15902 21100
rect 16408 21060 16436 21100
rect 16574 21060 16580 21072
rect 15764 21032 16436 21060
rect 16535 21032 16580 21060
rect 16574 21020 16580 21032
rect 16632 21020 16638 21072
rect 16684 21060 16712 21100
rect 17328 21100 21364 21128
rect 17328 21060 17356 21100
rect 21358 21088 21364 21100
rect 21416 21088 21422 21140
rect 25225 21131 25283 21137
rect 25225 21097 25237 21131
rect 25271 21128 25283 21131
rect 25314 21128 25320 21140
rect 25271 21100 25320 21128
rect 25271 21097 25283 21100
rect 25225 21091 25283 21097
rect 25314 21088 25320 21100
rect 25372 21088 25378 21140
rect 26602 21128 26608 21140
rect 26563 21100 26608 21128
rect 26602 21088 26608 21100
rect 26660 21088 26666 21140
rect 28074 21128 28080 21140
rect 27540 21100 28080 21128
rect 17494 21060 17500 21072
rect 16684 21032 17356 21060
rect 17455 21032 17500 21060
rect 17494 21020 17500 21032
rect 17552 21020 17558 21072
rect 17681 21063 17739 21069
rect 17681 21029 17693 21063
rect 17727 21060 17739 21063
rect 18046 21060 18052 21072
rect 17727 21032 18052 21060
rect 17727 21029 17739 21032
rect 17681 21023 17739 21029
rect 18046 21020 18052 21032
rect 18104 21020 18110 21072
rect 18141 21063 18199 21069
rect 18141 21029 18153 21063
rect 18187 21060 18199 21063
rect 19794 21060 19800 21072
rect 18187 21032 19800 21060
rect 18187 21029 18199 21032
rect 18141 21023 18199 21029
rect 19794 21020 19800 21032
rect 19852 21020 19858 21072
rect 19996 21032 20392 21060
rect 4985 20995 5043 21001
rect 4856 20964 4936 20992
rect 4856 20952 4862 20964
rect 2746 20896 4844 20924
rect 2777 20859 2835 20865
rect 2777 20825 2789 20859
rect 2823 20856 2835 20859
rect 3050 20856 3056 20868
rect 2823 20828 3056 20856
rect 2823 20825 2835 20828
rect 2777 20819 2835 20825
rect 3050 20816 3056 20828
rect 3108 20816 3114 20868
rect 3789 20859 3847 20865
rect 3789 20856 3801 20859
rect 3160 20828 3801 20856
rect 1302 20748 1308 20800
rect 1360 20788 1366 20800
rect 3160 20788 3188 20828
rect 3789 20825 3801 20828
rect 3835 20825 3847 20859
rect 3789 20819 3847 20825
rect 3973 20859 4031 20865
rect 3973 20825 3985 20859
rect 4019 20856 4031 20859
rect 4338 20856 4344 20868
rect 4019 20828 4344 20856
rect 4019 20825 4031 20828
rect 3973 20819 4031 20825
rect 4338 20816 4344 20828
rect 4396 20816 4402 20868
rect 1360 20760 3188 20788
rect 1360 20748 1366 20760
rect 3878 20748 3884 20800
rect 3936 20788 3942 20800
rect 4706 20788 4712 20800
rect 3936 20760 4712 20788
rect 3936 20748 3942 20760
rect 4706 20748 4712 20760
rect 4764 20748 4770 20800
rect 4816 20788 4844 20896
rect 4908 20865 4936 20964
rect 4985 20961 4997 20995
rect 5031 20961 5043 20995
rect 4985 20955 5043 20961
rect 5169 20995 5227 21001
rect 5169 20961 5181 20995
rect 5215 20992 5227 20995
rect 5442 20992 5448 21004
rect 5215 20964 5448 20992
rect 5215 20961 5227 20964
rect 5169 20955 5227 20961
rect 5442 20952 5448 20964
rect 5500 20952 5506 21004
rect 6273 20995 6331 21001
rect 6273 20961 6285 20995
rect 6319 20992 6331 20995
rect 6362 20992 6368 21004
rect 6319 20964 6368 20992
rect 6319 20961 6331 20964
rect 6273 20955 6331 20961
rect 6362 20952 6368 20964
rect 6420 20952 6426 21004
rect 6454 20952 6460 21004
rect 6512 20992 6518 21004
rect 6638 20992 6644 21004
rect 6512 20964 6644 20992
rect 6512 20952 6518 20964
rect 6638 20952 6644 20964
rect 6696 20952 6702 21004
rect 9306 20992 9312 21004
rect 8036 20964 9312 20992
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 6549 20927 6607 20933
rect 6549 20924 6561 20927
rect 5592 20896 6561 20924
rect 5592 20884 5598 20896
rect 6549 20893 6561 20896
rect 6595 20893 6607 20927
rect 6549 20887 6607 20893
rect 7009 20927 7067 20933
rect 7009 20893 7021 20927
rect 7055 20924 7067 20927
rect 8036 20924 8064 20964
rect 9306 20952 9312 20964
rect 9364 20952 9370 21004
rect 9398 20952 9404 21004
rect 9456 20992 9462 21004
rect 11793 20995 11851 21001
rect 11793 20992 11805 20995
rect 9456 20964 11805 20992
rect 9456 20952 9462 20964
rect 11793 20961 11805 20964
rect 11839 20961 11851 20995
rect 12710 20992 12716 21004
rect 12623 20964 12716 20992
rect 11793 20955 11851 20961
rect 12710 20952 12716 20964
rect 12768 20992 12774 21004
rect 13354 20992 13360 21004
rect 12768 20964 13360 20992
rect 12768 20952 12774 20964
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 14642 20992 14648 21004
rect 14603 20964 14648 20992
rect 14642 20952 14648 20964
rect 14700 20952 14706 21004
rect 14921 20995 14979 21001
rect 14921 20961 14933 20995
rect 14967 20992 14979 20995
rect 16206 20992 16212 21004
rect 14967 20964 16212 20992
rect 14967 20961 14979 20964
rect 14921 20955 14979 20961
rect 16206 20952 16212 20964
rect 16264 20952 16270 21004
rect 16301 20995 16359 21001
rect 16301 20961 16313 20995
rect 16347 20992 16359 20995
rect 16482 20992 16488 21004
rect 16347 20964 16488 20992
rect 16347 20961 16359 20964
rect 16301 20955 16359 20961
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 16758 20992 16764 21004
rect 16719 20964 16764 20992
rect 16758 20952 16764 20964
rect 16816 20952 16822 21004
rect 18506 20952 18512 21004
rect 18564 20992 18570 21004
rect 18874 20992 18880 21004
rect 18564 20964 18880 20992
rect 18564 20952 18570 20964
rect 18874 20952 18880 20964
rect 18932 20992 18938 21004
rect 19996 20992 20024 21032
rect 18932 20964 20024 20992
rect 18932 20952 18938 20964
rect 7055 20896 8064 20924
rect 7055 20893 7067 20896
rect 7009 20887 7067 20893
rect 7944 20868 7972 20896
rect 8294 20884 8300 20936
rect 8352 20924 8358 20936
rect 8941 20927 8999 20933
rect 8941 20924 8953 20927
rect 8352 20896 8953 20924
rect 8352 20884 8358 20896
rect 8941 20893 8953 20896
rect 8987 20893 8999 20927
rect 10778 20924 10784 20936
rect 10739 20896 10784 20924
rect 8941 20887 8999 20893
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 12066 20924 12072 20936
rect 12027 20896 12072 20924
rect 12066 20884 12072 20896
rect 12124 20884 12130 20936
rect 12802 20924 12808 20936
rect 12763 20896 12808 20924
rect 12802 20884 12808 20896
rect 12860 20884 12866 20936
rect 12897 20927 12955 20933
rect 12897 20893 12909 20927
rect 12943 20924 12955 20927
rect 13170 20924 13176 20936
rect 12943 20896 13176 20924
rect 12943 20893 12955 20896
rect 12897 20887 12955 20893
rect 13170 20884 13176 20896
rect 13228 20884 13234 20936
rect 18325 20927 18383 20933
rect 18325 20893 18337 20927
rect 18371 20924 18383 20927
rect 19150 20924 19156 20936
rect 18371 20896 19156 20924
rect 18371 20893 18383 20896
rect 18325 20887 18383 20893
rect 19150 20884 19156 20896
rect 19208 20884 19214 20936
rect 19886 20924 19892 20936
rect 19260 20896 19892 20924
rect 4893 20859 4951 20865
rect 4893 20825 4905 20859
rect 4939 20856 4951 20859
rect 6454 20856 6460 20868
rect 4939 20828 6460 20856
rect 4939 20825 4951 20828
rect 4893 20819 4951 20825
rect 6454 20816 6460 20828
rect 6512 20816 6518 20868
rect 7282 20865 7288 20868
rect 7276 20819 7288 20865
rect 7340 20856 7346 20868
rect 7340 20828 7376 20856
rect 7282 20816 7288 20819
rect 7340 20816 7346 20828
rect 7926 20816 7932 20868
rect 7984 20816 7990 20868
rect 8386 20816 8392 20868
rect 8444 20856 8450 20868
rect 8846 20856 8852 20868
rect 8444 20828 8852 20856
rect 8444 20816 8450 20828
rect 8846 20816 8852 20828
rect 8904 20816 8910 20868
rect 9125 20859 9183 20865
rect 9125 20825 9137 20859
rect 9171 20856 9183 20859
rect 9766 20856 9772 20868
rect 9171 20828 9772 20856
rect 9171 20825 9183 20828
rect 9125 20819 9183 20825
rect 9766 20816 9772 20828
rect 9824 20816 9830 20868
rect 11606 20816 11612 20868
rect 11664 20856 11670 20868
rect 13538 20856 13544 20868
rect 11664 20828 13544 20856
rect 11664 20816 11670 20828
rect 13538 20816 13544 20828
rect 13596 20816 13602 20868
rect 15286 20816 15292 20868
rect 15344 20856 15350 20868
rect 15381 20859 15439 20865
rect 15381 20856 15393 20859
rect 15344 20828 15393 20856
rect 15344 20816 15350 20828
rect 15381 20825 15393 20828
rect 15427 20856 15439 20859
rect 15470 20856 15476 20868
rect 15427 20828 15476 20856
rect 15427 20825 15439 20828
rect 15381 20819 15439 20825
rect 15470 20816 15476 20828
rect 15528 20856 15534 20868
rect 16574 20856 16580 20868
rect 15528 20828 16580 20856
rect 15528 20816 15534 20828
rect 16574 20816 16580 20828
rect 16632 20816 16638 20868
rect 17126 20816 17132 20868
rect 17184 20856 17190 20868
rect 17221 20859 17279 20865
rect 17221 20856 17233 20859
rect 17184 20828 17233 20856
rect 17184 20816 17190 20828
rect 17221 20825 17233 20828
rect 17267 20856 17279 20859
rect 19058 20856 19064 20868
rect 17267 20828 19064 20856
rect 17267 20825 17279 20828
rect 17221 20819 17279 20825
rect 19058 20816 19064 20828
rect 19116 20816 19122 20868
rect 13170 20788 13176 20800
rect 4816 20760 13176 20788
rect 13170 20748 13176 20760
rect 13228 20748 13234 20800
rect 13354 20748 13360 20800
rect 13412 20788 13418 20800
rect 19260 20788 19288 20896
rect 19886 20884 19892 20896
rect 19944 20884 19950 20936
rect 20364 20933 20392 21032
rect 23198 21020 23204 21072
rect 23256 21060 23262 21072
rect 24026 21060 24032 21072
rect 23256 21032 24032 21060
rect 23256 21020 23262 21032
rect 24026 21020 24032 21032
rect 24084 21020 24090 21072
rect 20438 20952 20444 21004
rect 20496 20992 20502 21004
rect 22646 20992 22652 21004
rect 20496 20964 22652 20992
rect 20496 20952 20502 20964
rect 22646 20952 22652 20964
rect 22704 20952 22710 21004
rect 26620 20992 26648 21088
rect 27540 21069 27568 21100
rect 28074 21088 28080 21100
rect 28132 21088 28138 21140
rect 27525 21063 27583 21069
rect 27525 21029 27537 21063
rect 27571 21029 27583 21063
rect 27525 21023 27583 21029
rect 27157 20995 27215 21001
rect 27157 20992 27169 20995
rect 26620 20964 27169 20992
rect 27157 20961 27169 20964
rect 27203 20961 27215 20995
rect 27157 20955 27215 20961
rect 27617 20995 27675 21001
rect 27617 20961 27629 20995
rect 27663 20992 27675 20995
rect 32214 20992 32220 21004
rect 27663 20964 32220 20992
rect 27663 20961 27675 20964
rect 27617 20955 27675 20961
rect 32214 20952 32220 20964
rect 32272 20952 32278 21004
rect 20349 20927 20407 20933
rect 20349 20893 20361 20927
rect 20395 20924 20407 20927
rect 25958 20924 25964 20936
rect 20395 20896 25964 20924
rect 20395 20893 20407 20896
rect 20349 20887 20407 20893
rect 25958 20884 25964 20896
rect 26016 20884 26022 20936
rect 19334 20816 19340 20868
rect 19392 20856 19398 20868
rect 19392 20828 19437 20856
rect 19392 20816 19398 20828
rect 19978 20816 19984 20868
rect 20036 20856 20042 20868
rect 23109 20859 23167 20865
rect 23109 20856 23121 20859
rect 20036 20828 23121 20856
rect 20036 20816 20042 20828
rect 23109 20825 23121 20828
rect 23155 20825 23167 20859
rect 23109 20819 23167 20825
rect 23198 20816 23204 20868
rect 23256 20856 23262 20868
rect 24762 20856 24768 20868
rect 23256 20828 24768 20856
rect 23256 20816 23262 20828
rect 24762 20816 24768 20828
rect 24820 20816 24826 20868
rect 25682 20816 25688 20868
rect 25740 20856 25746 20868
rect 26878 20856 26884 20868
rect 25740 20828 26884 20856
rect 25740 20816 25746 20828
rect 26878 20816 26884 20828
rect 26936 20816 26942 20868
rect 13412 20760 19288 20788
rect 19889 20791 19947 20797
rect 13412 20748 13418 20760
rect 19889 20757 19901 20791
rect 19935 20788 19947 20791
rect 20530 20788 20536 20800
rect 19935 20760 20536 20788
rect 19935 20757 19947 20760
rect 19889 20751 19947 20757
rect 20530 20748 20536 20760
rect 20588 20748 20594 20800
rect 20898 20788 20904 20800
rect 20859 20760 20904 20788
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 21450 20788 21456 20800
rect 21411 20760 21456 20788
rect 21450 20748 21456 20760
rect 21508 20748 21514 20800
rect 22097 20791 22155 20797
rect 22097 20757 22109 20791
rect 22143 20788 22155 20791
rect 22186 20788 22192 20800
rect 22143 20760 22192 20788
rect 22143 20757 22155 20760
rect 22097 20751 22155 20757
rect 22186 20748 22192 20760
rect 22244 20788 22250 20800
rect 22462 20788 22468 20800
rect 22244 20760 22468 20788
rect 22244 20748 22250 20760
rect 22462 20748 22468 20760
rect 22520 20748 22526 20800
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 23290 20788 23296 20800
rect 22704 20760 23296 20788
rect 22704 20748 22710 20760
rect 23290 20748 23296 20760
rect 23348 20748 23354 20800
rect 23658 20788 23664 20800
rect 23619 20760 23664 20788
rect 23658 20748 23664 20760
rect 23716 20748 23722 20800
rect 24486 20788 24492 20800
rect 24447 20760 24492 20788
rect 24486 20748 24492 20760
rect 24544 20748 24550 20800
rect 29086 20748 29092 20800
rect 29144 20788 29150 20800
rect 29549 20791 29607 20797
rect 29549 20788 29561 20791
rect 29144 20760 29561 20788
rect 29144 20748 29150 20760
rect 29549 20757 29561 20760
rect 29595 20757 29607 20791
rect 29549 20751 29607 20757
rect 1104 20698 44896 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 44896 20698
rect 1104 20624 44896 20646
rect 1210 20544 1216 20596
rect 1268 20584 1274 20596
rect 3237 20587 3295 20593
rect 3237 20584 3249 20587
rect 1268 20556 3249 20584
rect 1268 20544 1274 20556
rect 3237 20553 3249 20556
rect 3283 20553 3295 20587
rect 3237 20547 3295 20553
rect 4338 20544 4344 20596
rect 4396 20584 4402 20596
rect 6362 20584 6368 20596
rect 4396 20556 6368 20584
rect 4396 20544 4402 20556
rect 6362 20544 6368 20556
rect 6420 20544 6426 20596
rect 6546 20584 6552 20596
rect 6507 20556 6552 20584
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 6638 20544 6644 20596
rect 6696 20584 6702 20596
rect 7006 20584 7012 20596
rect 6696 20556 7012 20584
rect 6696 20544 6702 20556
rect 7006 20544 7012 20556
rect 7064 20544 7070 20596
rect 7558 20544 7564 20596
rect 7616 20584 7622 20596
rect 9122 20584 9128 20596
rect 7616 20556 9128 20584
rect 7616 20544 7622 20556
rect 9122 20544 9128 20556
rect 9180 20544 9186 20596
rect 9582 20544 9588 20596
rect 9640 20584 9646 20596
rect 11698 20584 11704 20596
rect 9640 20556 11704 20584
rect 9640 20544 9646 20556
rect 11698 20544 11704 20556
rect 11756 20544 11762 20596
rect 14200 20556 17632 20584
rect 2133 20519 2191 20525
rect 2133 20485 2145 20519
rect 2179 20516 2191 20519
rect 11514 20516 11520 20528
rect 2179 20488 11520 20516
rect 2179 20485 2191 20488
rect 2133 20479 2191 20485
rect 11514 20476 11520 20488
rect 11572 20476 11578 20528
rect 14200 20516 14228 20556
rect 11624 20488 14228 20516
rect 15657 20519 15715 20525
rect 1397 20451 1455 20457
rect 1397 20417 1409 20451
rect 1443 20448 1455 20451
rect 2314 20448 2320 20460
rect 1443 20420 2320 20448
rect 1443 20417 1455 20420
rect 1397 20411 1455 20417
rect 2314 20408 2320 20420
rect 2372 20448 2378 20460
rect 2498 20448 2504 20460
rect 2372 20420 2504 20448
rect 2372 20408 2378 20420
rect 2498 20408 2504 20420
rect 2556 20408 2562 20460
rect 2590 20408 2596 20460
rect 2648 20448 2654 20460
rect 3602 20448 3608 20460
rect 2648 20420 3608 20448
rect 2648 20408 2654 20420
rect 3602 20408 3608 20420
rect 3660 20408 3666 20460
rect 4246 20448 4252 20460
rect 4207 20420 4252 20448
rect 4246 20408 4252 20420
rect 4304 20408 4310 20460
rect 5166 20448 5172 20460
rect 4356 20420 5172 20448
rect 2038 20340 2044 20392
rect 2096 20380 2102 20392
rect 2777 20383 2835 20389
rect 2777 20380 2789 20383
rect 2096 20352 2789 20380
rect 2096 20340 2102 20352
rect 2777 20349 2789 20352
rect 2823 20380 2835 20383
rect 4356 20380 4384 20420
rect 5166 20408 5172 20420
rect 5224 20408 5230 20460
rect 5534 20448 5540 20460
rect 5495 20420 5540 20448
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 5810 20448 5816 20460
rect 5771 20420 5816 20448
rect 5810 20408 5816 20420
rect 5868 20408 5874 20460
rect 6638 20448 6644 20460
rect 6599 20420 6644 20448
rect 6638 20408 6644 20420
rect 6696 20408 6702 20460
rect 6748 20420 7328 20448
rect 4522 20380 4528 20392
rect 2823 20352 4384 20380
rect 4483 20352 4528 20380
rect 2823 20349 2835 20352
rect 2777 20343 2835 20349
rect 4522 20340 4528 20352
rect 4580 20340 4586 20392
rect 6178 20340 6184 20392
rect 6236 20380 6242 20392
rect 6748 20380 6776 20420
rect 6236 20352 6776 20380
rect 7193 20383 7251 20389
rect 6236 20340 6242 20352
rect 7193 20349 7205 20383
rect 7239 20349 7251 20383
rect 7193 20343 7251 20349
rect 2314 20312 2320 20324
rect 2275 20284 2320 20312
rect 2314 20272 2320 20284
rect 2372 20272 2378 20324
rect 3142 20312 3148 20324
rect 3103 20284 3148 20312
rect 3142 20272 3148 20284
rect 3200 20272 3206 20324
rect 3418 20272 3424 20324
rect 3476 20312 3482 20324
rect 7208 20312 7236 20343
rect 3476 20284 7236 20312
rect 7300 20312 7328 20420
rect 9122 20408 9128 20460
rect 9180 20448 9186 20460
rect 9306 20448 9312 20460
rect 9180 20420 9312 20448
rect 9180 20408 9186 20420
rect 9306 20408 9312 20420
rect 9364 20448 9370 20460
rect 9766 20448 9772 20460
rect 9364 20420 9674 20448
rect 9727 20420 9772 20448
rect 9364 20408 9370 20420
rect 8846 20380 8852 20392
rect 8807 20352 8852 20380
rect 8846 20340 8852 20352
rect 8904 20340 8910 20392
rect 9033 20383 9091 20389
rect 9033 20349 9045 20383
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 9493 20383 9551 20389
rect 9493 20349 9505 20383
rect 9539 20349 9551 20383
rect 9493 20343 9551 20349
rect 9048 20312 9076 20343
rect 7300 20284 9076 20312
rect 3476 20272 3482 20284
rect 1581 20247 1639 20253
rect 1581 20213 1593 20247
rect 1627 20244 1639 20247
rect 2682 20244 2688 20256
rect 1627 20216 2688 20244
rect 1627 20213 1639 20216
rect 1581 20207 1639 20213
rect 2682 20204 2688 20216
rect 2740 20244 2746 20256
rect 3050 20244 3056 20256
rect 2740 20216 3056 20244
rect 2740 20204 2746 20216
rect 3050 20204 3056 20216
rect 3108 20204 3114 20256
rect 4798 20204 4804 20256
rect 4856 20244 4862 20256
rect 9508 20244 9536 20343
rect 9646 20312 9674 20420
rect 9766 20408 9772 20420
rect 9824 20408 9830 20460
rect 10686 20408 10692 20460
rect 10744 20448 10750 20460
rect 10965 20451 11023 20457
rect 10965 20448 10977 20451
rect 10744 20420 10977 20448
rect 10744 20408 10750 20420
rect 10965 20417 10977 20420
rect 11011 20417 11023 20451
rect 11624 20448 11652 20488
rect 15657 20485 15669 20519
rect 15703 20516 15715 20519
rect 16022 20516 16028 20528
rect 15703 20488 16028 20516
rect 15703 20485 15715 20488
rect 15657 20479 15715 20485
rect 16022 20476 16028 20488
rect 16080 20476 16086 20528
rect 17604 20525 17632 20556
rect 18046 20544 18052 20596
rect 18104 20584 18110 20596
rect 18966 20584 18972 20596
rect 18104 20556 18644 20584
rect 18927 20556 18972 20584
rect 18104 20544 18110 20556
rect 17589 20519 17647 20525
rect 17589 20485 17601 20519
rect 17635 20516 17647 20519
rect 18322 20516 18328 20528
rect 17635 20488 18328 20516
rect 17635 20485 17647 20488
rect 17589 20479 17647 20485
rect 18322 20476 18328 20488
rect 18380 20476 18386 20528
rect 18506 20516 18512 20528
rect 18467 20488 18512 20516
rect 18506 20476 18512 20488
rect 18564 20476 18570 20528
rect 18616 20516 18644 20556
rect 18966 20544 18972 20556
rect 19024 20544 19030 20596
rect 20438 20584 20444 20596
rect 20399 20556 20444 20584
rect 20438 20544 20444 20556
rect 20496 20544 20502 20596
rect 20806 20544 20812 20596
rect 20864 20584 20870 20596
rect 20993 20587 21051 20593
rect 20993 20584 21005 20587
rect 20864 20556 21005 20584
rect 20864 20544 20870 20556
rect 20993 20553 21005 20556
rect 21039 20553 21051 20587
rect 22646 20584 22652 20596
rect 22607 20556 22652 20584
rect 20993 20547 21051 20553
rect 22646 20544 22652 20556
rect 22704 20544 22710 20596
rect 24210 20584 24216 20596
rect 24171 20556 24216 20584
rect 24210 20544 24216 20556
rect 24268 20544 24274 20596
rect 25774 20584 25780 20596
rect 25735 20556 25780 20584
rect 25774 20544 25780 20556
rect 25832 20544 25838 20596
rect 28350 20584 28356 20596
rect 28311 20556 28356 20584
rect 28350 20544 28356 20556
rect 28408 20544 28414 20596
rect 29730 20584 29736 20596
rect 29691 20556 29736 20584
rect 29730 20544 29736 20556
rect 29788 20544 29794 20596
rect 19429 20519 19487 20525
rect 19429 20516 19441 20519
rect 18616 20488 19441 20516
rect 19429 20485 19441 20488
rect 19475 20485 19487 20519
rect 19429 20479 19487 20485
rect 22741 20519 22799 20525
rect 22741 20485 22753 20519
rect 22787 20516 22799 20519
rect 24486 20516 24492 20528
rect 22787 20488 24492 20516
rect 22787 20485 22799 20488
rect 22741 20479 22799 20485
rect 24486 20476 24492 20488
rect 24544 20476 24550 20528
rect 24949 20519 25007 20525
rect 24949 20485 24961 20519
rect 24995 20516 25007 20519
rect 25314 20516 25320 20528
rect 24995 20488 25320 20516
rect 24995 20485 25007 20488
rect 24949 20479 25007 20485
rect 25314 20476 25320 20488
rect 25372 20476 25378 20528
rect 27525 20519 27583 20525
rect 27525 20485 27537 20519
rect 27571 20516 27583 20519
rect 27706 20516 27712 20528
rect 27571 20488 27712 20516
rect 27571 20485 27583 20488
rect 27525 20479 27583 20485
rect 27706 20476 27712 20488
rect 27764 20476 27770 20528
rect 10965 20411 11023 20417
rect 11072 20420 11652 20448
rect 10410 20340 10416 20392
rect 10468 20380 10474 20392
rect 11072 20380 11100 20420
rect 12986 20408 12992 20460
rect 13044 20448 13050 20460
rect 13449 20451 13507 20457
rect 13449 20448 13461 20451
rect 13044 20420 13461 20448
rect 13044 20408 13050 20420
rect 13449 20417 13461 20420
rect 13495 20417 13507 20451
rect 13449 20411 13507 20417
rect 13814 20408 13820 20460
rect 13872 20448 13878 20460
rect 14826 20448 14832 20460
rect 13872 20420 14832 20448
rect 13872 20408 13878 20420
rect 14826 20408 14832 20420
rect 14884 20408 14890 20460
rect 14921 20451 14979 20457
rect 14921 20417 14933 20451
rect 14967 20448 14979 20451
rect 15010 20448 15016 20460
rect 14967 20420 15016 20448
rect 14967 20417 14979 20420
rect 14921 20411 14979 20417
rect 15010 20408 15016 20420
rect 15068 20408 15074 20460
rect 18138 20448 18144 20460
rect 15948 20420 18144 20448
rect 10468 20352 11100 20380
rect 10468 20340 10474 20352
rect 11146 20340 11152 20392
rect 11204 20380 11210 20392
rect 12069 20383 12127 20389
rect 12069 20380 12081 20383
rect 11204 20352 12081 20380
rect 11204 20340 11210 20352
rect 12069 20349 12081 20352
rect 12115 20349 12127 20383
rect 12069 20343 12127 20349
rect 12345 20383 12403 20389
rect 12345 20349 12357 20383
rect 12391 20380 12403 20383
rect 13538 20380 13544 20392
rect 12391 20352 13544 20380
rect 12391 20349 12403 20352
rect 12345 20343 12403 20349
rect 13538 20340 13544 20352
rect 13596 20340 13602 20392
rect 13630 20340 13636 20392
rect 13688 20380 13694 20392
rect 13725 20383 13783 20389
rect 13725 20380 13737 20383
rect 13688 20352 13737 20380
rect 13688 20340 13694 20352
rect 13725 20349 13737 20352
rect 13771 20349 13783 20383
rect 13725 20343 13783 20349
rect 14642 20340 14648 20392
rect 14700 20380 14706 20392
rect 15197 20383 15255 20389
rect 15197 20380 15209 20383
rect 14700 20352 15209 20380
rect 14700 20340 14706 20352
rect 15197 20349 15209 20352
rect 15243 20349 15255 20383
rect 15197 20343 15255 20349
rect 10781 20315 10839 20321
rect 10781 20312 10793 20315
rect 9646 20284 10793 20312
rect 10781 20281 10793 20284
rect 10827 20312 10839 20315
rect 15948 20312 15976 20420
rect 18138 20408 18144 20420
rect 18196 20408 18202 20460
rect 20898 20448 20904 20460
rect 18248 20420 20904 20448
rect 16114 20380 16120 20392
rect 16040 20352 16120 20380
rect 16040 20321 16068 20352
rect 16114 20340 16120 20352
rect 16172 20340 16178 20392
rect 17218 20340 17224 20392
rect 17276 20380 17282 20392
rect 17494 20380 17500 20392
rect 17276 20352 17500 20380
rect 17276 20340 17282 20352
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 10827 20284 15976 20312
rect 16025 20315 16083 20321
rect 10827 20281 10839 20284
rect 10781 20275 10839 20281
rect 16025 20281 16037 20315
rect 16071 20281 16083 20315
rect 16025 20275 16083 20281
rect 17313 20315 17371 20321
rect 17313 20281 17325 20315
rect 17359 20312 17371 20315
rect 17954 20312 17960 20324
rect 17359 20284 17960 20312
rect 17359 20281 17371 20284
rect 17313 20275 17371 20281
rect 17954 20272 17960 20284
rect 18012 20272 18018 20324
rect 18248 20321 18276 20420
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 24118 20448 24124 20460
rect 24031 20420 24124 20448
rect 24118 20408 24124 20420
rect 24176 20408 24182 20460
rect 25685 20451 25743 20457
rect 25685 20417 25697 20451
rect 25731 20448 25743 20451
rect 25774 20448 25780 20460
rect 25731 20420 25780 20448
rect 25731 20417 25743 20420
rect 25685 20411 25743 20417
rect 25774 20408 25780 20420
rect 25832 20408 25838 20460
rect 27246 20408 27252 20460
rect 27304 20448 27310 20460
rect 28905 20451 28963 20457
rect 28905 20448 28917 20451
rect 27304 20420 28917 20448
rect 27304 20408 27310 20420
rect 28905 20417 28917 20420
rect 28951 20417 28963 20451
rect 29086 20448 29092 20460
rect 29047 20420 29092 20448
rect 28905 20411 28963 20417
rect 29086 20408 29092 20420
rect 29144 20408 29150 20460
rect 19518 20340 19524 20392
rect 19576 20380 19582 20392
rect 21634 20380 21640 20392
rect 19576 20352 21640 20380
rect 19576 20340 19582 20352
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 24136 20380 24164 20408
rect 33594 20380 33600 20392
rect 24136 20352 33600 20380
rect 33594 20340 33600 20352
rect 33652 20340 33658 20392
rect 18233 20315 18291 20321
rect 18233 20281 18245 20315
rect 18279 20281 18291 20315
rect 18233 20275 18291 20281
rect 19153 20315 19211 20321
rect 19153 20281 19165 20315
rect 19199 20312 19211 20315
rect 21821 20315 21879 20321
rect 21821 20312 21833 20315
rect 19199 20284 21833 20312
rect 19199 20281 19211 20284
rect 19153 20275 19211 20281
rect 21821 20281 21833 20284
rect 21867 20312 21879 20315
rect 21910 20312 21916 20324
rect 21867 20284 21916 20312
rect 21867 20281 21879 20284
rect 21821 20275 21879 20281
rect 21910 20272 21916 20284
rect 21968 20272 21974 20324
rect 4856 20216 9536 20244
rect 16117 20247 16175 20253
rect 4856 20204 4862 20216
rect 16117 20213 16129 20247
rect 16163 20244 16175 20247
rect 16482 20244 16488 20256
rect 16163 20216 16488 20244
rect 16163 20213 16175 20216
rect 16117 20207 16175 20213
rect 16482 20204 16488 20216
rect 16540 20204 16546 20256
rect 17126 20244 17132 20256
rect 17087 20216 17132 20244
rect 17126 20204 17132 20216
rect 17184 20204 17190 20256
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 18049 20247 18107 20253
rect 18049 20244 18061 20247
rect 17276 20216 18061 20244
rect 17276 20204 17282 20216
rect 18049 20213 18061 20216
rect 18095 20213 18107 20247
rect 18049 20207 18107 20213
rect 18690 20204 18696 20256
rect 18748 20244 18754 20256
rect 19889 20247 19947 20253
rect 19889 20244 19901 20247
rect 18748 20216 19901 20244
rect 18748 20204 18754 20216
rect 19889 20213 19901 20216
rect 19935 20213 19947 20247
rect 19889 20207 19947 20213
rect 20898 20204 20904 20256
rect 20956 20244 20962 20256
rect 23293 20247 23351 20253
rect 23293 20244 23305 20247
rect 20956 20216 23305 20244
rect 20956 20204 20962 20216
rect 23293 20213 23305 20216
rect 23339 20213 23351 20247
rect 24854 20244 24860 20256
rect 24815 20216 24860 20244
rect 23293 20207 23351 20213
rect 24854 20204 24860 20216
rect 24912 20204 24918 20256
rect 27430 20244 27436 20256
rect 27391 20216 27436 20244
rect 27430 20204 27436 20216
rect 27488 20204 27494 20256
rect 33597 20247 33655 20253
rect 33597 20213 33609 20247
rect 33643 20244 33655 20247
rect 33778 20244 33784 20256
rect 33643 20216 33784 20244
rect 33643 20213 33655 20216
rect 33597 20207 33655 20213
rect 33778 20204 33784 20216
rect 33836 20204 33842 20256
rect 1104 20154 44896 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 44896 20154
rect 1104 20080 44896 20102
rect 2041 20043 2099 20049
rect 2041 20009 2053 20043
rect 2087 20040 2099 20043
rect 2130 20040 2136 20052
rect 2087 20012 2136 20040
rect 2087 20009 2099 20012
rect 2041 20003 2099 20009
rect 2130 20000 2136 20012
rect 2188 20000 2194 20052
rect 3234 20040 3240 20052
rect 3195 20012 3240 20040
rect 3234 20000 3240 20012
rect 3292 20000 3298 20052
rect 4706 20000 4712 20052
rect 4764 20040 4770 20052
rect 5166 20040 5172 20052
rect 4764 20012 5172 20040
rect 4764 20000 4770 20012
rect 5166 20000 5172 20012
rect 5224 20000 5230 20052
rect 6638 20000 6644 20052
rect 6696 20040 6702 20052
rect 9674 20040 9680 20052
rect 6696 20012 9680 20040
rect 6696 20000 6702 20012
rect 9674 20000 9680 20012
rect 9732 20040 9738 20052
rect 10686 20040 10692 20052
rect 9732 20012 10692 20040
rect 9732 20000 9738 20012
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 18138 20000 18144 20052
rect 18196 20040 18202 20052
rect 18414 20040 18420 20052
rect 18196 20012 18420 20040
rect 18196 20000 18202 20012
rect 18414 20000 18420 20012
rect 18472 20040 18478 20052
rect 18693 20043 18751 20049
rect 18693 20040 18705 20043
rect 18472 20012 18705 20040
rect 18472 20000 18478 20012
rect 18693 20009 18705 20012
rect 18739 20009 18751 20043
rect 18693 20003 18751 20009
rect 18966 20000 18972 20052
rect 19024 20040 19030 20052
rect 19150 20040 19156 20052
rect 19024 20012 19156 20040
rect 19024 20000 19030 20012
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 20438 20000 20444 20052
rect 20496 20040 20502 20052
rect 22186 20040 22192 20052
rect 20496 20012 22192 20040
rect 20496 20000 20502 20012
rect 22186 20000 22192 20012
rect 22244 20000 22250 20052
rect 25590 20000 25596 20052
rect 25648 20040 25654 20052
rect 25685 20043 25743 20049
rect 25685 20040 25697 20043
rect 25648 20012 25697 20040
rect 25648 20000 25654 20012
rect 25685 20009 25697 20012
rect 25731 20009 25743 20043
rect 28166 20040 28172 20052
rect 25685 20003 25743 20009
rect 25792 20012 28172 20040
rect 1946 19972 1952 19984
rect 1907 19944 1952 19972
rect 1946 19932 1952 19944
rect 2004 19932 2010 19984
rect 2498 19932 2504 19984
rect 2556 19972 2562 19984
rect 6178 19972 6184 19984
rect 2556 19944 6184 19972
rect 2556 19932 2562 19944
rect 6178 19932 6184 19944
rect 6236 19932 6242 19984
rect 6362 19932 6368 19984
rect 6420 19972 6426 19984
rect 6420 19944 7420 19972
rect 6420 19932 6426 19944
rect 1581 19907 1639 19913
rect 1581 19873 1593 19907
rect 1627 19904 1639 19907
rect 2038 19904 2044 19916
rect 1627 19876 2044 19904
rect 1627 19873 1639 19876
rect 1581 19867 1639 19873
rect 2038 19864 2044 19876
rect 2096 19864 2102 19916
rect 2685 19907 2743 19913
rect 2685 19873 2697 19907
rect 2731 19904 2743 19907
rect 2866 19904 2872 19916
rect 2731 19876 2872 19904
rect 2731 19873 2743 19876
rect 2685 19867 2743 19873
rect 2866 19864 2872 19876
rect 2924 19904 2930 19916
rect 3786 19904 3792 19916
rect 2924 19876 3792 19904
rect 2924 19864 2930 19876
rect 3786 19864 3792 19876
rect 3844 19864 3850 19916
rect 4525 19907 4583 19913
rect 4525 19873 4537 19907
rect 4571 19904 4583 19907
rect 4890 19904 4896 19916
rect 4571 19876 4896 19904
rect 4571 19873 4583 19876
rect 4525 19867 4583 19873
rect 4890 19864 4896 19876
rect 4948 19864 4954 19916
rect 5813 19907 5871 19913
rect 5276 19876 5764 19904
rect 3326 19836 3332 19848
rect 2056 19808 3332 19836
rect 2056 19780 2084 19808
rect 3326 19796 3332 19808
rect 3384 19796 3390 19848
rect 4706 19796 4712 19848
rect 4764 19836 4770 19848
rect 4801 19839 4859 19845
rect 4801 19836 4813 19839
rect 4764 19808 4813 19836
rect 4764 19796 4770 19808
rect 4801 19805 4813 19808
rect 4847 19805 4859 19839
rect 4801 19799 4859 19805
rect 2038 19728 2044 19780
rect 2096 19728 2102 19780
rect 2777 19771 2835 19777
rect 2777 19737 2789 19771
rect 2823 19768 2835 19771
rect 5276 19768 5304 19876
rect 5350 19796 5356 19848
rect 5408 19796 5414 19848
rect 2823 19740 5304 19768
rect 2823 19737 2835 19740
rect 2777 19731 2835 19737
rect 2869 19703 2927 19709
rect 2869 19669 2881 19703
rect 2915 19700 2927 19703
rect 3326 19700 3332 19712
rect 2915 19672 3332 19700
rect 2915 19669 2927 19672
rect 2869 19663 2927 19669
rect 3326 19660 3332 19672
rect 3384 19660 3390 19712
rect 4154 19660 4160 19712
rect 4212 19700 4218 19712
rect 5368 19700 5396 19796
rect 5736 19768 5764 19876
rect 5813 19873 5825 19907
rect 5859 19904 5871 19907
rect 6730 19904 6736 19916
rect 5859 19876 6736 19904
rect 5859 19873 5871 19876
rect 5813 19867 5871 19873
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 7282 19904 7288 19916
rect 7243 19876 7288 19904
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 7392 19904 7420 19944
rect 8846 19932 8852 19984
rect 8904 19972 8910 19984
rect 16758 19972 16764 19984
rect 8904 19944 16764 19972
rect 8904 19932 8910 19944
rect 16758 19932 16764 19944
rect 16816 19932 16822 19984
rect 16945 19975 17003 19981
rect 16945 19941 16957 19975
rect 16991 19972 17003 19975
rect 17402 19972 17408 19984
rect 16991 19944 17408 19972
rect 16991 19941 17003 19944
rect 16945 19935 17003 19941
rect 17402 19932 17408 19944
rect 17460 19932 17466 19984
rect 17862 19932 17868 19984
rect 17920 19972 17926 19984
rect 17957 19975 18015 19981
rect 17957 19972 17969 19975
rect 17920 19944 17969 19972
rect 17920 19932 17926 19944
rect 17957 19941 17969 19944
rect 18003 19941 18015 19975
rect 17957 19935 18015 19941
rect 19889 19975 19947 19981
rect 19889 19941 19901 19975
rect 19935 19972 19947 19975
rect 25792 19972 25820 20012
rect 28166 20000 28172 20012
rect 28224 20000 28230 20052
rect 32766 20040 32772 20052
rect 32727 20012 32772 20040
rect 32766 20000 32772 20012
rect 32824 20000 32830 20052
rect 37826 20040 37832 20052
rect 35866 20012 37832 20040
rect 19935 19944 21128 19972
rect 19935 19941 19947 19944
rect 19889 19935 19947 19941
rect 9398 19904 9404 19916
rect 7392 19876 9404 19904
rect 9398 19864 9404 19876
rect 9456 19864 9462 19916
rect 10781 19907 10839 19913
rect 10781 19873 10793 19907
rect 10827 19904 10839 19907
rect 11054 19904 11060 19916
rect 10827 19876 11060 19904
rect 10827 19873 10839 19876
rect 10781 19867 10839 19873
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 11790 19904 11796 19916
rect 11751 19876 11796 19904
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 13262 19904 13268 19916
rect 13223 19876 13268 19904
rect 13262 19864 13268 19876
rect 13320 19864 13326 19916
rect 14366 19904 14372 19916
rect 14327 19876 14372 19904
rect 14366 19864 14372 19876
rect 14424 19864 14430 19916
rect 15102 19864 15108 19916
rect 15160 19904 15166 19916
rect 15933 19907 15991 19913
rect 15933 19904 15945 19907
rect 15160 19876 15945 19904
rect 15160 19864 15166 19876
rect 15933 19873 15945 19876
rect 15979 19873 15991 19907
rect 16206 19904 16212 19916
rect 16167 19876 16212 19904
rect 15933 19867 15991 19873
rect 16206 19864 16212 19876
rect 16264 19864 16270 19916
rect 16482 19864 16488 19916
rect 16540 19904 16546 19916
rect 18230 19904 18236 19916
rect 16540 19876 18236 19904
rect 16540 19864 16546 19876
rect 18230 19864 18236 19876
rect 18288 19904 18294 19916
rect 20901 19907 20959 19913
rect 18288 19876 18644 19904
rect 18288 19864 18294 19876
rect 18616 19848 18644 19876
rect 20901 19873 20913 19907
rect 20947 19904 20959 19907
rect 20990 19904 20996 19916
rect 20947 19876 20996 19904
rect 20947 19873 20959 19876
rect 20901 19867 20959 19873
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 21100 19904 21128 19944
rect 22066 19944 25820 19972
rect 27065 19975 27123 19981
rect 22066 19904 22094 19944
rect 27065 19941 27077 19975
rect 27111 19972 27123 19975
rect 27154 19972 27160 19984
rect 27111 19944 27160 19972
rect 27111 19941 27123 19944
rect 27065 19935 27123 19941
rect 27154 19932 27160 19944
rect 27212 19932 27218 19984
rect 28442 19932 28448 19984
rect 28500 19972 28506 19984
rect 28810 19972 28816 19984
rect 28500 19944 28816 19972
rect 28500 19932 28506 19944
rect 28810 19932 28816 19944
rect 28868 19932 28874 19984
rect 30650 19972 30656 19984
rect 30611 19944 30656 19972
rect 30650 19932 30656 19944
rect 30708 19932 30714 19984
rect 35866 19972 35894 20012
rect 37826 20000 37832 20012
rect 37884 20000 37890 20052
rect 31772 19944 35894 19972
rect 36081 19975 36139 19981
rect 21100 19876 22094 19904
rect 22189 19907 22247 19913
rect 22189 19873 22201 19907
rect 22235 19904 22247 19907
rect 22830 19904 22836 19916
rect 22235 19876 22836 19904
rect 22235 19873 22247 19876
rect 22189 19867 22247 19873
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 27801 19907 27859 19913
rect 27801 19873 27813 19907
rect 27847 19904 27859 19907
rect 31772 19904 31800 19944
rect 36081 19941 36093 19975
rect 36127 19972 36139 19975
rect 43622 19972 43628 19984
rect 36127 19944 43628 19972
rect 36127 19941 36139 19944
rect 36081 19935 36139 19941
rect 43622 19932 43628 19944
rect 43680 19932 43686 19984
rect 27847 19876 31800 19904
rect 35345 19907 35403 19913
rect 27847 19873 27859 19876
rect 27801 19867 27859 19873
rect 35345 19873 35357 19907
rect 35391 19904 35403 19907
rect 43530 19904 43536 19916
rect 35391 19876 43536 19904
rect 35391 19873 35403 19876
rect 35345 19867 35403 19873
rect 43530 19864 43536 19876
rect 43588 19864 43594 19916
rect 6086 19836 6092 19848
rect 6047 19808 6092 19836
rect 6086 19796 6092 19808
rect 6144 19796 6150 19848
rect 6362 19796 6368 19848
rect 6420 19836 6426 19848
rect 6549 19839 6607 19845
rect 6549 19836 6561 19839
rect 6420 19808 6561 19836
rect 6420 19796 6426 19808
rect 6549 19805 6561 19808
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 8846 19796 8852 19848
rect 8904 19836 8910 19848
rect 8941 19839 8999 19845
rect 8941 19836 8953 19839
rect 8904 19808 8953 19836
rect 8904 19796 8910 19808
rect 8941 19805 8953 19808
rect 8987 19805 8999 19839
rect 8941 19799 8999 19805
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19836 12127 19839
rect 12342 19836 12348 19848
rect 12115 19808 12348 19836
rect 12115 19805 12127 19808
rect 12069 19799 12127 19805
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 13538 19836 13544 19848
rect 13499 19808 13544 19836
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 14090 19836 14096 19848
rect 14051 19808 14096 19836
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14826 19796 14832 19848
rect 14884 19836 14890 19848
rect 14884 19808 17816 19836
rect 14884 19796 14890 19808
rect 5810 19768 5816 19780
rect 5736 19740 5816 19768
rect 5810 19728 5816 19740
rect 5868 19728 5874 19780
rect 6730 19768 6736 19780
rect 6691 19740 6736 19768
rect 6730 19728 6736 19740
rect 6788 19728 6794 19780
rect 9122 19768 9128 19780
rect 9083 19740 9128 19768
rect 9122 19728 9128 19740
rect 9180 19728 9186 19780
rect 16206 19728 16212 19780
rect 16264 19768 16270 19780
rect 16850 19768 16856 19780
rect 16264 19740 16856 19768
rect 16264 19728 16270 19740
rect 16850 19728 16856 19740
rect 16908 19768 16914 19780
rect 17221 19771 17279 19777
rect 16908 19740 17172 19768
rect 16908 19728 16914 19740
rect 4212 19672 5396 19700
rect 4212 19660 4218 19672
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 7098 19700 7104 19712
rect 5592 19672 7104 19700
rect 5592 19660 5598 19672
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 7190 19660 7196 19712
rect 7248 19700 7254 19712
rect 8754 19700 8760 19712
rect 7248 19672 8760 19700
rect 7248 19660 7254 19672
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 13538 19660 13544 19712
rect 13596 19700 13602 19712
rect 16574 19700 16580 19712
rect 13596 19672 16580 19700
rect 13596 19660 13602 19672
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 16666 19660 16672 19712
rect 16724 19700 16730 19712
rect 16761 19703 16819 19709
rect 16761 19700 16773 19703
rect 16724 19672 16773 19700
rect 16724 19660 16730 19672
rect 16761 19669 16773 19672
rect 16807 19669 16819 19703
rect 17144 19700 17172 19740
rect 17221 19737 17233 19771
rect 17267 19768 17279 19771
rect 17494 19768 17500 19780
rect 17267 19740 17500 19768
rect 17267 19737 17279 19740
rect 17221 19731 17279 19737
rect 17494 19728 17500 19740
rect 17552 19728 17558 19780
rect 17681 19771 17739 19777
rect 17681 19737 17693 19771
rect 17727 19737 17739 19771
rect 17788 19768 17816 19808
rect 18598 19796 18604 19848
rect 18656 19796 18662 19848
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19836 19763 19839
rect 20162 19836 20168 19848
rect 19751 19808 20168 19836
rect 19751 19805 19763 19808
rect 19705 19799 19763 19805
rect 20162 19796 20168 19808
rect 20220 19796 20226 19848
rect 20622 19836 20628 19848
rect 20583 19808 20628 19836
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 21266 19796 21272 19848
rect 21324 19836 21330 19848
rect 21913 19839 21971 19845
rect 21913 19836 21925 19839
rect 21324 19808 21925 19836
rect 21324 19796 21330 19808
rect 21913 19805 21925 19808
rect 21959 19805 21971 19839
rect 21913 19799 21971 19805
rect 23293 19839 23351 19845
rect 23293 19805 23305 19839
rect 23339 19836 23351 19839
rect 23382 19836 23388 19848
rect 23339 19808 23388 19836
rect 23339 19805 23351 19808
rect 23293 19799 23351 19805
rect 23382 19796 23388 19808
rect 23440 19796 23446 19848
rect 24857 19839 24915 19845
rect 24857 19805 24869 19839
rect 24903 19836 24915 19839
rect 24946 19836 24952 19848
rect 24903 19808 24952 19836
rect 24903 19805 24915 19808
rect 24857 19799 24915 19805
rect 24946 19796 24952 19808
rect 25004 19836 25010 19848
rect 26237 19839 26295 19845
rect 26237 19836 26249 19839
rect 25004 19808 26249 19836
rect 25004 19796 25010 19808
rect 26237 19805 26249 19808
rect 26283 19805 26295 19839
rect 26237 19799 26295 19805
rect 28350 19796 28356 19848
rect 28408 19836 28414 19848
rect 28537 19839 28595 19845
rect 28537 19836 28549 19839
rect 28408 19808 28549 19836
rect 28408 19796 28414 19808
rect 28537 19805 28549 19808
rect 28583 19805 28595 19839
rect 28537 19799 28595 19805
rect 29730 19796 29736 19848
rect 29788 19836 29794 19848
rect 30009 19839 30067 19845
rect 30009 19836 30021 19839
rect 29788 19808 30021 19836
rect 29788 19796 29794 19808
rect 30009 19805 30021 19808
rect 30055 19805 30067 19839
rect 33410 19836 33416 19848
rect 30009 19799 30067 19805
rect 30300 19808 33416 19836
rect 21542 19768 21548 19780
rect 17788 19740 21548 19768
rect 17681 19731 17739 19737
rect 17696 19700 17724 19731
rect 21542 19728 21548 19740
rect 21600 19728 21606 19780
rect 23474 19768 23480 19780
rect 23435 19740 23480 19768
rect 23474 19728 23480 19740
rect 23532 19728 23538 19780
rect 25038 19768 25044 19780
rect 24999 19740 25044 19768
rect 25038 19728 25044 19740
rect 25096 19728 25102 19780
rect 25593 19771 25651 19777
rect 25593 19737 25605 19771
rect 25639 19737 25651 19771
rect 26878 19768 26884 19780
rect 26839 19740 26884 19768
rect 25593 19731 25651 19737
rect 18138 19700 18144 19712
rect 17144 19672 17724 19700
rect 18099 19672 18144 19700
rect 16761 19663 16819 19669
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 18322 19660 18328 19712
rect 18380 19700 18386 19712
rect 21174 19700 21180 19712
rect 18380 19672 21180 19700
rect 18380 19660 18386 19672
rect 21174 19660 21180 19672
rect 21232 19660 21238 19712
rect 21634 19660 21640 19712
rect 21692 19700 21698 19712
rect 24762 19700 24768 19712
rect 21692 19672 24768 19700
rect 21692 19660 21698 19672
rect 24762 19660 24768 19672
rect 24820 19660 24826 19712
rect 25608 19700 25636 19731
rect 26878 19728 26884 19740
rect 26936 19728 26942 19780
rect 27614 19768 27620 19780
rect 27575 19740 27620 19768
rect 27614 19728 27620 19740
rect 27672 19728 27678 19780
rect 28442 19728 28448 19780
rect 28500 19768 28506 19780
rect 30190 19768 30196 19780
rect 28500 19740 30052 19768
rect 30151 19740 30196 19768
rect 28500 19728 28506 19740
rect 27154 19700 27160 19712
rect 25608 19672 27160 19700
rect 27154 19660 27160 19672
rect 27212 19660 27218 19712
rect 28626 19700 28632 19712
rect 28587 19672 28632 19700
rect 28626 19660 28632 19672
rect 28684 19660 28690 19712
rect 30024 19700 30052 19740
rect 30190 19728 30196 19740
rect 30248 19728 30254 19780
rect 30300 19700 30328 19808
rect 33410 19796 33416 19808
rect 33468 19796 33474 19848
rect 33965 19839 34023 19845
rect 33965 19805 33977 19839
rect 34011 19836 34023 19839
rect 43346 19836 43352 19848
rect 34011 19808 43352 19836
rect 34011 19805 34023 19808
rect 33965 19799 34023 19805
rect 43346 19796 43352 19808
rect 43404 19796 43410 19848
rect 30837 19771 30895 19777
rect 30837 19737 30849 19771
rect 30883 19737 30895 19771
rect 30837 19731 30895 19737
rect 32677 19771 32735 19777
rect 32677 19737 32689 19771
rect 32723 19737 32735 19771
rect 33778 19768 33784 19780
rect 33739 19740 33784 19768
rect 32677 19731 32735 19737
rect 30024 19672 30328 19700
rect 30852 19700 30880 19731
rect 31386 19700 31392 19712
rect 30852 19672 31392 19700
rect 31386 19660 31392 19672
rect 31444 19660 31450 19712
rect 32030 19700 32036 19712
rect 31991 19672 32036 19700
rect 32030 19660 32036 19672
rect 32088 19700 32094 19712
rect 32692 19700 32720 19731
rect 33778 19728 33784 19740
rect 33836 19728 33842 19780
rect 34606 19728 34612 19780
rect 34664 19768 34670 19780
rect 35161 19771 35219 19777
rect 35161 19768 35173 19771
rect 34664 19740 35173 19768
rect 34664 19728 34670 19740
rect 35161 19737 35173 19740
rect 35207 19737 35219 19771
rect 35161 19731 35219 19737
rect 35618 19728 35624 19780
rect 35676 19768 35682 19780
rect 35897 19771 35955 19777
rect 35897 19768 35909 19771
rect 35676 19740 35909 19768
rect 35676 19728 35682 19740
rect 35897 19737 35909 19740
rect 35943 19737 35955 19771
rect 35897 19731 35955 19737
rect 32088 19672 32720 19700
rect 32088 19660 32094 19672
rect 1104 19610 44896 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 44896 19610
rect 1104 19536 44896 19558
rect 1946 19456 1952 19508
rect 2004 19496 2010 19508
rect 2041 19499 2099 19505
rect 2041 19496 2053 19499
rect 2004 19468 2053 19496
rect 2004 19456 2010 19468
rect 2041 19465 2053 19468
rect 2087 19465 2099 19499
rect 2498 19496 2504 19508
rect 2459 19468 2504 19496
rect 2041 19459 2099 19465
rect 2498 19456 2504 19468
rect 2556 19456 2562 19508
rect 3973 19499 4031 19505
rect 3973 19465 3985 19499
rect 4019 19496 4031 19499
rect 5626 19496 5632 19508
rect 4019 19468 5632 19496
rect 4019 19465 4031 19468
rect 3973 19459 4031 19465
rect 5626 19456 5632 19468
rect 5684 19456 5690 19508
rect 5810 19496 5816 19508
rect 5771 19468 5816 19496
rect 5810 19456 5816 19468
rect 5868 19456 5874 19508
rect 5920 19468 8708 19496
rect 2314 19388 2320 19440
rect 2372 19428 2378 19440
rect 4700 19431 4758 19437
rect 2372 19400 4476 19428
rect 2372 19388 2378 19400
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19360 1455 19363
rect 1854 19360 1860 19372
rect 1443 19332 1860 19360
rect 1443 19329 1455 19332
rect 1397 19323 1455 19329
rect 1854 19320 1860 19332
rect 1912 19360 1918 19372
rect 2130 19360 2136 19372
rect 1912 19332 2136 19360
rect 1912 19320 1918 19332
rect 2130 19320 2136 19332
rect 2188 19320 2194 19372
rect 2406 19360 2412 19372
rect 2319 19332 2412 19360
rect 2406 19320 2412 19332
rect 2464 19360 2470 19372
rect 3418 19360 3424 19372
rect 2464 19332 3424 19360
rect 2464 19320 2470 19332
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 3694 19360 3700 19372
rect 3651 19332 3700 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 3694 19320 3700 19332
rect 3752 19360 3758 19372
rect 4448 19369 4476 19400
rect 4700 19397 4712 19431
rect 4746 19428 4758 19431
rect 5534 19428 5540 19440
rect 4746 19400 5540 19428
rect 4746 19397 4758 19400
rect 4700 19391 4758 19397
rect 5534 19388 5540 19400
rect 5592 19388 5598 19440
rect 5718 19388 5724 19440
rect 5776 19428 5782 19440
rect 5920 19428 5948 19468
rect 8478 19428 8484 19440
rect 5776 19400 5948 19428
rect 8439 19400 8484 19428
rect 5776 19388 5782 19400
rect 8478 19388 8484 19400
rect 8536 19388 8542 19440
rect 4433 19363 4491 19369
rect 3752 19332 4108 19360
rect 3752 19320 3758 19332
rect 2682 19292 2688 19304
rect 2595 19264 2688 19292
rect 2682 19252 2688 19264
rect 2740 19292 2746 19304
rect 3329 19295 3387 19301
rect 3329 19292 3341 19295
rect 2740 19264 3341 19292
rect 2740 19252 2746 19264
rect 3329 19261 3341 19264
rect 3375 19261 3387 19295
rect 3329 19255 3387 19261
rect 3513 19295 3571 19301
rect 3513 19261 3525 19295
rect 3559 19292 3571 19295
rect 3786 19292 3792 19304
rect 3559 19264 3792 19292
rect 3559 19261 3571 19264
rect 3513 19255 3571 19261
rect 3344 19224 3372 19255
rect 3786 19252 3792 19264
rect 3844 19252 3850 19304
rect 4080 19292 4108 19332
rect 4433 19329 4445 19363
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 4338 19292 4344 19304
rect 4080 19264 4344 19292
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 4154 19224 4160 19236
rect 3344 19196 4160 19224
rect 4154 19184 4160 19196
rect 4212 19184 4218 19236
rect 4246 19184 4252 19236
rect 4304 19184 4310 19236
rect 1581 19159 1639 19165
rect 1581 19125 1593 19159
rect 1627 19156 1639 19159
rect 1946 19156 1952 19168
rect 1627 19128 1952 19156
rect 1627 19125 1639 19128
rect 1581 19119 1639 19125
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 3326 19116 3332 19168
rect 3384 19156 3390 19168
rect 4264 19156 4292 19184
rect 3384 19128 4292 19156
rect 4448 19156 4476 19323
rect 6454 19320 6460 19372
rect 6512 19360 6518 19372
rect 8680 19369 8708 19468
rect 8938 19456 8944 19508
rect 8996 19496 9002 19508
rect 13955 19499 14013 19505
rect 13955 19496 13967 19499
rect 8996 19468 13967 19496
rect 8996 19456 9002 19468
rect 13955 19465 13967 19468
rect 14001 19465 14013 19499
rect 18601 19499 18659 19505
rect 18601 19496 18613 19499
rect 13955 19459 14013 19465
rect 14108 19468 18613 19496
rect 8754 19388 8760 19440
rect 8812 19428 8818 19440
rect 9125 19431 9183 19437
rect 9125 19428 9137 19431
rect 8812 19400 9137 19428
rect 8812 19388 8818 19400
rect 9125 19397 9137 19400
rect 9171 19397 9183 19431
rect 9125 19391 9183 19397
rect 10781 19431 10839 19437
rect 10781 19397 10793 19431
rect 10827 19428 10839 19431
rect 13538 19428 13544 19440
rect 10827 19400 13544 19428
rect 10827 19397 10839 19400
rect 10781 19391 10839 19397
rect 13538 19388 13544 19400
rect 13596 19388 13602 19440
rect 14108 19428 14136 19468
rect 18601 19465 18613 19468
rect 18647 19465 18659 19499
rect 18601 19459 18659 19465
rect 19426 19456 19432 19508
rect 19484 19496 19490 19508
rect 19705 19499 19763 19505
rect 19484 19468 19656 19496
rect 19484 19456 19490 19468
rect 19628 19440 19656 19468
rect 19705 19465 19717 19499
rect 19751 19496 19763 19499
rect 28442 19496 28448 19508
rect 19751 19468 24716 19496
rect 19751 19465 19763 19468
rect 19705 19459 19763 19465
rect 13648 19400 14136 19428
rect 6825 19363 6883 19369
rect 6825 19360 6837 19363
rect 6512 19332 6837 19360
rect 6512 19320 6518 19332
rect 6825 19329 6837 19332
rect 6871 19329 6883 19363
rect 6825 19323 6883 19329
rect 8665 19363 8723 19369
rect 8665 19329 8677 19363
rect 8711 19329 8723 19363
rect 8665 19323 8723 19329
rect 10965 19363 11023 19369
rect 10965 19329 10977 19363
rect 11011 19360 11023 19363
rect 11784 19363 11842 19369
rect 11011 19332 11045 19360
rect 11011 19329 11023 19332
rect 10965 19323 11023 19329
rect 11784 19329 11796 19363
rect 11830 19360 11842 19363
rect 11830 19332 13584 19360
rect 11830 19329 11842 19332
rect 11784 19323 11842 19329
rect 5626 19252 5632 19304
rect 5684 19292 5690 19304
rect 9398 19292 9404 19304
rect 5684 19264 9404 19292
rect 5684 19252 5690 19264
rect 9398 19252 9404 19264
rect 9456 19292 9462 19304
rect 10980 19292 11008 19323
rect 13556 19304 13584 19332
rect 11514 19292 11520 19304
rect 9456 19264 11008 19292
rect 11475 19264 11520 19292
rect 9456 19252 9462 19264
rect 10888 19236 10916 19264
rect 11514 19252 11520 19264
rect 11572 19252 11578 19304
rect 13538 19252 13544 19304
rect 13596 19252 13602 19304
rect 13648 19236 13676 19400
rect 14734 19388 14740 19440
rect 14792 19428 14798 19440
rect 19242 19428 19248 19440
rect 14792 19400 15976 19428
rect 14792 19388 14798 19400
rect 15010 19360 15016 19372
rect 13740 19332 15016 19360
rect 6086 19184 6092 19236
rect 6144 19224 6150 19236
rect 6638 19224 6644 19236
rect 6144 19196 6644 19224
rect 6144 19184 6150 19196
rect 6638 19184 6644 19196
rect 6696 19184 6702 19236
rect 8110 19184 8116 19236
rect 8168 19224 8174 19236
rect 9582 19224 9588 19236
rect 8168 19196 9588 19224
rect 8168 19184 8174 19196
rect 9582 19184 9588 19196
rect 9640 19184 9646 19236
rect 10870 19184 10876 19236
rect 10928 19184 10934 19236
rect 13630 19184 13636 19236
rect 13688 19184 13694 19236
rect 4614 19156 4620 19168
rect 4448 19128 4620 19156
rect 3384 19116 3390 19128
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 5902 19116 5908 19168
rect 5960 19156 5966 19168
rect 9766 19156 9772 19168
rect 5960 19128 9772 19156
rect 5960 19116 5966 19128
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 12897 19159 12955 19165
rect 12897 19125 12909 19159
rect 12943 19156 12955 19159
rect 13262 19156 13268 19168
rect 12943 19128 13268 19156
rect 12943 19125 12955 19128
rect 12897 19119 12955 19125
rect 13262 19116 13268 19128
rect 13320 19116 13326 19168
rect 13538 19116 13544 19168
rect 13596 19156 13602 19168
rect 13740 19156 13768 19332
rect 15010 19320 15016 19332
rect 15068 19320 15074 19372
rect 15194 19360 15200 19372
rect 15155 19332 15200 19360
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 15948 19369 15976 19400
rect 16684 19400 19248 19428
rect 15933 19363 15991 19369
rect 15933 19329 15945 19363
rect 15979 19360 15991 19363
rect 16022 19360 16028 19372
rect 15979 19332 16028 19360
rect 15979 19329 15991 19332
rect 15933 19323 15991 19329
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 16114 19320 16120 19372
rect 16172 19320 16178 19372
rect 16684 19369 16712 19400
rect 19242 19388 19248 19400
rect 19300 19388 19306 19440
rect 19610 19388 19616 19440
rect 19668 19388 19674 19440
rect 19978 19388 19984 19440
rect 20036 19428 20042 19440
rect 20257 19431 20315 19437
rect 20257 19428 20269 19431
rect 20036 19400 20269 19428
rect 20036 19388 20042 19400
rect 20257 19397 20269 19400
rect 20303 19397 20315 19431
rect 20257 19391 20315 19397
rect 20438 19388 20444 19440
rect 20496 19388 20502 19440
rect 21082 19428 21088 19440
rect 21043 19400 21088 19428
rect 21082 19388 21088 19400
rect 21140 19388 21146 19440
rect 21358 19388 21364 19440
rect 21416 19428 21422 19440
rect 23566 19428 23572 19440
rect 21416 19400 23572 19428
rect 21416 19388 21422 19400
rect 23566 19388 23572 19400
rect 23624 19388 23630 19440
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19329 16727 19363
rect 16936 19363 16994 19369
rect 16936 19360 16948 19363
rect 16669 19323 16727 19329
rect 16776 19332 16948 19360
rect 14185 19295 14243 19301
rect 14185 19261 14197 19295
rect 14231 19292 14243 19295
rect 15102 19292 15108 19304
rect 14231 19264 15108 19292
rect 14231 19261 14243 19264
rect 14185 19255 14243 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15286 19252 15292 19304
rect 15344 19292 15350 19304
rect 15473 19295 15531 19301
rect 15473 19292 15485 19295
rect 15344 19264 15485 19292
rect 15344 19252 15350 19264
rect 15473 19261 15485 19264
rect 15519 19261 15531 19295
rect 15473 19255 15531 19261
rect 16132 19233 16160 19320
rect 16482 19252 16488 19304
rect 16540 19292 16546 19304
rect 16776 19292 16804 19332
rect 16936 19329 16948 19332
rect 16982 19360 16994 19363
rect 18322 19360 18328 19372
rect 16982 19332 18328 19360
rect 16982 19329 16994 19332
rect 16936 19323 16994 19329
rect 18322 19320 18328 19332
rect 18380 19320 18386 19372
rect 18506 19360 18512 19372
rect 18432 19332 18512 19360
rect 18432 19292 18460 19332
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 18785 19363 18843 19369
rect 18785 19329 18797 19363
rect 18831 19360 18843 19363
rect 19426 19360 19432 19372
rect 18831 19332 19432 19360
rect 18831 19329 18843 19332
rect 18785 19323 18843 19329
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 19886 19320 19892 19372
rect 19944 19360 19950 19372
rect 20456 19360 20484 19388
rect 19944 19332 20484 19360
rect 22097 19363 22155 19369
rect 19944 19320 19950 19332
rect 22097 19329 22109 19363
rect 22143 19360 22155 19363
rect 22738 19360 22744 19372
rect 22143 19332 22744 19360
rect 22143 19329 22155 19332
rect 22097 19323 22155 19329
rect 22738 19320 22744 19332
rect 22796 19320 22802 19372
rect 23658 19320 23664 19372
rect 23716 19360 23722 19372
rect 24581 19363 24639 19369
rect 24581 19360 24593 19363
rect 23716 19332 24593 19360
rect 23716 19320 23722 19332
rect 24581 19329 24593 19332
rect 24627 19329 24639 19363
rect 24688 19360 24716 19468
rect 25332 19468 28448 19496
rect 25332 19437 25360 19468
rect 28442 19456 28448 19468
rect 28500 19456 28506 19508
rect 28718 19496 28724 19508
rect 28679 19468 28724 19496
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 29454 19496 29460 19508
rect 29415 19468 29460 19496
rect 29454 19456 29460 19468
rect 29512 19456 29518 19508
rect 33134 19496 33140 19508
rect 33095 19468 33140 19496
rect 33134 19456 33140 19468
rect 33192 19456 33198 19508
rect 25317 19431 25375 19437
rect 25317 19397 25329 19431
rect 25363 19397 25375 19431
rect 25317 19391 25375 19397
rect 26053 19431 26111 19437
rect 26053 19397 26065 19431
rect 26099 19428 26111 19431
rect 33318 19428 33324 19440
rect 26099 19400 33324 19428
rect 26099 19397 26111 19400
rect 26053 19391 26111 19397
rect 33318 19388 33324 19400
rect 33376 19388 33382 19440
rect 26694 19360 26700 19372
rect 24688 19332 26700 19360
rect 24581 19323 24639 19329
rect 26694 19320 26700 19332
rect 26752 19320 26758 19372
rect 27338 19320 27344 19372
rect 27396 19360 27402 19372
rect 27433 19363 27491 19369
rect 27433 19360 27445 19363
rect 27396 19332 27445 19360
rect 27396 19320 27402 19332
rect 27433 19329 27445 19332
rect 27479 19329 27491 19363
rect 27433 19323 27491 19329
rect 28169 19363 28227 19369
rect 28169 19329 28181 19363
rect 28215 19360 28227 19363
rect 28813 19363 28871 19369
rect 28813 19360 28825 19363
rect 28215 19332 28825 19360
rect 28215 19329 28227 19332
rect 28169 19323 28227 19329
rect 28813 19329 28825 19332
rect 28859 19360 28871 19363
rect 28902 19360 28908 19372
rect 28859 19332 28908 19360
rect 28859 19329 28871 19332
rect 28813 19323 28871 19329
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 29549 19363 29607 19369
rect 29549 19329 29561 19363
rect 29595 19360 29607 19363
rect 30190 19360 30196 19372
rect 29595 19332 30196 19360
rect 29595 19329 29607 19332
rect 29549 19323 29607 19329
rect 30190 19320 30196 19332
rect 30248 19320 30254 19372
rect 31754 19320 31760 19372
rect 31812 19360 31818 19372
rect 32030 19360 32036 19372
rect 31812 19332 32036 19360
rect 31812 19320 31818 19332
rect 32030 19320 32036 19332
rect 32088 19320 32094 19372
rect 32398 19320 32404 19372
rect 32456 19360 32462 19372
rect 33045 19363 33103 19369
rect 33045 19360 33057 19363
rect 32456 19332 33057 19360
rect 32456 19320 32462 19332
rect 33045 19329 33057 19332
rect 33091 19329 33103 19363
rect 33045 19323 33103 19329
rect 33962 19320 33968 19372
rect 34020 19360 34026 19372
rect 34241 19363 34299 19369
rect 34241 19360 34253 19363
rect 34020 19332 34253 19360
rect 34020 19320 34026 19332
rect 34241 19329 34253 19332
rect 34287 19329 34299 19363
rect 34241 19323 34299 19329
rect 16540 19264 16804 19292
rect 18064 19264 18460 19292
rect 16540 19252 16546 19264
rect 18064 19233 18092 19264
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 19245 19295 19303 19301
rect 19245 19292 19257 19295
rect 19208 19264 19257 19292
rect 19208 19252 19214 19264
rect 19245 19261 19257 19264
rect 19291 19261 19303 19295
rect 19245 19255 19303 19261
rect 19610 19252 19616 19304
rect 19668 19292 19674 19304
rect 19978 19292 19984 19304
rect 19668 19264 19984 19292
rect 19668 19252 19674 19264
rect 19978 19252 19984 19264
rect 20036 19292 20042 19304
rect 20441 19295 20499 19301
rect 20441 19292 20453 19295
rect 20036 19264 20453 19292
rect 20036 19252 20042 19264
rect 20441 19261 20453 19264
rect 20487 19261 20499 19295
rect 21818 19292 21824 19304
rect 21779 19264 21824 19292
rect 20441 19255 20499 19261
rect 21818 19252 21824 19264
rect 21876 19252 21882 19304
rect 23198 19292 23204 19304
rect 23159 19264 23204 19292
rect 23198 19252 23204 19264
rect 23256 19252 23262 19304
rect 25498 19292 25504 19304
rect 25459 19264 25504 19292
rect 25498 19252 25504 19264
rect 25556 19252 25562 19304
rect 26237 19295 26295 19301
rect 26237 19261 26249 19295
rect 26283 19292 26295 19295
rect 34425 19295 34483 19301
rect 26283 19264 31754 19292
rect 26283 19261 26295 19264
rect 26237 19255 26295 19261
rect 16117 19227 16175 19233
rect 16117 19193 16129 19227
rect 16163 19193 16175 19227
rect 16117 19187 16175 19193
rect 18049 19227 18107 19233
rect 18049 19193 18061 19227
rect 18095 19193 18107 19227
rect 18049 19187 18107 19193
rect 18230 19184 18236 19236
rect 18288 19224 18294 19236
rect 18782 19224 18788 19236
rect 18288 19196 18788 19224
rect 18288 19184 18294 19196
rect 18782 19184 18788 19196
rect 18840 19184 18846 19236
rect 19518 19224 19524 19236
rect 19479 19196 19524 19224
rect 19518 19184 19524 19196
rect 19576 19184 19582 19236
rect 19794 19184 19800 19236
rect 19852 19224 19858 19236
rect 20254 19224 20260 19236
rect 19852 19196 20260 19224
rect 19852 19184 19858 19196
rect 20254 19184 20260 19196
rect 20312 19184 20318 19236
rect 23753 19227 23811 19233
rect 23753 19224 23765 19227
rect 20364 19196 23765 19224
rect 13596 19128 13768 19156
rect 13596 19116 13602 19128
rect 18874 19116 18880 19168
rect 18932 19156 18938 19168
rect 19150 19156 19156 19168
rect 18932 19128 19156 19156
rect 18932 19116 18938 19128
rect 19150 19116 19156 19128
rect 19208 19116 19214 19168
rect 19610 19116 19616 19168
rect 19668 19156 19674 19168
rect 20364 19156 20392 19196
rect 23753 19193 23765 19196
rect 23799 19193 23811 19227
rect 27614 19224 27620 19236
rect 27575 19196 27620 19224
rect 23753 19187 23811 19193
rect 27614 19184 27620 19196
rect 27672 19184 27678 19236
rect 31018 19224 31024 19236
rect 27816 19196 31024 19224
rect 19668 19128 20392 19156
rect 19668 19116 19674 19128
rect 20438 19116 20444 19168
rect 20496 19156 20502 19168
rect 20898 19156 20904 19168
rect 20496 19128 20904 19156
rect 20496 19116 20502 19128
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 20993 19159 21051 19165
rect 20993 19125 21005 19159
rect 21039 19156 21051 19159
rect 21358 19156 21364 19168
rect 21039 19128 21364 19156
rect 21039 19125 21051 19128
rect 20993 19119 21051 19125
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 24673 19159 24731 19165
rect 24673 19125 24685 19159
rect 24719 19156 24731 19159
rect 27816 19156 27844 19196
rect 31018 19184 31024 19196
rect 31076 19184 31082 19236
rect 31726 19224 31754 19264
rect 34425 19261 34437 19295
rect 34471 19292 34483 19295
rect 35342 19292 35348 19304
rect 34471 19264 35348 19292
rect 34471 19261 34483 19264
rect 34425 19255 34483 19261
rect 35342 19252 35348 19264
rect 35400 19252 35406 19304
rect 34238 19224 34244 19236
rect 31726 19196 34244 19224
rect 34238 19184 34244 19196
rect 34296 19184 34302 19236
rect 24719 19128 27844 19156
rect 24719 19125 24731 19128
rect 24673 19119 24731 19125
rect 28166 19116 28172 19168
rect 28224 19156 28230 19168
rect 28718 19156 28724 19168
rect 28224 19128 28724 19156
rect 28224 19116 28230 19128
rect 28718 19116 28724 19128
rect 28776 19116 28782 19168
rect 30190 19156 30196 19168
rect 30151 19128 30196 19156
rect 30190 19116 30196 19128
rect 30248 19116 30254 19168
rect 32398 19156 32404 19168
rect 32359 19128 32404 19156
rect 32398 19116 32404 19128
rect 32456 19116 32462 19168
rect 34606 19116 34612 19168
rect 34664 19156 34670 19168
rect 34885 19159 34943 19165
rect 34885 19156 34897 19159
rect 34664 19128 34897 19156
rect 34664 19116 34670 19128
rect 34885 19125 34897 19128
rect 34931 19125 34943 19159
rect 35618 19156 35624 19168
rect 35579 19128 35624 19156
rect 34885 19119 34943 19125
rect 35618 19116 35624 19128
rect 35676 19116 35682 19168
rect 1104 19066 44896 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 44896 19066
rect 1104 18992 44896 19014
rect 2038 18952 2044 18964
rect 1999 18924 2044 18952
rect 2038 18912 2044 18924
rect 2096 18912 2102 18964
rect 3142 18912 3148 18964
rect 3200 18952 3206 18964
rect 3237 18955 3295 18961
rect 3237 18952 3249 18955
rect 3200 18924 3249 18952
rect 3200 18912 3206 18924
rect 3237 18921 3249 18924
rect 3283 18921 3295 18955
rect 3237 18915 3295 18921
rect 4706 18912 4712 18964
rect 4764 18952 4770 18964
rect 4764 18924 6592 18952
rect 4764 18912 4770 18924
rect 3694 18844 3700 18896
rect 3752 18884 3758 18896
rect 5902 18884 5908 18896
rect 3752 18856 5908 18884
rect 3752 18844 3758 18856
rect 5902 18844 5908 18856
rect 5960 18844 5966 18896
rect 1026 18776 1032 18828
rect 1084 18816 1090 18828
rect 1857 18819 1915 18825
rect 1857 18816 1869 18819
rect 1084 18788 1869 18816
rect 1084 18776 1090 18788
rect 1857 18785 1869 18788
rect 1903 18785 1915 18819
rect 2682 18816 2688 18828
rect 2643 18788 2688 18816
rect 1857 18779 1915 18785
rect 2682 18776 2688 18788
rect 2740 18776 2746 18828
rect 2777 18819 2835 18825
rect 2777 18785 2789 18819
rect 2823 18816 2835 18819
rect 5626 18816 5632 18828
rect 2823 18788 5632 18816
rect 2823 18785 2835 18788
rect 2777 18779 2835 18785
rect 5626 18776 5632 18788
rect 5684 18776 5690 18828
rect 6564 18825 6592 18924
rect 9582 18912 9588 18964
rect 9640 18952 9646 18964
rect 13722 18952 13728 18964
rect 9640 18924 13728 18952
rect 9640 18912 9646 18924
rect 13722 18912 13728 18924
rect 13780 18912 13786 18964
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 16390 18952 16396 18964
rect 14148 18924 16396 18952
rect 14148 18912 14154 18924
rect 16390 18912 16396 18924
rect 16448 18912 16454 18964
rect 17972 18924 20116 18952
rect 9674 18884 9680 18896
rect 7024 18856 9680 18884
rect 6089 18819 6147 18825
rect 6089 18785 6101 18819
rect 6135 18785 6147 18819
rect 6089 18779 6147 18785
rect 6549 18819 6607 18825
rect 6549 18785 6561 18819
rect 6595 18785 6607 18819
rect 6549 18779 6607 18785
rect 1118 18708 1124 18760
rect 1176 18748 1182 18760
rect 1765 18751 1823 18757
rect 1765 18748 1777 18751
rect 1176 18720 1777 18748
rect 1176 18708 1182 18720
rect 1765 18717 1777 18720
rect 1811 18717 1823 18751
rect 2038 18748 2044 18760
rect 1999 18720 2044 18748
rect 1765 18711 1823 18717
rect 2038 18708 2044 18720
rect 2096 18708 2102 18760
rect 2869 18751 2927 18757
rect 2869 18717 2881 18751
rect 2915 18748 2927 18751
rect 3234 18748 3240 18760
rect 2915 18720 3240 18748
rect 2915 18717 2927 18720
rect 2869 18711 2927 18717
rect 3234 18708 3240 18720
rect 3292 18708 3298 18760
rect 4249 18751 4307 18757
rect 4249 18717 4261 18751
rect 4295 18748 4307 18751
rect 4522 18748 4528 18760
rect 4295 18720 4528 18748
rect 4295 18717 4307 18720
rect 4249 18711 4307 18717
rect 4522 18708 4528 18720
rect 4580 18708 4586 18760
rect 6104 18748 6132 18779
rect 7024 18748 7052 18856
rect 9674 18844 9680 18856
rect 9732 18844 9738 18896
rect 10428 18856 11376 18884
rect 8202 18816 8208 18828
rect 8163 18788 8208 18816
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 9030 18776 9036 18828
rect 9088 18816 9094 18828
rect 10428 18816 10456 18856
rect 10594 18816 10600 18828
rect 9088 18788 10456 18816
rect 10555 18788 10600 18816
rect 9088 18776 9094 18788
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 6104 18720 7052 18748
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 11241 18751 11299 18757
rect 11241 18717 11253 18751
rect 11287 18717 11299 18751
rect 11348 18748 11376 18856
rect 13538 18844 13544 18896
rect 13596 18884 13602 18896
rect 17034 18884 17040 18896
rect 13596 18856 16160 18884
rect 13596 18844 13602 18856
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11701 18819 11759 18825
rect 11701 18816 11713 18819
rect 11572 18788 11713 18816
rect 11572 18776 11578 18788
rect 11701 18785 11713 18788
rect 11747 18785 11759 18819
rect 11701 18779 11759 18785
rect 14093 18819 14151 18825
rect 14093 18785 14105 18819
rect 14139 18816 14151 18819
rect 14274 18816 14280 18828
rect 14139 18788 14280 18816
rect 14139 18785 14151 18788
rect 14093 18779 14151 18785
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 15930 18816 15936 18828
rect 15891 18788 15936 18816
rect 15930 18776 15936 18788
rect 15988 18776 15994 18828
rect 14366 18748 14372 18760
rect 11348 18720 14228 18748
rect 14327 18720 14372 18748
rect 11241 18711 11299 18717
rect 4706 18640 4712 18692
rect 4764 18680 4770 18692
rect 5905 18683 5963 18689
rect 5905 18680 5917 18683
rect 4764 18652 5917 18680
rect 4764 18640 4770 18652
rect 5905 18649 5917 18652
rect 5951 18649 5963 18683
rect 5905 18643 5963 18649
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18612 1639 18615
rect 2682 18612 2688 18624
rect 1627 18584 2688 18612
rect 1627 18581 1639 18584
rect 1581 18575 1639 18581
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 3786 18572 3792 18624
rect 3844 18612 3850 18624
rect 8404 18612 8432 18711
rect 10410 18640 10416 18692
rect 10468 18680 10474 18692
rect 10870 18680 10876 18692
rect 10468 18652 10876 18680
rect 10468 18640 10474 18652
rect 10870 18640 10876 18652
rect 10928 18640 10934 18692
rect 11054 18680 11060 18692
rect 11015 18652 11060 18680
rect 11054 18640 11060 18652
rect 11112 18640 11118 18692
rect 3844 18584 8432 18612
rect 3844 18572 3850 18584
rect 9490 18572 9496 18624
rect 9548 18612 9554 18624
rect 10502 18612 10508 18624
rect 9548 18584 10508 18612
rect 9548 18572 9554 18584
rect 10502 18572 10508 18584
rect 10560 18612 10566 18624
rect 11256 18612 11284 18711
rect 11968 18683 12026 18689
rect 11968 18649 11980 18683
rect 12014 18680 12026 18683
rect 13538 18680 13544 18692
rect 12014 18652 13544 18680
rect 12014 18649 12026 18652
rect 11968 18643 12026 18649
rect 13538 18640 13544 18652
rect 13596 18640 13602 18692
rect 14200 18680 14228 18720
rect 14366 18708 14372 18720
rect 14424 18708 14430 18760
rect 16132 18748 16160 18856
rect 16224 18856 17040 18884
rect 16224 18825 16252 18856
rect 17034 18844 17040 18856
rect 17092 18844 17098 18896
rect 16209 18819 16267 18825
rect 16209 18785 16221 18819
rect 16255 18785 16267 18819
rect 16209 18779 16267 18785
rect 16853 18819 16911 18825
rect 16853 18785 16865 18819
rect 16899 18816 16911 18819
rect 17862 18816 17868 18828
rect 16899 18788 17868 18816
rect 16899 18785 16911 18788
rect 16853 18779 16911 18785
rect 17862 18776 17868 18788
rect 17920 18776 17926 18828
rect 16132 18720 17448 18748
rect 17126 18680 17132 18692
rect 14200 18652 17132 18680
rect 10560 18584 11284 18612
rect 10560 18572 10566 18584
rect 12710 18572 12716 18624
rect 12768 18612 12774 18624
rect 13081 18615 13139 18621
rect 13081 18612 13093 18615
rect 12768 18584 13093 18612
rect 12768 18572 12774 18584
rect 13081 18581 13093 18584
rect 13127 18581 13139 18615
rect 13081 18575 13139 18581
rect 13170 18572 13176 18624
rect 13228 18612 13234 18624
rect 14734 18612 14740 18624
rect 13228 18584 14740 18612
rect 13228 18572 13234 18584
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 17052 18621 17080 18652
rect 17126 18640 17132 18652
rect 17184 18640 17190 18692
rect 17420 18680 17448 18720
rect 17494 18708 17500 18760
rect 17552 18748 17558 18760
rect 17678 18748 17684 18760
rect 17552 18720 17684 18748
rect 17552 18708 17558 18720
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 17972 18748 18000 18924
rect 20088 18896 20116 18924
rect 20254 18912 20260 18964
rect 20312 18952 20318 18964
rect 21542 18952 21548 18964
rect 20312 18924 20576 18952
rect 21503 18924 21548 18952
rect 20312 18912 20318 18924
rect 18138 18884 18144 18896
rect 18099 18856 18144 18884
rect 18138 18844 18144 18856
rect 18196 18844 18202 18896
rect 19518 18884 19524 18896
rect 18248 18856 19524 18884
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18248 18816 18276 18856
rect 19518 18844 19524 18856
rect 19576 18844 19582 18896
rect 19613 18887 19671 18893
rect 19613 18853 19625 18887
rect 19659 18884 19671 18887
rect 19794 18884 19800 18896
rect 19659 18856 19800 18884
rect 19659 18853 19671 18856
rect 19613 18847 19671 18853
rect 19794 18844 19800 18856
rect 19852 18844 19858 18896
rect 20070 18844 20076 18896
rect 20128 18844 20134 18896
rect 20346 18844 20352 18896
rect 20404 18884 20410 18896
rect 20441 18887 20499 18893
rect 20441 18884 20453 18887
rect 20404 18856 20453 18884
rect 20404 18844 20410 18856
rect 20441 18853 20453 18856
rect 20487 18853 20499 18887
rect 20548 18884 20576 18924
rect 21542 18912 21548 18924
rect 21600 18912 21606 18964
rect 22189 18955 22247 18961
rect 22189 18921 22201 18955
rect 22235 18952 22247 18955
rect 22554 18952 22560 18964
rect 22235 18924 22560 18952
rect 22235 18921 22247 18924
rect 22189 18915 22247 18921
rect 22554 18912 22560 18924
rect 22612 18912 22618 18964
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 24302 18952 24308 18964
rect 23532 18924 24308 18952
rect 23532 18912 23538 18924
rect 24302 18912 24308 18924
rect 24360 18952 24366 18964
rect 24397 18955 24455 18961
rect 24397 18952 24409 18955
rect 24360 18924 24409 18952
rect 24360 18912 24366 18924
rect 24397 18921 24409 18924
rect 24443 18921 24455 18955
rect 24946 18952 24952 18964
rect 24907 18924 24952 18952
rect 24397 18915 24455 18921
rect 24946 18912 24952 18924
rect 25004 18912 25010 18964
rect 27246 18952 27252 18964
rect 27207 18924 27252 18952
rect 27246 18912 27252 18924
rect 27304 18912 27310 18964
rect 27614 18912 27620 18964
rect 27672 18952 27678 18964
rect 36262 18952 36268 18964
rect 27672 18924 36268 18952
rect 27672 18912 27678 18924
rect 36262 18912 36268 18924
rect 36320 18912 36326 18964
rect 21450 18884 21456 18896
rect 20548 18856 21456 18884
rect 20441 18847 20499 18853
rect 21450 18844 21456 18856
rect 21508 18844 21514 18896
rect 30098 18844 30104 18896
rect 30156 18884 30162 18896
rect 35618 18884 35624 18896
rect 30156 18856 35624 18884
rect 30156 18844 30162 18856
rect 35618 18844 35624 18856
rect 35676 18844 35682 18896
rect 19705 18819 19763 18825
rect 18104 18788 18276 18816
rect 19306 18788 19656 18816
rect 18104 18776 18110 18788
rect 19306 18748 19334 18788
rect 19628 18760 19656 18788
rect 19705 18785 19717 18819
rect 19751 18785 19763 18819
rect 30558 18816 30564 18828
rect 19705 18779 19763 18785
rect 20180 18788 30564 18816
rect 17797 18720 18000 18748
rect 18708 18720 19334 18748
rect 17797 18680 17825 18720
rect 17420 18652 17825 18680
rect 17865 18683 17923 18689
rect 17865 18649 17877 18683
rect 17911 18680 17923 18683
rect 18046 18680 18052 18692
rect 17911 18652 18052 18680
rect 17911 18649 17923 18652
rect 17865 18643 17923 18649
rect 18046 18640 18052 18652
rect 18104 18640 18110 18692
rect 18708 18680 18736 18720
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 19720 18748 19748 18779
rect 19720 18744 20024 18748
rect 20180 18744 20208 18788
rect 30558 18776 30564 18788
rect 30616 18776 30622 18828
rect 19720 18720 20208 18744
rect 19996 18716 20208 18720
rect 20257 18751 20315 18757
rect 20257 18717 20269 18751
rect 20303 18748 20315 18751
rect 20438 18748 20444 18760
rect 20303 18720 20444 18748
rect 20303 18717 20315 18720
rect 20257 18711 20315 18717
rect 20438 18708 20444 18720
rect 20496 18708 20502 18760
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 20864 18720 21097 18748
rect 20864 18708 20870 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 21542 18708 21548 18760
rect 21600 18748 21606 18760
rect 21729 18751 21787 18757
rect 21729 18748 21741 18751
rect 21600 18720 21741 18748
rect 21600 18708 21606 18720
rect 21729 18717 21741 18720
rect 21775 18717 21787 18751
rect 22370 18748 22376 18760
rect 22331 18720 22376 18748
rect 21729 18711 21787 18717
rect 22370 18708 22376 18720
rect 22428 18708 22434 18760
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 22796 18720 23029 18748
rect 22796 18708 22802 18720
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 24762 18708 24768 18760
rect 24820 18748 24826 18760
rect 30742 18748 30748 18760
rect 24820 18720 30748 18748
rect 24820 18708 24826 18720
rect 30742 18708 30748 18720
rect 30800 18708 30806 18760
rect 18156 18652 18736 18680
rect 16945 18615 17003 18621
rect 16945 18612 16957 18615
rect 16724 18584 16957 18612
rect 16724 18572 16730 18584
rect 16945 18581 16957 18584
rect 16991 18581 17003 18615
rect 16945 18575 17003 18581
rect 17037 18615 17095 18621
rect 17037 18581 17049 18615
rect 17083 18581 17095 18615
rect 17037 18575 17095 18581
rect 17405 18615 17463 18621
rect 17405 18581 17417 18615
rect 17451 18612 17463 18615
rect 18156 18612 18184 18652
rect 18782 18640 18788 18692
rect 18840 18680 18846 18692
rect 19245 18683 19303 18689
rect 19245 18680 19257 18683
rect 18840 18652 19257 18680
rect 18840 18640 18846 18652
rect 19245 18649 19257 18652
rect 19291 18649 19303 18683
rect 19245 18643 19303 18649
rect 19794 18640 19800 18692
rect 19852 18680 19858 18692
rect 21634 18680 21640 18692
rect 19852 18652 21640 18680
rect 19852 18640 19858 18652
rect 21634 18640 21640 18652
rect 21692 18640 21698 18692
rect 22646 18640 22652 18692
rect 22704 18680 22710 18692
rect 24780 18680 24808 18708
rect 22704 18652 24808 18680
rect 25593 18683 25651 18689
rect 22704 18640 22710 18652
rect 25593 18649 25605 18683
rect 25639 18680 25651 18683
rect 26970 18680 26976 18692
rect 25639 18652 26976 18680
rect 25639 18649 25651 18652
rect 25593 18643 25651 18649
rect 26970 18640 26976 18652
rect 27028 18640 27034 18692
rect 27157 18683 27215 18689
rect 27157 18649 27169 18683
rect 27203 18649 27215 18683
rect 27157 18643 27215 18649
rect 18322 18612 18328 18624
rect 17451 18584 18184 18612
rect 18283 18584 18328 18612
rect 17451 18581 17463 18584
rect 17405 18575 17463 18581
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 18506 18572 18512 18624
rect 18564 18612 18570 18624
rect 20901 18615 20959 18621
rect 20901 18612 20913 18615
rect 18564 18584 20913 18612
rect 18564 18572 18570 18584
rect 20901 18581 20913 18584
rect 20947 18581 20959 18615
rect 20901 18575 20959 18581
rect 20990 18572 20996 18624
rect 21048 18612 21054 18624
rect 22833 18615 22891 18621
rect 22833 18612 22845 18615
rect 21048 18584 22845 18612
rect 21048 18572 21054 18584
rect 22833 18581 22845 18584
rect 22879 18581 22891 18615
rect 22833 18575 22891 18581
rect 23569 18615 23627 18621
rect 23569 18581 23581 18615
rect 23615 18612 23627 18615
rect 24486 18612 24492 18624
rect 23615 18584 24492 18612
rect 23615 18581 23627 18584
rect 23569 18575 23627 18581
rect 24486 18572 24492 18584
rect 24544 18572 24550 18624
rect 26602 18612 26608 18624
rect 26563 18584 26608 18612
rect 26602 18572 26608 18584
rect 26660 18612 26666 18624
rect 27172 18612 27200 18643
rect 30190 18640 30196 18692
rect 30248 18680 30254 18692
rect 43990 18680 43996 18692
rect 30248 18652 43996 18680
rect 30248 18640 30254 18652
rect 43990 18640 43996 18652
rect 44048 18640 44054 18692
rect 33962 18612 33968 18624
rect 26660 18584 27200 18612
rect 33923 18584 33968 18612
rect 26660 18572 26666 18584
rect 33962 18572 33968 18584
rect 34020 18572 34026 18624
rect 1104 18522 44896 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 44896 18522
rect 1104 18448 44896 18470
rect 2317 18411 2375 18417
rect 2317 18377 2329 18411
rect 2363 18408 2375 18411
rect 4154 18408 4160 18420
rect 2363 18380 4160 18408
rect 2363 18377 2375 18380
rect 2317 18371 2375 18377
rect 4154 18368 4160 18380
rect 4212 18368 4218 18420
rect 9122 18408 9128 18420
rect 4264 18380 9128 18408
rect 4264 18340 4292 18380
rect 9122 18368 9128 18380
rect 9180 18368 9186 18420
rect 9214 18368 9220 18420
rect 9272 18408 9278 18420
rect 11974 18408 11980 18420
rect 9272 18380 11980 18408
rect 9272 18368 9278 18380
rect 11974 18368 11980 18380
rect 12032 18368 12038 18420
rect 14366 18408 14372 18420
rect 12406 18380 14372 18408
rect 3712 18312 4292 18340
rect 4700 18343 4758 18349
rect 3712 18281 3740 18312
rect 4700 18309 4712 18343
rect 4746 18340 4758 18343
rect 4982 18340 4988 18352
rect 4746 18312 4988 18340
rect 4746 18309 4758 18312
rect 4700 18303 4758 18309
rect 4982 18300 4988 18312
rect 5040 18300 5046 18352
rect 5442 18300 5448 18352
rect 5500 18340 5506 18352
rect 7834 18340 7840 18352
rect 5500 18312 7840 18340
rect 5500 18300 5506 18312
rect 7834 18300 7840 18312
rect 7892 18300 7898 18352
rect 8297 18343 8355 18349
rect 8297 18309 8309 18343
rect 8343 18340 8355 18343
rect 12406 18340 12434 18380
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 16022 18408 16028 18420
rect 15983 18380 16028 18408
rect 16022 18368 16028 18380
rect 16080 18368 16086 18420
rect 16669 18411 16727 18417
rect 16669 18377 16681 18411
rect 16715 18408 16727 18411
rect 17310 18408 17316 18420
rect 16715 18380 17316 18408
rect 16715 18377 16727 18380
rect 16669 18371 16727 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 18230 18368 18236 18420
rect 18288 18408 18294 18420
rect 18288 18380 18333 18408
rect 18288 18368 18294 18380
rect 18874 18368 18880 18420
rect 18932 18408 18938 18420
rect 20806 18408 20812 18420
rect 18932 18380 20812 18408
rect 18932 18368 18938 18380
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 21358 18408 21364 18420
rect 20916 18380 21364 18408
rect 20916 18340 20944 18380
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 21450 18368 21456 18420
rect 21508 18408 21514 18420
rect 22373 18411 22431 18417
rect 22373 18408 22385 18411
rect 21508 18380 22385 18408
rect 21508 18368 21514 18380
rect 22373 18377 22385 18380
rect 22419 18377 22431 18411
rect 22922 18408 22928 18420
rect 22883 18380 22928 18408
rect 22373 18371 22431 18377
rect 8343 18312 12434 18340
rect 14108 18312 20944 18340
rect 21177 18343 21235 18349
rect 8343 18309 8355 18312
rect 8297 18303 8355 18309
rect 14108 18284 14136 18312
rect 21177 18309 21189 18343
rect 21223 18340 21235 18343
rect 21726 18340 21732 18352
rect 21223 18312 21732 18340
rect 21223 18309 21235 18312
rect 21177 18303 21235 18309
rect 21726 18300 21732 18312
rect 21784 18300 21790 18352
rect 22278 18340 22284 18352
rect 22239 18312 22284 18340
rect 22278 18300 22284 18312
rect 22336 18300 22342 18352
rect 22388 18340 22416 18371
rect 22922 18368 22928 18380
rect 22980 18368 22986 18420
rect 23566 18408 23572 18420
rect 23527 18380 23572 18408
rect 23566 18368 23572 18380
rect 23624 18368 23630 18420
rect 24762 18408 24768 18420
rect 24723 18380 24768 18408
rect 24762 18368 24768 18380
rect 24820 18368 24826 18420
rect 24946 18368 24952 18420
rect 25004 18408 25010 18420
rect 25777 18411 25835 18417
rect 25777 18408 25789 18411
rect 25004 18380 25789 18408
rect 25004 18368 25010 18380
rect 25777 18377 25789 18380
rect 25823 18377 25835 18411
rect 25777 18371 25835 18377
rect 27430 18368 27436 18420
rect 27488 18408 27494 18420
rect 28074 18408 28080 18420
rect 27488 18380 28080 18408
rect 27488 18368 27494 18380
rect 28074 18368 28080 18380
rect 28132 18368 28138 18420
rect 29270 18408 29276 18420
rect 29231 18380 29276 18408
rect 29270 18368 29276 18380
rect 29328 18368 29334 18420
rect 28353 18343 28411 18349
rect 22388 18312 28304 18340
rect 3697 18275 3755 18281
rect 3697 18241 3709 18275
rect 3743 18241 3755 18275
rect 3970 18272 3976 18284
rect 3931 18244 3976 18272
rect 3697 18235 3755 18241
rect 3970 18232 3976 18244
rect 4028 18232 4034 18284
rect 4430 18272 4436 18284
rect 4391 18244 4436 18272
rect 4430 18232 4436 18244
rect 4488 18232 4494 18284
rect 5626 18232 5632 18284
rect 5684 18272 5690 18284
rect 6270 18272 6276 18284
rect 5684 18244 6276 18272
rect 5684 18232 5690 18244
rect 6270 18232 6276 18244
rect 6328 18272 6334 18284
rect 6328 18244 7052 18272
rect 6328 18232 6334 18244
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18173 2191 18207
rect 2133 18167 2191 18173
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18204 2283 18207
rect 6914 18204 6920 18216
rect 2271 18176 4476 18204
rect 6875 18176 6920 18204
rect 2271 18173 2283 18176
rect 2225 18167 2283 18173
rect 2148 18136 2176 18167
rect 2866 18136 2872 18148
rect 2148 18108 2872 18136
rect 2866 18096 2872 18108
rect 2924 18096 2930 18148
rect 1489 18071 1547 18077
rect 1489 18037 1501 18071
rect 1535 18068 1547 18071
rect 2590 18068 2596 18080
rect 1535 18040 2596 18068
rect 1535 18037 1547 18040
rect 1489 18031 1547 18037
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 2685 18071 2743 18077
rect 2685 18037 2697 18071
rect 2731 18068 2743 18071
rect 3326 18068 3332 18080
rect 2731 18040 3332 18068
rect 2731 18037 2743 18040
rect 2685 18031 2743 18037
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 4448 18068 4476 18176
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 7024 18204 7052 18244
rect 11330 18232 11336 18284
rect 11388 18272 11394 18284
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 11388 18244 11529 18272
rect 11388 18232 11394 18244
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 14090 18272 14096 18284
rect 14003 18244 14096 18272
rect 11517 18235 11575 18241
rect 14090 18232 14096 18244
rect 14148 18232 14154 18284
rect 14360 18275 14418 18281
rect 14360 18241 14372 18275
rect 14406 18272 14418 18275
rect 16482 18272 16488 18284
rect 14406 18244 16488 18272
rect 14406 18241 14418 18244
rect 14360 18235 14418 18241
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 16666 18232 16672 18284
rect 16724 18272 16730 18284
rect 17037 18275 17095 18281
rect 17037 18272 17049 18275
rect 16724 18244 17049 18272
rect 16724 18232 16730 18244
rect 17037 18241 17049 18244
rect 17083 18241 17095 18275
rect 17037 18235 17095 18241
rect 17126 18232 17132 18284
rect 17184 18272 17190 18284
rect 17402 18272 17408 18284
rect 17184 18244 17408 18272
rect 17184 18232 17190 18244
rect 17402 18232 17408 18244
rect 17460 18232 17466 18284
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 17512 18244 18337 18272
rect 8481 18207 8539 18213
rect 8481 18204 8493 18207
rect 7024 18176 8493 18204
rect 8481 18173 8493 18176
rect 8527 18173 8539 18207
rect 9030 18204 9036 18216
rect 8991 18176 9036 18204
rect 8481 18167 8539 18173
rect 9030 18164 9036 18176
rect 9088 18164 9094 18216
rect 10597 18207 10655 18213
rect 10597 18173 10609 18207
rect 10643 18173 10655 18207
rect 10597 18167 10655 18173
rect 10781 18207 10839 18213
rect 10781 18173 10793 18207
rect 10827 18204 10839 18207
rect 11701 18207 11759 18213
rect 10827 18176 11376 18204
rect 11701 18188 11713 18207
rect 10827 18173 10839 18176
rect 10781 18167 10839 18173
rect 5813 18139 5871 18145
rect 5813 18105 5825 18139
rect 5859 18136 5871 18139
rect 5859 18108 6592 18136
rect 5859 18105 5871 18108
rect 5813 18099 5871 18105
rect 6362 18068 6368 18080
rect 4448 18040 6368 18068
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 6564 18068 6592 18108
rect 8846 18068 8852 18080
rect 6564 18040 8852 18068
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 10612 18068 10640 18167
rect 11348 18148 11376 18176
rect 11624 18173 11713 18188
rect 11747 18173 11759 18207
rect 11624 18167 11759 18173
rect 11624 18160 11744 18167
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 12492 18176 12537 18204
rect 12492 18164 12498 18176
rect 15286 18164 15292 18216
rect 15344 18204 15350 18216
rect 16850 18204 16856 18216
rect 15344 18176 16856 18204
rect 15344 18164 15350 18176
rect 16850 18164 16856 18176
rect 16908 18164 16914 18216
rect 17218 18204 17224 18216
rect 17179 18176 17224 18204
rect 17218 18164 17224 18176
rect 17276 18164 17282 18216
rect 17310 18164 17316 18216
rect 17368 18204 17374 18216
rect 17512 18204 17540 18244
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 18325 18235 18383 18241
rect 18782 18232 18788 18284
rect 18840 18272 18846 18284
rect 19981 18275 20039 18281
rect 19981 18272 19993 18275
rect 18840 18244 19993 18272
rect 18840 18232 18846 18244
rect 19981 18241 19993 18244
rect 20027 18241 20039 18275
rect 20901 18275 20959 18281
rect 20901 18272 20913 18275
rect 19981 18235 20039 18241
rect 20088 18244 20913 18272
rect 17368 18176 17540 18204
rect 17368 18164 17374 18176
rect 17862 18164 17868 18216
rect 17920 18204 17926 18216
rect 18417 18207 18475 18213
rect 18417 18204 18429 18207
rect 17920 18176 18429 18204
rect 17920 18164 17926 18176
rect 18417 18173 18429 18176
rect 18463 18204 18475 18207
rect 19518 18204 19524 18216
rect 18463 18176 19334 18204
rect 19479 18176 19524 18204
rect 18463 18173 18475 18176
rect 18417 18167 18475 18173
rect 11146 18136 11152 18148
rect 10980 18108 11152 18136
rect 10980 18068 11008 18108
rect 11146 18096 11152 18108
rect 11204 18096 11210 18148
rect 11330 18096 11336 18148
rect 11388 18096 11394 18148
rect 11422 18096 11428 18148
rect 11480 18136 11486 18148
rect 11624 18136 11652 18160
rect 11480 18108 11652 18136
rect 11480 18096 11486 18108
rect 12158 18096 12164 18148
rect 12216 18136 12222 18148
rect 12986 18136 12992 18148
rect 12216 18108 12992 18136
rect 12216 18096 12222 18108
rect 12986 18096 12992 18108
rect 13044 18096 13050 18148
rect 18506 18136 18512 18148
rect 15396 18108 18512 18136
rect 10612 18040 11008 18068
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 15396 18068 15424 18108
rect 18506 18096 18512 18108
rect 18564 18096 18570 18148
rect 19150 18136 19156 18148
rect 19111 18108 19156 18136
rect 19150 18096 19156 18108
rect 19208 18096 19214 18148
rect 19306 18136 19334 18176
rect 19518 18164 19524 18176
rect 19576 18164 19582 18216
rect 19702 18164 19708 18216
rect 19760 18204 19766 18216
rect 20088 18204 20116 18244
rect 20901 18241 20913 18244
rect 20947 18241 20959 18275
rect 20901 18235 20959 18241
rect 20438 18204 20444 18216
rect 19760 18176 20116 18204
rect 20399 18176 20444 18204
rect 19760 18164 19766 18176
rect 20438 18164 20444 18176
rect 20496 18164 20502 18216
rect 20916 18204 20944 18235
rect 20990 18232 20996 18284
rect 21048 18272 21054 18284
rect 21048 18244 21093 18272
rect 21048 18232 21054 18244
rect 23014 18232 23020 18284
rect 23072 18272 23078 18284
rect 23109 18275 23167 18281
rect 23109 18272 23121 18275
rect 23072 18244 23121 18272
rect 23072 18232 23078 18244
rect 23109 18241 23121 18244
rect 23155 18241 23167 18275
rect 23109 18235 23167 18241
rect 24026 18232 24032 18284
rect 24084 18272 24090 18284
rect 24213 18275 24271 18281
rect 24213 18272 24225 18275
rect 24084 18244 24225 18272
rect 24084 18232 24090 18244
rect 24213 18241 24225 18244
rect 24259 18272 24271 18275
rect 24762 18272 24768 18284
rect 24259 18244 24768 18272
rect 24259 18241 24271 18244
rect 24213 18235 24271 18241
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 25314 18272 25320 18284
rect 25227 18244 25320 18272
rect 25314 18232 25320 18244
rect 25372 18272 25378 18284
rect 27246 18272 27252 18284
rect 25372 18244 27252 18272
rect 25372 18232 25378 18244
rect 27246 18232 27252 18244
rect 27304 18232 27310 18284
rect 27617 18275 27675 18281
rect 27617 18241 27629 18275
rect 27663 18272 27675 18275
rect 28166 18272 28172 18284
rect 27663 18244 28172 18272
rect 27663 18241 27675 18244
rect 27617 18235 27675 18241
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 21358 18204 21364 18216
rect 20916 18176 21364 18204
rect 21358 18164 21364 18176
rect 21416 18164 21422 18216
rect 23290 18164 23296 18216
rect 23348 18204 23354 18216
rect 26326 18204 26332 18216
rect 23348 18176 26332 18204
rect 23348 18164 23354 18176
rect 26326 18164 26332 18176
rect 26384 18164 26390 18216
rect 28276 18204 28304 18312
rect 28353 18309 28365 18343
rect 28399 18340 28411 18343
rect 28994 18340 29000 18352
rect 28399 18312 29000 18340
rect 28399 18309 28411 18312
rect 28353 18303 28411 18309
rect 28994 18300 29000 18312
rect 29052 18300 29058 18352
rect 29181 18343 29239 18349
rect 29181 18309 29193 18343
rect 29227 18309 29239 18343
rect 29181 18303 29239 18309
rect 30193 18343 30251 18349
rect 30193 18309 30205 18343
rect 30239 18340 30251 18343
rect 30282 18340 30288 18352
rect 30239 18312 30288 18340
rect 30239 18309 30251 18312
rect 30193 18303 30251 18309
rect 29196 18216 29224 18303
rect 30282 18300 30288 18312
rect 30340 18300 30346 18352
rect 29914 18232 29920 18284
rect 29972 18272 29978 18284
rect 30009 18275 30067 18281
rect 30009 18272 30021 18275
rect 29972 18244 30021 18272
rect 29972 18232 29978 18244
rect 30009 18241 30021 18244
rect 30055 18241 30067 18275
rect 30009 18235 30067 18241
rect 28350 18204 28356 18216
rect 28276 18176 28356 18204
rect 28350 18164 28356 18176
rect 28408 18164 28414 18216
rect 29178 18164 29184 18216
rect 29236 18164 29242 18216
rect 19978 18136 19984 18148
rect 19306 18108 19984 18136
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 20349 18139 20407 18145
rect 20349 18105 20361 18139
rect 20395 18136 20407 18139
rect 20530 18136 20536 18148
rect 20395 18108 20536 18136
rect 20395 18105 20407 18108
rect 20349 18099 20407 18105
rect 20530 18096 20536 18108
rect 20588 18096 20594 18148
rect 20640 18108 22040 18136
rect 11112 18040 15424 18068
rect 15473 18071 15531 18077
rect 11112 18028 11118 18040
rect 15473 18037 15485 18071
rect 15519 18068 15531 18071
rect 16482 18068 16488 18080
rect 15519 18040 16488 18068
rect 15519 18037 15531 18040
rect 15473 18031 15531 18037
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 16942 18028 16948 18080
rect 17000 18068 17006 18080
rect 17865 18071 17923 18077
rect 17865 18068 17877 18071
rect 17000 18040 17877 18068
rect 17000 18028 17006 18040
rect 17865 18037 17877 18040
rect 17911 18037 17923 18071
rect 17865 18031 17923 18037
rect 18138 18028 18144 18080
rect 18196 18068 18202 18080
rect 19061 18071 19119 18077
rect 19061 18068 19073 18071
rect 18196 18040 19073 18068
rect 18196 18028 18202 18040
rect 19061 18037 19073 18040
rect 19107 18037 19119 18071
rect 19061 18031 19119 18037
rect 19518 18028 19524 18080
rect 19576 18068 19582 18080
rect 20640 18068 20668 18108
rect 19576 18040 20668 18068
rect 21177 18071 21235 18077
rect 19576 18028 19582 18040
rect 21177 18037 21189 18071
rect 21223 18068 21235 18071
rect 21910 18068 21916 18080
rect 21223 18040 21916 18068
rect 21223 18037 21235 18040
rect 21177 18031 21235 18037
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 22012 18068 22040 18108
rect 24026 18096 24032 18148
rect 24084 18136 24090 18148
rect 31754 18136 31760 18148
rect 24084 18108 31760 18136
rect 24084 18096 24090 18108
rect 31754 18096 31760 18108
rect 31812 18096 31818 18148
rect 25314 18068 25320 18080
rect 22012 18040 25320 18068
rect 25314 18028 25320 18040
rect 25372 18028 25378 18080
rect 27062 18068 27068 18080
rect 27023 18040 27068 18068
rect 27062 18028 27068 18040
rect 27120 18028 27126 18080
rect 27246 18028 27252 18080
rect 27304 18068 27310 18080
rect 30834 18068 30840 18080
rect 27304 18040 30840 18068
rect 27304 18028 27310 18040
rect 30834 18028 30840 18040
rect 30892 18028 30898 18080
rect 1104 17978 44896 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 44896 17978
rect 1104 17904 44896 17926
rect 1578 17864 1584 17876
rect 1539 17836 1584 17864
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 1820 17836 3801 17864
rect 1820 17824 1826 17836
rect 3789 17833 3801 17836
rect 3835 17833 3847 17867
rect 6730 17864 6736 17876
rect 3789 17827 3847 17833
rect 4724 17836 6736 17864
rect 4724 17796 4752 17836
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 9858 17824 9864 17876
rect 9916 17864 9922 17876
rect 11054 17864 11060 17876
rect 9916 17836 11060 17864
rect 9916 17824 9922 17836
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 11238 17824 11244 17876
rect 11296 17864 11302 17876
rect 12066 17864 12072 17876
rect 11296 17836 12072 17864
rect 11296 17824 11302 17836
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 13170 17864 13176 17876
rect 12406 17836 13176 17864
rect 2976 17768 4752 17796
rect 6089 17799 6147 17805
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17728 1639 17731
rect 2222 17728 2228 17740
rect 1627 17700 2228 17728
rect 1627 17697 1639 17700
rect 1581 17691 1639 17697
rect 2222 17688 2228 17700
rect 2280 17688 2286 17740
rect 2976 17737 3004 17768
rect 6089 17765 6101 17799
rect 6135 17796 6147 17799
rect 6178 17796 6184 17808
rect 6135 17768 6184 17796
rect 6135 17765 6147 17768
rect 6089 17759 6147 17765
rect 6178 17756 6184 17768
rect 6236 17756 6242 17808
rect 6638 17756 6644 17808
rect 6696 17796 6702 17808
rect 12406 17796 12434 17836
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 13354 17824 13360 17876
rect 13412 17864 13418 17876
rect 14458 17864 14464 17876
rect 13412 17836 14464 17864
rect 13412 17824 13418 17836
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 14734 17824 14740 17876
rect 14792 17864 14798 17876
rect 16942 17864 16948 17876
rect 14792 17836 16948 17864
rect 14792 17824 14798 17836
rect 16942 17824 16948 17836
rect 17000 17824 17006 17876
rect 17126 17864 17132 17876
rect 17087 17836 17132 17864
rect 17126 17824 17132 17836
rect 17184 17824 17190 17876
rect 17402 17824 17408 17876
rect 17460 17864 17466 17876
rect 18414 17864 18420 17876
rect 17460 17836 18420 17864
rect 17460 17824 17466 17836
rect 18414 17824 18420 17836
rect 18472 17824 18478 17876
rect 18509 17867 18567 17873
rect 18509 17833 18521 17867
rect 18555 17864 18567 17867
rect 19150 17864 19156 17876
rect 18555 17836 19156 17864
rect 18555 17833 18567 17836
rect 18509 17827 18567 17833
rect 6696 17768 12434 17796
rect 15473 17799 15531 17805
rect 6696 17756 6702 17768
rect 15473 17765 15485 17799
rect 15519 17796 15531 17799
rect 18524 17796 18552 17827
rect 19150 17824 19156 17836
rect 19208 17824 19214 17876
rect 19242 17824 19248 17876
rect 19300 17864 19306 17876
rect 19518 17864 19524 17876
rect 19300 17836 19524 17864
rect 19300 17824 19306 17836
rect 19518 17824 19524 17836
rect 19576 17824 19582 17876
rect 20438 17864 20444 17876
rect 19727 17836 20444 17864
rect 15519 17768 18552 17796
rect 19613 17799 19671 17805
rect 15519 17765 15531 17768
rect 15473 17759 15531 17765
rect 19613 17765 19625 17799
rect 19659 17796 19671 17799
rect 19727 17796 19755 17836
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 20898 17864 20904 17876
rect 20859 17836 20904 17864
rect 20898 17824 20904 17836
rect 20956 17824 20962 17876
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 24397 17867 24455 17873
rect 24397 17864 24409 17867
rect 22244 17836 24409 17864
rect 22244 17824 22250 17836
rect 24397 17833 24409 17836
rect 24443 17833 24455 17867
rect 24397 17827 24455 17833
rect 25593 17867 25651 17873
rect 25593 17833 25605 17867
rect 25639 17864 25651 17867
rect 25682 17864 25688 17876
rect 25639 17836 25688 17864
rect 25639 17833 25651 17836
rect 25593 17827 25651 17833
rect 19659 17768 19755 17796
rect 19659 17765 19671 17768
rect 19613 17759 19671 17765
rect 19794 17756 19800 17808
rect 19852 17796 19858 17808
rect 20165 17799 20223 17805
rect 20165 17796 20177 17799
rect 19852 17768 20177 17796
rect 19852 17756 19858 17768
rect 20165 17765 20177 17768
rect 20211 17765 20223 17799
rect 21637 17799 21695 17805
rect 21637 17796 21649 17799
rect 20165 17759 20223 17765
rect 20272 17768 21649 17796
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17697 3019 17731
rect 3694 17728 3700 17740
rect 2961 17691 3019 17697
rect 3068 17700 3700 17728
rect 1394 17660 1400 17672
rect 1355 17632 1400 17660
rect 1394 17620 1400 17632
rect 1452 17620 1458 17672
rect 1670 17660 1676 17672
rect 1631 17632 1676 17660
rect 1670 17620 1676 17632
rect 1728 17620 1734 17672
rect 2866 17620 2872 17672
rect 2924 17660 2930 17672
rect 3068 17660 3096 17700
rect 3694 17688 3700 17700
rect 3752 17728 3758 17740
rect 3881 17731 3939 17737
rect 3881 17728 3893 17731
rect 3752 17700 3893 17728
rect 3752 17688 3758 17700
rect 3881 17697 3893 17700
rect 3927 17697 3939 17731
rect 3881 17691 3939 17697
rect 3988 17700 4568 17728
rect 2924 17632 3096 17660
rect 3237 17663 3295 17669
rect 2924 17620 2930 17632
rect 3237 17629 3249 17663
rect 3283 17660 3295 17663
rect 3988 17660 4016 17700
rect 3283 17632 4016 17660
rect 3283 17629 3295 17632
rect 3237 17623 3295 17629
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 4540 17660 4568 17700
rect 4614 17688 4620 17740
rect 4672 17728 4678 17740
rect 4709 17731 4767 17737
rect 4709 17728 4721 17731
rect 4672 17700 4721 17728
rect 4672 17688 4678 17700
rect 4709 17697 4721 17700
rect 4755 17697 4767 17731
rect 4709 17691 4767 17697
rect 5810 17688 5816 17740
rect 5868 17728 5874 17740
rect 6549 17731 6607 17737
rect 6549 17728 6561 17731
rect 5868 17700 6561 17728
rect 5868 17688 5874 17700
rect 6549 17697 6561 17700
rect 6595 17697 6607 17731
rect 6549 17691 6607 17697
rect 6730 17688 6736 17740
rect 6788 17728 6794 17740
rect 7009 17731 7067 17737
rect 7009 17728 7021 17731
rect 6788 17700 7021 17728
rect 6788 17688 6794 17700
rect 7009 17697 7021 17700
rect 7055 17697 7067 17731
rect 7009 17691 7067 17697
rect 7098 17688 7104 17740
rect 7156 17728 7162 17740
rect 10502 17728 10508 17740
rect 7156 17700 10508 17728
rect 7156 17688 7162 17700
rect 10502 17688 10508 17700
rect 10560 17728 10566 17740
rect 12158 17728 12164 17740
rect 10560 17700 12164 17728
rect 10560 17688 10566 17700
rect 12158 17688 12164 17700
rect 12216 17688 12222 17740
rect 12434 17728 12440 17740
rect 12395 17700 12440 17728
rect 12434 17688 12440 17700
rect 12492 17688 12498 17740
rect 12897 17731 12955 17737
rect 12897 17697 12909 17731
rect 12943 17728 12955 17731
rect 13630 17728 13636 17740
rect 12943 17700 13636 17728
rect 12943 17697 12955 17700
rect 12897 17691 12955 17697
rect 13630 17688 13636 17700
rect 13688 17688 13694 17740
rect 14090 17728 14096 17740
rect 14051 17700 14096 17728
rect 14090 17688 14096 17700
rect 14148 17688 14154 17740
rect 16114 17728 16120 17740
rect 16075 17700 16120 17728
rect 16114 17688 16120 17700
rect 16172 17728 16178 17740
rect 17218 17728 17224 17740
rect 16172 17700 17224 17728
rect 16172 17688 16178 17700
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17728 17831 17731
rect 17862 17728 17868 17740
rect 17819 17700 17868 17728
rect 17819 17697 17831 17700
rect 17773 17691 17831 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 18690 17728 18696 17740
rect 18432 17700 18696 17728
rect 5442 17660 5448 17672
rect 4120 17632 4165 17660
rect 4540 17632 5448 17660
rect 4120 17620 4126 17632
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 5534 17620 5540 17672
rect 5592 17620 5598 17672
rect 6178 17620 6184 17672
rect 6236 17660 6242 17672
rect 6454 17660 6460 17672
rect 6236 17632 6460 17660
rect 6236 17620 6242 17632
rect 6454 17620 6460 17632
rect 6512 17620 6518 17672
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 10870 17660 10876 17672
rect 10827 17632 10876 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13127 17632 13860 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 3050 17552 3056 17604
rect 3108 17592 3114 17604
rect 3326 17592 3332 17604
rect 3108 17564 3332 17592
rect 3108 17552 3114 17564
rect 3326 17552 3332 17564
rect 3384 17592 3390 17604
rect 3789 17595 3847 17601
rect 3789 17592 3801 17595
rect 3384 17564 3801 17592
rect 3384 17552 3390 17564
rect 3789 17561 3801 17564
rect 3835 17561 3847 17595
rect 4976 17595 5034 17601
rect 3789 17555 3847 17561
rect 3896 17564 4936 17592
rect 1854 17524 1860 17536
rect 1815 17496 1860 17524
rect 1854 17484 1860 17496
rect 1912 17484 1918 17536
rect 3694 17484 3700 17536
rect 3752 17524 3758 17536
rect 3896 17524 3924 17564
rect 3752 17496 3924 17524
rect 4249 17527 4307 17533
rect 3752 17484 3758 17496
rect 4249 17493 4261 17527
rect 4295 17524 4307 17527
rect 4798 17524 4804 17536
rect 4295 17496 4804 17524
rect 4295 17493 4307 17496
rect 4249 17487 4307 17493
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 4908 17524 4936 17564
rect 4976 17561 4988 17595
rect 5022 17592 5034 17595
rect 5074 17592 5080 17604
rect 5022 17564 5080 17592
rect 5022 17561 5034 17564
rect 4976 17555 5034 17561
rect 5074 17552 5080 17564
rect 5132 17552 5138 17604
rect 5552 17592 5580 17620
rect 6733 17595 6791 17601
rect 6733 17592 6745 17595
rect 5552 17564 6745 17592
rect 6733 17561 6745 17564
rect 6779 17561 6791 17595
rect 6733 17555 6791 17561
rect 7098 17552 7104 17604
rect 7156 17592 7162 17604
rect 7926 17592 7932 17604
rect 7156 17564 7932 17592
rect 7156 17552 7162 17564
rect 7926 17552 7932 17564
rect 7984 17552 7990 17604
rect 8941 17595 8999 17601
rect 8941 17561 8953 17595
rect 8987 17561 8999 17595
rect 8941 17555 8999 17561
rect 10597 17595 10655 17601
rect 10597 17561 10609 17595
rect 10643 17592 10655 17595
rect 11422 17592 11428 17604
rect 10643 17564 11428 17592
rect 10643 17561 10655 17564
rect 10597 17555 10655 17561
rect 8956 17524 8984 17555
rect 11422 17552 11428 17564
rect 11480 17552 11486 17604
rect 12342 17552 12348 17604
rect 12400 17592 12406 17604
rect 13354 17592 13360 17604
rect 12400 17564 13360 17592
rect 12400 17552 12406 17564
rect 13354 17552 13360 17564
rect 13412 17552 13418 17604
rect 13832 17592 13860 17632
rect 13906 17620 13912 17672
rect 13964 17660 13970 17672
rect 14349 17663 14407 17669
rect 14349 17660 14361 17663
rect 13964 17632 14361 17660
rect 13964 17620 13970 17632
rect 14349 17629 14361 17632
rect 14395 17629 14407 17663
rect 15654 17660 15660 17672
rect 14349 17623 14407 17629
rect 14476 17632 15660 17660
rect 14476 17592 14504 17632
rect 15654 17620 15660 17632
rect 15712 17660 15718 17672
rect 15838 17660 15844 17672
rect 15712 17632 15844 17660
rect 15712 17620 15718 17632
rect 15838 17620 15844 17632
rect 15896 17660 15902 17672
rect 17310 17660 17316 17672
rect 15896 17632 17316 17660
rect 15896 17620 15902 17632
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 17402 17620 17408 17672
rect 17460 17620 17466 17672
rect 17494 17620 17500 17672
rect 17552 17660 17558 17672
rect 18322 17660 18328 17672
rect 17552 17632 18328 17660
rect 17552 17620 17558 17632
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 16301 17595 16359 17601
rect 16301 17592 16313 17595
rect 13832 17564 14504 17592
rect 14568 17564 16313 17592
rect 4908 17496 8984 17524
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 14568 17524 14596 17564
rect 16301 17561 16313 17564
rect 16347 17561 16359 17595
rect 16301 17555 16359 17561
rect 17218 17552 17224 17604
rect 17276 17592 17282 17604
rect 17420 17592 17448 17620
rect 18432 17592 18460 17700
rect 18690 17688 18696 17700
rect 18748 17688 18754 17740
rect 18874 17688 18880 17740
rect 18932 17728 18938 17740
rect 18932 17700 19380 17728
rect 18932 17688 18938 17700
rect 19352 17660 19380 17700
rect 19518 17688 19524 17740
rect 19576 17728 19582 17740
rect 20272 17728 20300 17768
rect 21637 17765 21649 17768
rect 21683 17765 21695 17799
rect 21637 17759 21695 17765
rect 22557 17799 22615 17805
rect 22557 17765 22569 17799
rect 22603 17796 22615 17799
rect 22646 17796 22652 17808
rect 22603 17768 22652 17796
rect 22603 17765 22615 17768
rect 22557 17759 22615 17765
rect 22646 17756 22652 17768
rect 22704 17756 22710 17808
rect 23477 17799 23535 17805
rect 23477 17765 23489 17799
rect 23523 17796 23535 17799
rect 25608 17796 25636 17827
rect 25682 17824 25688 17836
rect 25740 17824 25746 17876
rect 26050 17864 26056 17876
rect 26011 17836 26056 17864
rect 26050 17824 26056 17836
rect 26108 17824 26114 17876
rect 27801 17867 27859 17873
rect 27801 17833 27813 17867
rect 27847 17864 27859 17867
rect 27890 17864 27896 17876
rect 27847 17836 27896 17864
rect 27847 17833 27859 17836
rect 27801 17827 27859 17833
rect 27890 17824 27896 17836
rect 27948 17824 27954 17876
rect 28258 17864 28264 17876
rect 28219 17836 28264 17864
rect 28258 17824 28264 17836
rect 28316 17824 28322 17876
rect 23523 17768 25636 17796
rect 23523 17765 23535 17768
rect 23477 17759 23535 17765
rect 19576 17700 20300 17728
rect 19576 17688 19582 17700
rect 21082 17688 21088 17740
rect 21140 17728 21146 17740
rect 22373 17731 22431 17737
rect 21140 17700 21864 17728
rect 21140 17688 21146 17700
rect 19794 17660 19800 17672
rect 19352 17654 19472 17660
rect 19536 17654 19800 17660
rect 19352 17632 19800 17654
rect 19444 17626 19564 17632
rect 19794 17620 19800 17632
rect 19852 17620 19858 17672
rect 19978 17620 19984 17672
rect 20036 17660 20042 17672
rect 20165 17663 20223 17669
rect 20165 17660 20177 17663
rect 20036 17632 20177 17660
rect 20036 17620 20042 17632
rect 20165 17629 20177 17632
rect 20211 17629 20223 17663
rect 20165 17623 20223 17629
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17660 20499 17663
rect 21177 17663 21235 17669
rect 20487 17632 21128 17660
rect 20487 17629 20499 17632
rect 20441 17623 20499 17629
rect 18506 17601 18512 17604
rect 17276 17564 17448 17592
rect 17972 17564 18460 17592
rect 18493 17595 18512 17601
rect 17276 17552 17282 17564
rect 17972 17536 18000 17564
rect 18493 17561 18505 17595
rect 18493 17555 18512 17561
rect 18506 17552 18512 17555
rect 18564 17552 18570 17604
rect 18693 17595 18751 17601
rect 18693 17561 18705 17595
rect 18739 17561 18751 17595
rect 18693 17555 18751 17561
rect 16206 17524 16212 17536
rect 9824 17496 14596 17524
rect 16167 17496 16212 17524
rect 9824 17484 9830 17496
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 16669 17527 16727 17533
rect 16669 17493 16681 17527
rect 16715 17524 16727 17527
rect 17310 17524 17316 17536
rect 16715 17496 17316 17524
rect 16715 17493 16727 17496
rect 16669 17487 16727 17493
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 17494 17524 17500 17536
rect 17455 17496 17500 17524
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 17589 17527 17647 17533
rect 17589 17493 17601 17527
rect 17635 17524 17647 17527
rect 17862 17524 17868 17536
rect 17635 17496 17868 17524
rect 17635 17493 17647 17496
rect 17589 17487 17647 17493
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 17954 17484 17960 17536
rect 18012 17484 18018 17536
rect 18046 17484 18052 17536
rect 18104 17524 18110 17536
rect 18325 17527 18383 17533
rect 18325 17524 18337 17527
rect 18104 17496 18337 17524
rect 18104 17484 18110 17496
rect 18325 17493 18337 17496
rect 18371 17493 18383 17527
rect 18708 17524 18736 17555
rect 18782 17552 18788 17604
rect 18840 17592 18846 17604
rect 19245 17595 19303 17601
rect 19245 17592 19257 17595
rect 18840 17564 19257 17592
rect 18840 17552 18846 17564
rect 19245 17561 19257 17564
rect 19291 17561 19303 17595
rect 20901 17595 20959 17601
rect 20901 17592 20913 17595
rect 19245 17555 19303 17561
rect 19352 17564 20913 17592
rect 18966 17524 18972 17536
rect 18708 17496 18972 17524
rect 18325 17487 18383 17493
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 19150 17484 19156 17536
rect 19208 17524 19214 17536
rect 19352 17524 19380 17564
rect 20901 17561 20913 17564
rect 20947 17561 20959 17595
rect 21100 17592 21128 17632
rect 21177 17629 21189 17663
rect 21223 17660 21235 17663
rect 21358 17660 21364 17672
rect 21223 17632 21364 17660
rect 21223 17629 21235 17632
rect 21177 17623 21235 17629
rect 21358 17620 21364 17632
rect 21416 17620 21422 17672
rect 21836 17669 21864 17700
rect 22373 17697 22385 17731
rect 22419 17728 22431 17731
rect 22922 17728 22928 17740
rect 22419 17700 22928 17728
rect 22419 17697 22431 17700
rect 22373 17691 22431 17697
rect 22922 17688 22928 17700
rect 22980 17688 22986 17740
rect 23293 17731 23351 17737
rect 23293 17697 23305 17731
rect 23339 17728 23351 17731
rect 25130 17728 25136 17740
rect 23339 17700 25136 17728
rect 23339 17697 23351 17700
rect 23293 17691 23351 17697
rect 25130 17688 25136 17700
rect 25188 17688 25194 17740
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17629 21879 17663
rect 26605 17663 26663 17669
rect 26605 17660 26617 17663
rect 21821 17623 21879 17629
rect 22756 17632 26617 17660
rect 21726 17592 21732 17604
rect 21100 17564 21732 17592
rect 20901 17555 20959 17561
rect 21726 17552 21732 17564
rect 21784 17552 21790 17604
rect 19208 17496 19380 17524
rect 19705 17527 19763 17533
rect 19208 17484 19214 17496
rect 19705 17493 19717 17527
rect 19751 17524 19763 17527
rect 20254 17524 20260 17536
rect 19751 17496 20260 17524
rect 19751 17493 19763 17496
rect 19705 17487 19763 17493
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 20349 17527 20407 17533
rect 20349 17493 20361 17527
rect 20395 17524 20407 17527
rect 20530 17524 20536 17536
rect 20395 17496 20536 17524
rect 20395 17493 20407 17496
rect 20349 17487 20407 17493
rect 20530 17484 20536 17496
rect 20588 17484 20594 17536
rect 20990 17484 20996 17536
rect 21048 17524 21054 17536
rect 21085 17527 21143 17533
rect 21085 17524 21097 17527
rect 21048 17496 21097 17524
rect 21048 17484 21054 17496
rect 21085 17493 21097 17496
rect 21131 17493 21143 17527
rect 21085 17487 21143 17493
rect 21358 17484 21364 17536
rect 21416 17524 21422 17536
rect 22756 17524 22784 17632
rect 26605 17629 26617 17632
rect 26651 17660 26663 17663
rect 27062 17660 27068 17672
rect 26651 17632 27068 17660
rect 26651 17629 26663 17632
rect 26605 17623 26663 17629
rect 27062 17620 27068 17632
rect 27120 17660 27126 17672
rect 27157 17663 27215 17669
rect 27157 17660 27169 17663
rect 27120 17632 27169 17660
rect 27120 17620 27126 17632
rect 27157 17629 27169 17632
rect 27203 17660 27215 17663
rect 27246 17660 27252 17672
rect 27203 17632 27252 17660
rect 27203 17629 27215 17632
rect 27157 17623 27215 17629
rect 27246 17620 27252 17632
rect 27304 17620 27310 17672
rect 22833 17595 22891 17601
rect 22833 17561 22845 17595
rect 22879 17592 22891 17595
rect 23014 17592 23020 17604
rect 22879 17564 23020 17592
rect 22879 17561 22891 17564
rect 22833 17555 22891 17561
rect 23014 17552 23020 17564
rect 23072 17592 23078 17604
rect 23753 17595 23811 17601
rect 23753 17592 23765 17595
rect 23072 17564 23765 17592
rect 23072 17552 23078 17564
rect 23753 17561 23765 17564
rect 23799 17561 23811 17595
rect 23753 17555 23811 17561
rect 21416 17496 22784 17524
rect 21416 17484 21422 17496
rect 23198 17484 23204 17536
rect 23256 17524 23262 17536
rect 23566 17524 23572 17536
rect 23256 17496 23572 17524
rect 23256 17484 23262 17496
rect 23566 17484 23572 17496
rect 23624 17484 23630 17536
rect 24946 17524 24952 17536
rect 24907 17496 24952 17524
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 28997 17527 29055 17533
rect 28997 17493 29009 17527
rect 29043 17524 29055 17527
rect 29178 17524 29184 17536
rect 29043 17496 29184 17524
rect 29043 17493 29055 17496
rect 28997 17487 29055 17493
rect 29178 17484 29184 17496
rect 29236 17484 29242 17536
rect 29825 17527 29883 17533
rect 29825 17493 29837 17527
rect 29871 17524 29883 17527
rect 29914 17524 29920 17536
rect 29871 17496 29920 17524
rect 29871 17493 29883 17496
rect 29825 17487 29883 17493
rect 29914 17484 29920 17496
rect 29972 17484 29978 17536
rect 1104 17434 44896 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 44896 17434
rect 1104 17360 44896 17382
rect 1765 17323 1823 17329
rect 1765 17289 1777 17323
rect 1811 17320 1823 17323
rect 2774 17320 2780 17332
rect 1811 17292 2780 17320
rect 1811 17289 1823 17292
rect 1765 17283 1823 17289
rect 2774 17280 2780 17292
rect 2832 17320 2838 17332
rect 3694 17320 3700 17332
rect 2832 17292 3700 17320
rect 2832 17280 2838 17292
rect 3694 17280 3700 17292
rect 3752 17280 3758 17332
rect 3973 17323 4031 17329
rect 3973 17289 3985 17323
rect 4019 17320 4031 17323
rect 5626 17320 5632 17332
rect 4019 17292 5632 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 5626 17280 5632 17292
rect 5684 17280 5690 17332
rect 5718 17280 5724 17332
rect 5776 17320 5782 17332
rect 5813 17323 5871 17329
rect 5813 17320 5825 17323
rect 5776 17292 5825 17320
rect 5776 17280 5782 17292
rect 5813 17289 5825 17292
rect 5859 17289 5871 17323
rect 5813 17283 5871 17289
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 10594 17320 10600 17332
rect 5960 17292 10600 17320
rect 5960 17280 5966 17292
rect 10594 17280 10600 17292
rect 10652 17280 10658 17332
rect 12250 17320 12256 17332
rect 11532 17292 12256 17320
rect 2860 17255 2918 17261
rect 2860 17221 2872 17255
rect 2906 17252 2918 17255
rect 3878 17252 3884 17264
rect 2906 17224 3884 17252
rect 2906 17221 2918 17224
rect 2860 17215 2918 17221
rect 3878 17212 3884 17224
rect 3936 17212 3942 17264
rect 4154 17212 4160 17264
rect 4212 17252 4218 17264
rect 4678 17255 4736 17261
rect 4678 17252 4690 17255
rect 4212 17224 4690 17252
rect 4212 17212 4218 17224
rect 4678 17221 4690 17224
rect 4724 17221 4736 17255
rect 4678 17215 4736 17221
rect 4798 17212 4804 17264
rect 4856 17252 4862 17264
rect 9125 17255 9183 17261
rect 9125 17252 9137 17255
rect 4856 17224 9137 17252
rect 4856 17212 4862 17224
rect 9125 17221 9137 17224
rect 9171 17221 9183 17255
rect 9125 17215 9183 17221
rect 10686 17212 10692 17264
rect 10744 17252 10750 17264
rect 11532 17261 11560 17292
rect 12250 17280 12256 17292
rect 12308 17320 12314 17332
rect 17494 17320 17500 17332
rect 12308 17292 17500 17320
rect 12308 17280 12314 17292
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 18598 17280 18604 17332
rect 18656 17320 18662 17332
rect 22278 17320 22284 17332
rect 18656 17292 22284 17320
rect 18656 17280 18662 17292
rect 22278 17280 22284 17292
rect 22336 17280 22342 17332
rect 23109 17323 23167 17329
rect 23109 17289 23121 17323
rect 23155 17320 23167 17323
rect 24026 17320 24032 17332
rect 23155 17292 24032 17320
rect 23155 17289 23167 17292
rect 23109 17283 23167 17289
rect 24026 17280 24032 17292
rect 24084 17280 24090 17332
rect 28626 17280 28632 17332
rect 28684 17320 28690 17332
rect 41598 17320 41604 17332
rect 28684 17292 41604 17320
rect 28684 17280 28690 17292
rect 41598 17280 41604 17292
rect 41656 17280 41662 17332
rect 10781 17255 10839 17261
rect 10781 17252 10793 17255
rect 10744 17224 10793 17252
rect 10744 17212 10750 17224
rect 10781 17221 10793 17224
rect 10827 17221 10839 17255
rect 10781 17215 10839 17221
rect 11517 17255 11575 17261
rect 11517 17221 11529 17255
rect 11563 17221 11575 17255
rect 11517 17215 11575 17221
rect 11790 17212 11796 17264
rect 11848 17252 11854 17264
rect 12342 17252 12348 17264
rect 11848 17224 12348 17252
rect 11848 17212 11854 17224
rect 12342 17212 12348 17224
rect 12400 17212 12406 17264
rect 13170 17252 13176 17264
rect 13131 17224 13176 17252
rect 13170 17212 13176 17224
rect 13228 17212 13234 17264
rect 14182 17212 14188 17264
rect 14240 17252 14246 17264
rect 14338 17255 14396 17261
rect 14338 17252 14350 17255
rect 14240 17224 14350 17252
rect 14240 17212 14246 17224
rect 14338 17221 14350 17224
rect 14384 17221 14396 17255
rect 17954 17252 17960 17264
rect 14338 17215 14396 17221
rect 16040 17224 17960 17252
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 2314 17144 2320 17196
rect 2372 17184 2378 17196
rect 2590 17184 2596 17196
rect 2372 17156 2596 17184
rect 2372 17144 2378 17156
rect 2590 17144 2596 17156
rect 2648 17144 2654 17196
rect 4430 17184 4436 17196
rect 4391 17156 4436 17184
rect 4430 17144 4436 17156
rect 4488 17144 4494 17196
rect 4540 17156 5488 17184
rect 750 17076 756 17128
rect 808 17116 814 17128
rect 1489 17119 1547 17125
rect 1489 17116 1501 17119
rect 808 17088 1501 17116
rect 808 17076 814 17088
rect 1489 17085 1501 17088
rect 1535 17085 1547 17119
rect 1489 17079 1547 17085
rect 3970 17076 3976 17128
rect 4028 17116 4034 17128
rect 4540 17116 4568 17156
rect 4028 17088 4568 17116
rect 5460 17116 5488 17156
rect 6086 17144 6092 17196
rect 6144 17184 6150 17196
rect 6457 17187 6515 17193
rect 6457 17184 6469 17187
rect 6144 17156 6469 17184
rect 6144 17144 6150 17156
rect 6457 17153 6469 17156
rect 6503 17153 6515 17187
rect 7098 17184 7104 17196
rect 7059 17156 7104 17184
rect 6457 17147 6515 17153
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 7190 17144 7196 17196
rect 7248 17144 7254 17196
rect 7368 17187 7426 17193
rect 7368 17153 7380 17187
rect 7414 17184 7426 17187
rect 8478 17184 8484 17196
rect 7414 17156 8484 17184
rect 7414 17153 7426 17156
rect 7368 17147 7426 17153
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 8846 17144 8852 17196
rect 8904 17150 8910 17196
rect 14090 17184 14096 17196
rect 14051 17156 14096 17184
rect 8904 17144 8972 17150
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 14200 17156 15240 17184
rect 7208 17116 7236 17144
rect 8864 17125 8972 17144
rect 8864 17122 8999 17125
rect 5460 17088 7236 17116
rect 8941 17119 8999 17122
rect 4028 17076 4034 17088
rect 8941 17085 8953 17119
rect 8987 17085 8999 17119
rect 8941 17079 8999 17085
rect 9122 17076 9128 17128
rect 9180 17116 9186 17128
rect 9858 17116 9864 17128
rect 9180 17088 9864 17116
rect 9180 17076 9186 17088
rect 9858 17076 9864 17088
rect 9916 17076 9922 17128
rect 13357 17119 13415 17125
rect 13357 17085 13369 17119
rect 13403 17116 13415 17119
rect 13814 17116 13820 17128
rect 13403 17088 13820 17116
rect 13403 17085 13415 17088
rect 13357 17079 13415 17085
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 14200 17116 14228 17156
rect 14108 17088 14228 17116
rect 2130 17048 2136 17060
rect 2091 17020 2136 17048
rect 2130 17008 2136 17020
rect 2188 17008 2194 17060
rect 8481 17051 8539 17057
rect 8481 17017 8493 17051
rect 8527 17048 8539 17051
rect 12434 17048 12440 17060
rect 8527 17020 12440 17048
rect 8527 17017 8539 17020
rect 8481 17011 8539 17017
rect 12434 17008 12440 17020
rect 12492 17008 12498 17060
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 14108 17048 14136 17088
rect 12584 17020 14136 17048
rect 15212 17048 15240 17156
rect 15286 17076 15292 17128
rect 15344 17116 15350 17128
rect 16040 17125 16068 17224
rect 17954 17212 17960 17224
rect 18012 17252 18018 17264
rect 18417 17255 18475 17261
rect 18417 17252 18429 17255
rect 18012 17224 18429 17252
rect 18012 17212 18018 17224
rect 18417 17221 18429 17224
rect 18463 17221 18475 17255
rect 18417 17215 18475 17221
rect 18782 17212 18788 17264
rect 18840 17252 18846 17264
rect 19337 17255 19395 17261
rect 18840 17224 19196 17252
rect 18840 17212 18846 17224
rect 16666 17184 16672 17196
rect 16627 17156 16672 17184
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 16758 17144 16764 17196
rect 16816 17184 16822 17196
rect 16945 17187 17003 17193
rect 16945 17184 16957 17187
rect 16816 17156 16957 17184
rect 16816 17144 16822 17156
rect 16945 17153 16957 17156
rect 16991 17153 17003 17187
rect 16945 17147 17003 17153
rect 17218 17144 17224 17196
rect 17276 17184 17282 17196
rect 18101 17187 18159 17193
rect 18101 17184 18113 17187
rect 17276 17156 18113 17184
rect 17276 17144 17282 17156
rect 18101 17153 18113 17156
rect 18147 17153 18159 17187
rect 18101 17147 18159 17153
rect 18233 17187 18291 17193
rect 18233 17153 18245 17187
rect 18279 17184 18291 17187
rect 18506 17184 18512 17196
rect 18279 17156 18512 17184
rect 18279 17153 18291 17156
rect 18233 17147 18291 17153
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 19061 17187 19119 17193
rect 19061 17184 19073 17187
rect 18800 17156 19073 17184
rect 18800 17128 18828 17156
rect 19061 17153 19073 17156
rect 19107 17153 19119 17187
rect 19168 17184 19196 17224
rect 19337 17221 19349 17255
rect 19383 17252 19395 17255
rect 19978 17252 19984 17264
rect 19383 17224 19984 17252
rect 19383 17221 19395 17224
rect 19337 17215 19395 17221
rect 19978 17212 19984 17224
rect 20036 17212 20042 17264
rect 20438 17212 20444 17264
rect 20496 17252 20502 17264
rect 20625 17255 20683 17261
rect 20625 17252 20637 17255
rect 20496 17224 20637 17252
rect 20496 17212 20502 17224
rect 20625 17221 20637 17224
rect 20671 17252 20683 17255
rect 26145 17255 26203 17261
rect 26145 17252 26157 17255
rect 20671 17224 26157 17252
rect 20671 17221 20683 17224
rect 20625 17215 20683 17221
rect 26145 17221 26157 17224
rect 26191 17221 26203 17255
rect 28077 17255 28135 17261
rect 28077 17252 28089 17255
rect 26145 17215 26203 17221
rect 27586 17224 28089 17252
rect 21266 17184 21272 17196
rect 19168 17156 20576 17184
rect 21227 17156 21272 17184
rect 19061 17147 19119 17153
rect 20548 17128 20576 17156
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 21726 17144 21732 17196
rect 21784 17184 21790 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21784 17156 22017 17184
rect 21784 17144 21790 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22097 17187 22155 17193
rect 22097 17153 22109 17187
rect 22143 17153 22155 17187
rect 22097 17147 22155 17153
rect 22281 17187 22339 17193
rect 22281 17153 22293 17187
rect 22327 17184 22339 17187
rect 22554 17184 22560 17196
rect 22327 17156 22560 17184
rect 22327 17153 22339 17156
rect 22281 17147 22339 17153
rect 16025 17119 16083 17125
rect 16025 17116 16037 17119
rect 15344 17088 16037 17116
rect 15344 17076 15350 17088
rect 16025 17085 16037 17088
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 18782 17076 18788 17128
rect 18840 17076 18846 17128
rect 19245 17119 19303 17125
rect 19245 17085 19257 17119
rect 19291 17116 19303 17119
rect 19610 17116 19616 17128
rect 19291 17088 19616 17116
rect 19291 17085 19303 17088
rect 19245 17079 19303 17085
rect 19610 17076 19616 17088
rect 19668 17076 19674 17128
rect 19794 17076 19800 17128
rect 19852 17116 19858 17128
rect 20165 17119 20223 17125
rect 20165 17116 20177 17119
rect 19852 17088 20177 17116
rect 19852 17076 19858 17088
rect 20165 17085 20177 17088
rect 20211 17085 20223 17119
rect 20165 17079 20223 17085
rect 20346 17076 20352 17128
rect 20404 17076 20410 17128
rect 20530 17076 20536 17128
rect 20588 17116 20594 17128
rect 22112 17116 22140 17147
rect 22554 17144 22560 17156
rect 22612 17144 22618 17196
rect 23474 17144 23480 17196
rect 23532 17184 23538 17196
rect 27586 17184 27614 17224
rect 28077 17221 28089 17224
rect 28123 17221 28135 17255
rect 28077 17215 28135 17221
rect 28994 17212 29000 17264
rect 29052 17252 29058 17264
rect 43898 17252 43904 17264
rect 29052 17224 43904 17252
rect 29052 17212 29058 17224
rect 43898 17212 43904 17224
rect 43956 17212 43962 17264
rect 23532 17156 27614 17184
rect 23532 17144 23538 17156
rect 27890 17144 27896 17196
rect 27948 17184 27954 17196
rect 28629 17187 28687 17193
rect 28629 17184 28641 17187
rect 27948 17156 28641 17184
rect 27948 17144 27954 17156
rect 28629 17153 28641 17156
rect 28675 17184 28687 17187
rect 29638 17184 29644 17196
rect 28675 17156 29644 17184
rect 28675 17153 28687 17156
rect 28629 17147 28687 17153
rect 29638 17144 29644 17156
rect 29696 17144 29702 17196
rect 23198 17116 23204 17128
rect 20588 17088 23204 17116
rect 20588 17076 20594 17088
rect 23198 17076 23204 17088
rect 23256 17076 23262 17128
rect 23569 17119 23627 17125
rect 23569 17085 23581 17119
rect 23615 17085 23627 17119
rect 23569 17079 23627 17085
rect 17957 17051 18015 17057
rect 17957 17048 17969 17051
rect 15212 17020 17969 17048
rect 12584 17008 12590 17020
rect 17957 17017 17969 17020
rect 18003 17017 18015 17051
rect 17957 17011 18015 17017
rect 18322 17008 18328 17060
rect 18380 17048 18386 17060
rect 18877 17051 18935 17057
rect 18877 17048 18889 17051
rect 18380 17020 18889 17048
rect 18380 17008 18386 17020
rect 18877 17017 18889 17020
rect 18923 17017 18935 17051
rect 20257 17051 20315 17057
rect 18877 17011 18935 17017
rect 19168 17020 20208 17048
rect 474 16940 480 16992
rect 532 16980 538 16992
rect 750 16980 756 16992
rect 532 16952 756 16980
rect 532 16940 538 16952
rect 750 16940 756 16952
rect 808 16940 814 16992
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 5718 16980 5724 16992
rect 3384 16952 5724 16980
rect 3384 16940 3390 16952
rect 5718 16940 5724 16952
rect 5776 16980 5782 16992
rect 5902 16980 5908 16992
rect 5776 16952 5908 16980
rect 5776 16940 5782 16952
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 6546 16980 6552 16992
rect 6052 16952 6552 16980
rect 6052 16940 6058 16952
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 6730 16940 6736 16992
rect 6788 16980 6794 16992
rect 10410 16980 10416 16992
rect 6788 16952 10416 16980
rect 6788 16940 6794 16952
rect 10410 16940 10416 16952
rect 10468 16940 10474 16992
rect 10594 16940 10600 16992
rect 10652 16980 10658 16992
rect 15286 16980 15292 16992
rect 10652 16952 15292 16980
rect 10652 16940 10658 16952
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 15473 16983 15531 16989
rect 15473 16949 15485 16983
rect 15519 16980 15531 16983
rect 16390 16980 16396 16992
rect 15519 16952 16396 16980
rect 15519 16949 15531 16952
rect 15473 16943 15531 16949
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 18417 16983 18475 16989
rect 18417 16980 18429 16983
rect 16724 16952 18429 16980
rect 16724 16940 16730 16952
rect 18417 16949 18429 16952
rect 18463 16980 18475 16983
rect 18506 16980 18512 16992
rect 18463 16952 18512 16980
rect 18463 16949 18475 16952
rect 18417 16943 18475 16949
rect 18506 16940 18512 16952
rect 18564 16940 18570 16992
rect 18966 16940 18972 16992
rect 19024 16980 19030 16992
rect 19168 16980 19196 17020
rect 19334 16980 19340 16992
rect 19024 16952 19196 16980
rect 19295 16952 19340 16980
rect 19024 16940 19030 16952
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 20180 16980 20208 17020
rect 20257 17017 20269 17051
rect 20303 17048 20315 17051
rect 20364 17048 20392 17076
rect 20303 17020 20392 17048
rect 21085 17051 21143 17057
rect 20303 17017 20315 17020
rect 20257 17011 20315 17017
rect 21085 17017 21097 17051
rect 21131 17048 21143 17051
rect 21174 17048 21180 17060
rect 21131 17020 21180 17048
rect 21131 17017 21143 17020
rect 21085 17011 21143 17017
rect 21174 17008 21180 17020
rect 21232 17048 21238 17060
rect 23293 17051 23351 17057
rect 21232 17020 22968 17048
rect 21232 17008 21238 17020
rect 22940 16992 22968 17020
rect 23293 17017 23305 17051
rect 23339 17048 23351 17051
rect 23382 17048 23388 17060
rect 23339 17020 23388 17048
rect 23339 17017 23351 17020
rect 23293 17011 23351 17017
rect 23382 17008 23388 17020
rect 23440 17008 23446 17060
rect 23584 17048 23612 17079
rect 24118 17076 24124 17128
rect 24176 17116 24182 17128
rect 24673 17119 24731 17125
rect 24673 17116 24685 17119
rect 24176 17088 24685 17116
rect 24176 17076 24182 17088
rect 24673 17085 24685 17088
rect 24719 17085 24731 17119
rect 24673 17079 24731 17085
rect 24762 17076 24768 17128
rect 24820 17116 24826 17128
rect 25593 17119 25651 17125
rect 25593 17116 25605 17119
rect 24820 17088 25605 17116
rect 24820 17076 24826 17088
rect 25593 17085 25605 17088
rect 25639 17085 25651 17119
rect 25593 17079 25651 17085
rect 29270 17076 29276 17128
rect 29328 17116 29334 17128
rect 30374 17116 30380 17128
rect 29328 17088 30380 17116
rect 29328 17076 29334 17088
rect 30374 17076 30380 17088
rect 30432 17076 30438 17128
rect 23492 17020 23612 17048
rect 25041 17051 25099 17057
rect 20990 16980 20996 16992
rect 20180 16952 20996 16980
rect 20990 16940 20996 16952
rect 21048 16980 21054 16992
rect 22186 16980 22192 16992
rect 21048 16952 22192 16980
rect 21048 16940 21054 16952
rect 22186 16940 22192 16952
rect 22244 16940 22250 16992
rect 22281 16983 22339 16989
rect 22281 16949 22293 16983
rect 22327 16980 22339 16983
rect 22646 16980 22652 16992
rect 22327 16952 22652 16980
rect 22327 16949 22339 16952
rect 22281 16943 22339 16949
rect 22646 16940 22652 16952
rect 22704 16940 22710 16992
rect 22922 16940 22928 16992
rect 22980 16940 22986 16992
rect 23014 16940 23020 16992
rect 23072 16980 23078 16992
rect 23492 16980 23520 17020
rect 25041 17017 25053 17051
rect 25087 17048 25099 17051
rect 26050 17048 26056 17060
rect 25087 17020 26056 17048
rect 25087 17017 25099 17020
rect 25041 17011 25099 17017
rect 26050 17008 26056 17020
rect 26108 17008 26114 17060
rect 24026 16980 24032 16992
rect 23072 16952 23520 16980
rect 23987 16952 24032 16980
rect 23072 16940 23078 16952
rect 24026 16940 24032 16952
rect 24084 16940 24090 16992
rect 25133 16983 25191 16989
rect 25133 16949 25145 16983
rect 25179 16980 25191 16983
rect 25406 16980 25412 16992
rect 25179 16952 25412 16980
rect 25179 16949 25191 16952
rect 25133 16943 25191 16949
rect 25406 16940 25412 16952
rect 25464 16940 25470 16992
rect 26970 16980 26976 16992
rect 26931 16952 26976 16980
rect 26970 16940 26976 16952
rect 27028 16940 27034 16992
rect 27617 16983 27675 16989
rect 27617 16949 27629 16983
rect 27663 16980 27675 16983
rect 28902 16980 28908 16992
rect 27663 16952 28908 16980
rect 27663 16949 27675 16952
rect 27617 16943 27675 16949
rect 28902 16940 28908 16952
rect 28960 16940 28966 16992
rect 29086 16940 29092 16992
rect 29144 16980 29150 16992
rect 37918 16980 37924 16992
rect 29144 16952 37924 16980
rect 29144 16940 29150 16952
rect 37918 16940 37924 16952
rect 37976 16940 37982 16992
rect 1104 16890 44896 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 44896 16890
rect 1104 16816 44896 16838
rect 1762 16776 1768 16788
rect 1723 16748 1768 16776
rect 1762 16736 1768 16748
rect 1820 16736 1826 16788
rect 2866 16776 2872 16788
rect 1872 16748 2872 16776
rect 1394 16600 1400 16652
rect 1452 16640 1458 16652
rect 1673 16643 1731 16649
rect 1673 16640 1685 16643
rect 1452 16612 1685 16640
rect 1452 16600 1458 16612
rect 1673 16609 1685 16612
rect 1719 16640 1731 16643
rect 1872 16640 1900 16748
rect 2866 16736 2872 16748
rect 2924 16736 2930 16788
rect 6730 16776 6736 16788
rect 5460 16748 6736 16776
rect 1949 16711 2007 16717
rect 1949 16677 1961 16711
rect 1995 16708 2007 16711
rect 1995 16680 2452 16708
rect 1995 16677 2007 16680
rect 1949 16671 2007 16677
rect 2424 16649 2452 16680
rect 1719 16612 1900 16640
rect 2409 16643 2467 16649
rect 1719 16609 1731 16612
rect 1673 16603 1731 16609
rect 2409 16609 2421 16643
rect 2455 16609 2467 16643
rect 2409 16603 2467 16609
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16640 4399 16643
rect 4706 16640 4712 16652
rect 4387 16612 4712 16640
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 1578 16532 1584 16584
rect 1636 16572 1642 16584
rect 1765 16575 1823 16581
rect 1765 16572 1777 16575
rect 1636 16544 1777 16572
rect 1636 16532 1642 16544
rect 1765 16541 1777 16544
rect 1811 16572 1823 16575
rect 3970 16572 3976 16584
rect 1811 16544 3976 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16572 4675 16575
rect 5460 16572 5488 16748
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 7098 16776 7104 16788
rect 6932 16748 7104 16776
rect 6932 16649 6960 16748
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 7248 16748 7972 16776
rect 7248 16736 7254 16748
rect 6457 16643 6515 16649
rect 6457 16609 6469 16643
rect 6503 16640 6515 16643
rect 6917 16643 6975 16649
rect 6917 16640 6929 16643
rect 6503 16612 6929 16640
rect 6503 16609 6515 16612
rect 6457 16603 6515 16609
rect 6917 16609 6929 16612
rect 6963 16609 6975 16643
rect 7944 16640 7972 16748
rect 8478 16736 8484 16788
rect 8536 16776 8542 16788
rect 9122 16776 9128 16788
rect 8536 16748 9128 16776
rect 8536 16736 8542 16748
rect 9122 16736 9128 16748
rect 9180 16736 9186 16788
rect 13630 16776 13636 16788
rect 11348 16748 13636 16776
rect 8202 16668 8208 16720
rect 8260 16708 8266 16720
rect 10134 16708 10140 16720
rect 8260 16680 10140 16708
rect 8260 16668 8266 16680
rect 10134 16668 10140 16680
rect 10192 16708 10198 16720
rect 10870 16708 10876 16720
rect 10192 16680 10876 16708
rect 10192 16668 10198 16680
rect 10870 16668 10876 16680
rect 10928 16668 10934 16720
rect 9033 16643 9091 16649
rect 9033 16640 9045 16643
rect 7944 16612 9045 16640
rect 6917 16603 6975 16609
rect 9033 16609 9045 16612
rect 9079 16640 9091 16643
rect 9306 16640 9312 16652
rect 9079 16612 9312 16640
rect 9079 16609 9091 16612
rect 9033 16603 9091 16609
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 9766 16640 9772 16652
rect 9727 16612 9772 16640
rect 9766 16600 9772 16612
rect 9824 16600 9830 16652
rect 11348 16649 11376 16748
rect 13630 16736 13636 16748
rect 13688 16736 13694 16788
rect 14366 16776 14372 16788
rect 14108 16748 14372 16776
rect 14108 16708 14136 16748
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 16666 16776 16672 16788
rect 14476 16748 16672 16776
rect 13096 16680 14136 16708
rect 14185 16711 14243 16717
rect 11333 16643 11391 16649
rect 11333 16609 11345 16643
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 11514 16600 11520 16652
rect 11572 16640 11578 16652
rect 11793 16643 11851 16649
rect 11793 16640 11805 16643
rect 11572 16612 11805 16640
rect 11572 16600 11578 16612
rect 11793 16609 11805 16612
rect 11839 16640 11851 16643
rect 11839 16612 12204 16640
rect 11839 16609 11851 16612
rect 11793 16603 11851 16609
rect 4663 16544 5488 16572
rect 6201 16575 6259 16581
rect 4663 16541 4675 16544
rect 4617 16535 4675 16541
rect 6201 16541 6213 16575
rect 6247 16572 6259 16575
rect 6822 16572 6828 16584
rect 6247 16544 6828 16572
rect 6247 16541 6259 16544
rect 6201 16535 6259 16541
rect 6822 16532 6828 16544
rect 6880 16532 6886 16584
rect 7184 16575 7242 16581
rect 7184 16541 7196 16575
rect 7230 16572 7242 16575
rect 7466 16572 7472 16584
rect 7230 16544 7472 16572
rect 7230 16541 7242 16544
rect 7184 16535 7242 16541
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 12066 16572 12072 16584
rect 12027 16544 12072 16572
rect 12066 16532 12072 16544
rect 12124 16532 12130 16584
rect 12176 16572 12204 16612
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 13096 16640 13124 16680
rect 14185 16677 14197 16711
rect 14231 16708 14243 16711
rect 14476 16708 14504 16748
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 17678 16736 17684 16788
rect 17736 16776 17742 16788
rect 18230 16776 18236 16788
rect 17736 16748 18236 16776
rect 17736 16736 17742 16748
rect 18230 16736 18236 16748
rect 18288 16736 18294 16788
rect 18782 16736 18788 16788
rect 18840 16736 18846 16788
rect 19334 16736 19340 16788
rect 19392 16776 19398 16788
rect 19429 16779 19487 16785
rect 19429 16776 19441 16779
rect 19392 16748 19441 16776
rect 19392 16736 19398 16748
rect 19429 16745 19441 16748
rect 19475 16745 19487 16779
rect 19429 16739 19487 16745
rect 19702 16736 19708 16788
rect 19760 16776 19766 16788
rect 20162 16776 20168 16788
rect 19760 16748 20168 16776
rect 19760 16736 19766 16748
rect 20162 16736 20168 16748
rect 20220 16736 20226 16788
rect 20625 16779 20683 16785
rect 20625 16745 20637 16779
rect 20671 16776 20683 16779
rect 20898 16776 20904 16788
rect 20671 16748 20904 16776
rect 20671 16745 20683 16748
rect 20625 16739 20683 16745
rect 20898 16736 20904 16748
rect 20956 16736 20962 16788
rect 23198 16736 23204 16788
rect 23256 16776 23262 16788
rect 25866 16776 25872 16788
rect 23256 16748 25636 16776
rect 25827 16748 25872 16776
rect 23256 16736 23262 16748
rect 14231 16680 14504 16708
rect 14231 16677 14243 16680
rect 14185 16671 14243 16677
rect 12492 16612 13124 16640
rect 12492 16600 12498 16612
rect 13170 16600 13176 16652
rect 13228 16640 13234 16652
rect 14200 16640 14228 16671
rect 13228 16612 14228 16640
rect 14645 16643 14703 16649
rect 13228 16600 13234 16612
rect 14645 16609 14657 16643
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 12986 16572 12992 16584
rect 12176 16544 12992 16572
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 14660 16572 14688 16603
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 16577 16643 16635 16649
rect 16577 16640 16589 16643
rect 16448 16612 16589 16640
rect 16448 16600 16454 16612
rect 16577 16609 16589 16612
rect 16623 16609 16635 16643
rect 16577 16603 16635 16609
rect 16666 16600 16672 16652
rect 16724 16640 16730 16652
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 16724 16612 16865 16640
rect 16724 16600 16730 16612
rect 16853 16609 16865 16612
rect 16899 16609 16911 16643
rect 16853 16603 16911 16609
rect 17586 16600 17592 16652
rect 17644 16640 17650 16652
rect 17865 16643 17923 16649
rect 17865 16640 17877 16643
rect 17644 16612 17877 16640
rect 17644 16600 17650 16612
rect 17865 16609 17877 16612
rect 17911 16609 17923 16643
rect 18138 16640 18144 16652
rect 18099 16612 18144 16640
rect 17865 16603 17923 16609
rect 18138 16600 18144 16612
rect 18196 16600 18202 16652
rect 18800 16640 18828 16736
rect 19150 16668 19156 16720
rect 19208 16708 19214 16720
rect 21361 16711 21419 16717
rect 21361 16708 21373 16711
rect 19208 16680 21373 16708
rect 19208 16668 19214 16680
rect 21361 16677 21373 16680
rect 21407 16677 21419 16711
rect 21361 16671 21419 16677
rect 22373 16711 22431 16717
rect 22373 16677 22385 16711
rect 22419 16708 22431 16711
rect 22462 16708 22468 16720
rect 22419 16680 22468 16708
rect 22419 16677 22431 16680
rect 22373 16671 22431 16677
rect 22462 16668 22468 16680
rect 22520 16668 22526 16720
rect 23477 16711 23535 16717
rect 23477 16677 23489 16711
rect 23523 16708 23535 16711
rect 24670 16708 24676 16720
rect 23523 16680 24676 16708
rect 23523 16677 23535 16680
rect 23477 16671 23535 16677
rect 24670 16668 24676 16680
rect 24728 16668 24734 16720
rect 25409 16711 25467 16717
rect 25409 16677 25421 16711
rect 25455 16708 25467 16711
rect 25498 16708 25504 16720
rect 25455 16680 25504 16708
rect 25455 16677 25467 16680
rect 25409 16671 25467 16677
rect 25498 16668 25504 16680
rect 25556 16668 25562 16720
rect 25608 16708 25636 16748
rect 25866 16736 25872 16748
rect 25924 16736 25930 16788
rect 27614 16776 27620 16788
rect 25976 16748 27620 16776
rect 25976 16708 26004 16748
rect 27614 16736 27620 16748
rect 27672 16736 27678 16788
rect 28169 16779 28227 16785
rect 28169 16745 28181 16779
rect 28215 16776 28227 16779
rect 28350 16776 28356 16788
rect 28215 16748 28356 16776
rect 28215 16745 28227 16748
rect 28169 16739 28227 16745
rect 28350 16736 28356 16748
rect 28408 16776 28414 16788
rect 28629 16779 28687 16785
rect 28629 16776 28641 16779
rect 28408 16748 28641 16776
rect 28408 16736 28414 16748
rect 28629 16745 28641 16748
rect 28675 16745 28687 16779
rect 28629 16739 28687 16745
rect 27062 16708 27068 16720
rect 25608 16680 26004 16708
rect 27023 16680 27068 16708
rect 27062 16668 27068 16680
rect 27120 16668 27126 16720
rect 29546 16708 29552 16720
rect 29507 16680 29552 16708
rect 29546 16668 29552 16680
rect 29604 16668 29610 16720
rect 19610 16640 19616 16652
rect 18800 16612 19472 16640
rect 19571 16612 19616 16640
rect 14734 16572 14740 16584
rect 14660 16544 14740 16572
rect 14734 16532 14740 16544
rect 14792 16532 14798 16584
rect 14918 16581 14924 16584
rect 14912 16535 14924 16581
rect 14976 16572 14982 16584
rect 14976 16544 15012 16572
rect 14918 16532 14924 16535
rect 14976 16532 14982 16544
rect 16482 16532 16488 16584
rect 16540 16572 16546 16584
rect 18322 16572 18328 16584
rect 16540 16544 18328 16572
rect 16540 16532 16546 16544
rect 18322 16532 18328 16544
rect 18380 16532 18386 16584
rect 19444 16581 19472 16612
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 20162 16600 20168 16652
rect 20220 16640 20226 16652
rect 20441 16643 20499 16649
rect 20441 16640 20453 16643
rect 20220 16612 20453 16640
rect 20220 16600 20226 16612
rect 20441 16609 20453 16612
rect 20487 16640 20499 16643
rect 21266 16640 21272 16652
rect 20487 16612 21272 16640
rect 20487 16609 20499 16612
rect 20441 16603 20499 16609
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 21542 16600 21548 16652
rect 21600 16640 21606 16652
rect 21600 16612 21645 16640
rect 21600 16600 21606 16612
rect 22094 16600 22100 16652
rect 22152 16640 22158 16652
rect 22554 16640 22560 16652
rect 22152 16612 22560 16640
rect 22152 16600 22158 16612
rect 22554 16600 22560 16612
rect 22612 16600 22618 16652
rect 22922 16600 22928 16652
rect 22980 16640 22986 16652
rect 24489 16643 24547 16649
rect 24489 16640 24501 16643
rect 22980 16612 24501 16640
rect 22980 16600 22986 16612
rect 24489 16609 24501 16612
rect 24535 16640 24547 16643
rect 25038 16640 25044 16652
rect 24535 16612 25044 16640
rect 24535 16609 24547 16612
rect 24489 16603 24547 16609
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 27617 16643 27675 16649
rect 27617 16640 27629 16643
rect 25240 16612 27629 16640
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16572 19763 16575
rect 19978 16572 19984 16584
rect 19751 16544 19984 16572
rect 19751 16541 19763 16544
rect 19705 16535 19763 16541
rect 1489 16507 1547 16513
rect 1489 16473 1501 16507
rect 1535 16504 1547 16507
rect 3326 16504 3332 16516
rect 1535 16476 3332 16504
rect 1535 16473 1547 16476
rect 1489 16467 1547 16473
rect 3326 16464 3332 16476
rect 3384 16464 3390 16516
rect 5442 16504 5448 16516
rect 3712 16476 5448 16504
rect 2639 16439 2697 16445
rect 2639 16405 2651 16439
rect 2685 16436 2697 16439
rect 3712 16436 3740 16476
rect 5442 16464 5448 16476
rect 5500 16464 5506 16516
rect 5626 16464 5632 16516
rect 5684 16504 5690 16516
rect 10226 16504 10232 16516
rect 5684 16476 10232 16504
rect 5684 16464 5690 16476
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 11149 16507 11207 16513
rect 11149 16473 11161 16507
rect 11195 16504 11207 16507
rect 11606 16504 11612 16516
rect 11195 16476 11612 16504
rect 11195 16473 11207 16476
rect 11149 16467 11207 16473
rect 11606 16464 11612 16476
rect 11664 16464 11670 16516
rect 15470 16464 15476 16516
rect 15528 16504 15534 16516
rect 15838 16504 15844 16516
rect 15528 16476 15844 16504
rect 15528 16464 15534 16476
rect 15838 16464 15844 16476
rect 15896 16464 15902 16516
rect 17862 16504 17868 16516
rect 16040 16476 17868 16504
rect 2685 16408 3740 16436
rect 2685 16405 2697 16408
rect 2639 16399 2697 16405
rect 3786 16396 3792 16448
rect 3844 16436 3850 16448
rect 5077 16439 5135 16445
rect 5077 16436 5089 16439
rect 3844 16408 5089 16436
rect 3844 16396 3850 16408
rect 5077 16405 5089 16408
rect 5123 16405 5135 16439
rect 5077 16399 5135 16405
rect 7374 16396 7380 16448
rect 7432 16436 7438 16448
rect 8202 16436 8208 16448
rect 7432 16408 8208 16436
rect 7432 16396 7438 16408
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 8297 16439 8355 16445
rect 8297 16405 8309 16439
rect 8343 16436 8355 16439
rect 8846 16436 8852 16448
rect 8343 16408 8852 16436
rect 8343 16405 8355 16408
rect 8297 16399 8355 16405
rect 8846 16396 8852 16408
rect 8904 16396 8910 16448
rect 13170 16436 13176 16448
rect 13131 16408 13176 16436
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 16040 16445 16068 16476
rect 17862 16464 17868 16476
rect 17920 16504 17926 16516
rect 19334 16504 19340 16516
rect 17920 16476 19340 16504
rect 17920 16464 17926 16476
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 19444 16504 19472 16535
rect 19978 16532 19984 16544
rect 20036 16532 20042 16584
rect 20254 16532 20260 16584
rect 20312 16572 20318 16584
rect 20349 16575 20407 16581
rect 20349 16572 20361 16575
rect 20312 16544 20361 16572
rect 20312 16532 20318 16544
rect 20349 16541 20361 16544
rect 20395 16541 20407 16575
rect 21174 16572 21180 16584
rect 20349 16535 20407 16541
rect 20456 16544 21180 16572
rect 20456 16504 20484 16544
rect 21174 16532 21180 16544
rect 21232 16532 21238 16584
rect 23290 16572 23296 16584
rect 23251 16544 23296 16572
rect 23290 16532 23296 16544
rect 23348 16532 23354 16584
rect 25240 16516 25268 16612
rect 27617 16609 27629 16612
rect 27663 16609 27675 16643
rect 27617 16603 27675 16609
rect 20622 16504 20628 16516
rect 19444 16476 20484 16504
rect 20583 16476 20628 16504
rect 20622 16464 20628 16476
rect 20680 16464 20686 16516
rect 21085 16507 21143 16513
rect 21085 16473 21097 16507
rect 21131 16504 21143 16507
rect 22002 16504 22008 16516
rect 21131 16476 22008 16504
rect 21131 16473 21143 16476
rect 21085 16467 21143 16473
rect 22002 16464 22008 16476
rect 22060 16464 22066 16516
rect 25222 16504 25228 16516
rect 22388 16476 24440 16504
rect 25183 16476 25228 16504
rect 16025 16439 16083 16445
rect 16025 16436 16037 16439
rect 13872 16408 16037 16436
rect 13872 16396 13878 16408
rect 16025 16405 16037 16408
rect 16071 16405 16083 16439
rect 16025 16399 16083 16405
rect 16114 16396 16120 16448
rect 16172 16436 16178 16448
rect 18598 16436 18604 16448
rect 16172 16408 18604 16436
rect 16172 16396 16178 16408
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 18690 16396 18696 16448
rect 18748 16436 18754 16448
rect 19245 16439 19303 16445
rect 19245 16436 19257 16439
rect 18748 16408 19257 16436
rect 18748 16396 18754 16408
rect 19245 16405 19257 16408
rect 19291 16405 19303 16439
rect 19245 16399 19303 16405
rect 20165 16439 20223 16445
rect 20165 16405 20177 16439
rect 20211 16436 20223 16439
rect 20254 16436 20260 16448
rect 20211 16408 20260 16436
rect 20211 16405 20223 16408
rect 20165 16399 20223 16405
rect 20254 16396 20260 16408
rect 20312 16396 20318 16448
rect 21266 16396 21272 16448
rect 21324 16436 21330 16448
rect 22388 16436 22416 16476
rect 21324 16408 22416 16436
rect 22465 16439 22523 16445
rect 21324 16396 21330 16408
rect 22465 16405 22477 16439
rect 22511 16436 22523 16439
rect 23290 16436 23296 16448
rect 22511 16408 23296 16436
rect 22511 16405 22523 16408
rect 22465 16399 22523 16405
rect 23290 16396 23296 16408
rect 23348 16396 23354 16448
rect 24412 16436 24440 16476
rect 25222 16464 25228 16476
rect 25280 16464 25286 16516
rect 26418 16436 26424 16448
rect 24412 16408 26424 16436
rect 26418 16396 26424 16408
rect 26476 16396 26482 16448
rect 1104 16346 44896 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 44896 16346
rect 1104 16272 44896 16294
rect 1670 16232 1676 16244
rect 1631 16204 1676 16232
rect 1670 16192 1676 16204
rect 1728 16192 1734 16244
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 3973 16235 4031 16241
rect 3973 16201 3985 16235
rect 4019 16201 4031 16235
rect 3973 16195 4031 16201
rect 842 16124 848 16176
rect 900 16164 906 16176
rect 2838 16167 2896 16173
rect 2838 16164 2850 16167
rect 900 16136 2850 16164
rect 900 16124 906 16136
rect 2838 16133 2850 16136
rect 2884 16133 2896 16167
rect 3988 16164 4016 16195
rect 4062 16192 4068 16244
rect 4120 16232 4126 16244
rect 4120 16204 8800 16232
rect 4120 16192 4126 16204
rect 5258 16164 5264 16176
rect 3988 16136 5264 16164
rect 2838 16127 2896 16133
rect 5258 16124 5264 16136
rect 5316 16124 5322 16176
rect 7926 16124 7932 16176
rect 7984 16164 7990 16176
rect 7984 16136 8708 16164
rect 7984 16124 7990 16136
rect 1302 16056 1308 16108
rect 1360 16096 1366 16108
rect 1765 16099 1823 16105
rect 1765 16096 1777 16099
rect 1360 16068 1777 16096
rect 1360 16056 1366 16068
rect 1765 16065 1777 16068
rect 1811 16096 1823 16099
rect 2590 16096 2596 16108
rect 1811 16068 2452 16096
rect 2551 16068 2596 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 2424 15892 2452 16068
rect 2590 16056 2596 16068
rect 2648 16056 2654 16108
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16096 4491 16099
rect 4522 16096 4528 16108
rect 4479 16068 4528 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 4522 16056 4528 16068
rect 4580 16056 4586 16108
rect 4700 16099 4758 16105
rect 4700 16065 4712 16099
rect 4746 16096 4758 16099
rect 5166 16096 5172 16108
rect 4746 16068 5172 16096
rect 4746 16065 4758 16068
rect 4700 16059 4758 16065
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 6454 16096 6460 16108
rect 6415 16068 6460 16096
rect 6454 16056 6460 16068
rect 6512 16056 6518 16108
rect 6549 16099 6607 16105
rect 6549 16065 6561 16099
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 8409 16099 8467 16105
rect 8409 16065 8421 16099
rect 8455 16096 8467 16099
rect 8570 16096 8576 16108
rect 8455 16068 8576 16096
rect 8455 16065 8467 16068
rect 8409 16059 8467 16065
rect 5813 15963 5871 15969
rect 5813 15929 5825 15963
rect 5859 15960 5871 15963
rect 6362 15960 6368 15972
rect 5859 15932 6368 15960
rect 5859 15929 5871 15932
rect 5813 15923 5871 15929
rect 6362 15920 6368 15932
rect 6420 15920 6426 15972
rect 6564 15960 6592 16059
rect 8570 16056 8576 16068
rect 8628 16056 8634 16108
rect 8680 16105 8708 16136
rect 8665 16099 8723 16105
rect 8665 16065 8677 16099
rect 8711 16065 8723 16099
rect 8772 16096 8800 16204
rect 9398 16192 9404 16244
rect 9456 16232 9462 16244
rect 11330 16232 11336 16244
rect 9456 16204 11336 16232
rect 9456 16192 9462 16204
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 11606 16232 11612 16244
rect 11567 16204 11612 16232
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 15749 16235 15807 16241
rect 15749 16232 15761 16235
rect 12452 16204 15761 16232
rect 8938 16124 8944 16176
rect 8996 16164 9002 16176
rect 8996 16136 11376 16164
rect 8996 16124 9002 16136
rect 9122 16096 9128 16108
rect 8772 16068 9128 16096
rect 8665 16059 8723 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 11348 16096 11376 16136
rect 12452 16096 12480 16204
rect 15749 16201 15761 16204
rect 15795 16201 15807 16235
rect 16666 16232 16672 16244
rect 16627 16204 16672 16232
rect 15749 16195 15807 16201
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 16942 16192 16948 16244
rect 17000 16232 17006 16244
rect 20898 16232 20904 16244
rect 17000 16204 20904 16232
rect 17000 16192 17006 16204
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 21818 16232 21824 16244
rect 21779 16204 21824 16232
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 23474 16232 23480 16244
rect 21928 16204 23480 16232
rect 12744 16167 12802 16173
rect 12744 16133 12756 16167
rect 12790 16164 12802 16167
rect 13078 16164 13084 16176
rect 12790 16136 13084 16164
rect 12790 16133 12802 16136
rect 12744 16127 12802 16133
rect 13078 16124 13084 16136
rect 13136 16124 13142 16176
rect 14090 16124 14096 16176
rect 14148 16164 14154 16176
rect 17770 16164 17776 16176
rect 17828 16173 17834 16176
rect 14148 16136 14964 16164
rect 17740 16136 17776 16164
rect 14148 16124 14154 16136
rect 12986 16096 12992 16108
rect 11348 16068 12480 16096
rect 12899 16068 12992 16096
rect 12986 16056 12992 16068
rect 13044 16096 13050 16108
rect 14108 16096 14136 16124
rect 13044 16068 14136 16096
rect 14665 16099 14723 16105
rect 13044 16056 13050 16068
rect 14665 16065 14677 16099
rect 14711 16096 14723 16099
rect 14826 16096 14832 16108
rect 14711 16068 14832 16096
rect 14711 16065 14723 16068
rect 14665 16059 14723 16065
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 14936 16105 14964 16136
rect 17770 16124 17776 16136
rect 17828 16127 17840 16173
rect 19242 16164 19248 16176
rect 18064 16136 19248 16164
rect 17828 16124 17834 16127
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 15838 16096 15844 16108
rect 15703 16068 15844 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 15838 16056 15844 16068
rect 15896 16096 15902 16108
rect 16114 16096 16120 16108
rect 15896 16068 16120 16096
rect 15896 16056 15902 16068
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 17954 16056 17960 16108
rect 18012 16096 18018 16108
rect 18064 16105 18092 16136
rect 19242 16124 19248 16136
rect 19300 16124 19306 16176
rect 20070 16124 20076 16176
rect 20128 16164 20134 16176
rect 20165 16167 20223 16173
rect 20165 16164 20177 16167
rect 20128 16136 20177 16164
rect 20128 16124 20134 16136
rect 20165 16133 20177 16136
rect 20211 16133 20223 16167
rect 21450 16164 21456 16176
rect 20165 16127 20223 16133
rect 20272 16136 21456 16164
rect 18049 16099 18107 16105
rect 18049 16096 18061 16099
rect 18012 16068 18061 16096
rect 18012 16056 18018 16068
rect 18049 16065 18061 16068
rect 18095 16065 18107 16099
rect 18874 16096 18880 16108
rect 18835 16068 18880 16096
rect 18049 16059 18107 16065
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 19886 16096 19892 16108
rect 19847 16068 19892 16096
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 20036 16068 20081 16096
rect 20036 16056 20042 16068
rect 10778 16028 10784 16040
rect 10739 16000 10784 16028
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 15997 11023 16031
rect 15470 16028 15476 16040
rect 15431 16000 15476 16028
rect 10965 15991 11023 15997
rect 6564 15932 7788 15960
rect 3878 15892 3884 15904
rect 2424 15864 3884 15892
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 6733 15895 6791 15901
rect 6733 15861 6745 15895
rect 6779 15892 6791 15895
rect 6914 15892 6920 15904
rect 6779 15864 6920 15892
rect 6779 15861 6791 15864
rect 6733 15855 6791 15861
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 7374 15892 7380 15904
rect 7331 15864 7380 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 7760 15892 7788 15932
rect 10134 15892 10140 15904
rect 7760 15864 10140 15892
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 10980 15892 11008 15991
rect 15470 15988 15476 16000
rect 15528 15988 15534 16040
rect 18598 16028 18604 16040
rect 18559 16000 18604 16028
rect 18598 15988 18604 16000
rect 18656 15988 18662 16040
rect 18785 16031 18843 16037
rect 18785 15997 18797 16031
rect 18831 16028 18843 16031
rect 19058 16028 19064 16040
rect 18831 16000 19064 16028
rect 18831 15997 18843 16000
rect 18785 15991 18843 15997
rect 19058 15988 19064 16000
rect 19116 16028 19122 16040
rect 20272 16028 20300 16136
rect 21450 16124 21456 16136
rect 21508 16164 21514 16176
rect 21928 16164 21956 16204
rect 23474 16192 23480 16204
rect 23532 16192 23538 16244
rect 23661 16235 23719 16241
rect 23661 16201 23673 16235
rect 23707 16232 23719 16235
rect 24394 16232 24400 16244
rect 23707 16204 24400 16232
rect 23707 16201 23719 16204
rect 23661 16195 23719 16201
rect 24394 16192 24400 16204
rect 24452 16192 24458 16244
rect 25038 16232 25044 16244
rect 24999 16204 25044 16232
rect 25038 16192 25044 16204
rect 25096 16192 25102 16244
rect 25314 16192 25320 16244
rect 25372 16232 25378 16244
rect 25593 16235 25651 16241
rect 25593 16232 25605 16235
rect 25372 16204 25605 16232
rect 25372 16192 25378 16204
rect 25593 16201 25605 16204
rect 25639 16232 25651 16235
rect 26786 16232 26792 16244
rect 25639 16204 26792 16232
rect 25639 16201 25651 16204
rect 25593 16195 25651 16201
rect 26786 16192 26792 16204
rect 26844 16192 26850 16244
rect 27614 16232 27620 16244
rect 27575 16204 27620 16232
rect 27614 16192 27620 16204
rect 27672 16232 27678 16244
rect 30377 16235 30435 16241
rect 30377 16232 30389 16235
rect 27672 16204 30389 16232
rect 27672 16192 27678 16204
rect 30377 16201 30389 16204
rect 30423 16201 30435 16235
rect 30377 16195 30435 16201
rect 21508 16136 21956 16164
rect 21508 16124 21514 16136
rect 22830 16124 22836 16176
rect 22888 16164 22894 16176
rect 23198 16164 23204 16176
rect 22888 16136 23204 16164
rect 22888 16124 22894 16136
rect 23198 16124 23204 16136
rect 23256 16124 23262 16176
rect 23290 16124 23296 16176
rect 23348 16164 23354 16176
rect 26145 16167 26203 16173
rect 23348 16136 24532 16164
rect 23348 16124 23354 16136
rect 20530 16056 20536 16108
rect 20588 16096 20594 16108
rect 20809 16099 20867 16105
rect 20588 16068 20668 16096
rect 20588 16056 20594 16068
rect 20640 16037 20668 16068
rect 20809 16065 20821 16099
rect 20855 16096 20867 16099
rect 20855 16068 21496 16096
rect 20855 16065 20867 16068
rect 20809 16059 20867 16065
rect 19116 16000 20300 16028
rect 20625 16031 20683 16037
rect 19116 15988 19122 16000
rect 20625 15997 20637 16031
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 20990 15988 20996 16040
rect 21048 16028 21054 16040
rect 21085 16031 21143 16037
rect 21085 16028 21097 16031
rect 21048 16000 21097 16028
rect 21048 15988 21054 16000
rect 21085 15997 21097 16000
rect 21131 15997 21143 16031
rect 21468 16028 21496 16068
rect 21542 16056 21548 16108
rect 21600 16096 21606 16108
rect 24504 16105 24532 16136
rect 26145 16133 26157 16167
rect 26191 16164 26203 16167
rect 26326 16164 26332 16176
rect 26191 16136 26332 16164
rect 26191 16133 26203 16136
rect 26145 16127 26203 16133
rect 26326 16124 26332 16136
rect 26384 16124 26390 16176
rect 23845 16099 23903 16105
rect 23845 16096 23857 16099
rect 21600 16068 23857 16096
rect 21600 16056 21606 16068
rect 23845 16065 23857 16068
rect 23891 16065 23903 16099
rect 23845 16059 23903 16065
rect 24489 16099 24547 16105
rect 24489 16065 24501 16099
rect 24535 16065 24547 16099
rect 24489 16059 24547 16065
rect 24946 16056 24952 16108
rect 25004 16096 25010 16108
rect 26970 16096 26976 16108
rect 25004 16068 26976 16096
rect 25004 16056 25010 16068
rect 26970 16056 26976 16068
rect 27028 16056 27034 16108
rect 22281 16031 22339 16037
rect 21468 16000 22094 16028
rect 21085 15991 21143 15997
rect 16117 15963 16175 15969
rect 16117 15929 16129 15963
rect 16163 15960 16175 15963
rect 16163 15932 17172 15960
rect 16163 15929 16175 15932
rect 16117 15923 16175 15929
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 10980 15864 13553 15892
rect 13541 15861 13553 15864
rect 13587 15892 13599 15895
rect 16482 15892 16488 15904
rect 13587 15864 16488 15892
rect 13587 15861 13599 15864
rect 13541 15855 13599 15861
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 17144 15892 17172 15932
rect 19150 15920 19156 15972
rect 19208 15960 19214 15972
rect 19245 15963 19303 15969
rect 19245 15960 19257 15963
rect 19208 15932 19257 15960
rect 19208 15920 19214 15932
rect 19245 15929 19257 15932
rect 19291 15929 19303 15963
rect 19245 15923 19303 15929
rect 19426 15920 19432 15972
rect 19484 15960 19490 15972
rect 19705 15963 19763 15969
rect 19705 15960 19717 15963
rect 19484 15932 19717 15960
rect 19484 15920 19490 15932
rect 19705 15929 19717 15932
rect 19751 15929 19763 15963
rect 19705 15923 19763 15929
rect 20088 15932 20668 15960
rect 17770 15892 17776 15904
rect 17144 15864 17776 15892
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 18414 15852 18420 15904
rect 18472 15892 18478 15904
rect 20088 15892 20116 15932
rect 18472 15864 20116 15892
rect 20165 15895 20223 15901
rect 18472 15852 18478 15864
rect 20165 15861 20177 15895
rect 20211 15892 20223 15895
rect 20530 15892 20536 15904
rect 20211 15864 20536 15892
rect 20211 15861 20223 15864
rect 20165 15855 20223 15861
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 20640 15892 20668 15932
rect 20714 15920 20720 15972
rect 20772 15960 20778 15972
rect 21913 15963 21971 15969
rect 21913 15960 21925 15963
rect 20772 15932 21925 15960
rect 20772 15920 20778 15932
rect 21913 15929 21925 15932
rect 21959 15929 21971 15963
rect 22066 15960 22094 16000
rect 22281 15997 22293 16031
rect 22327 16028 22339 16031
rect 22327 16000 22692 16028
rect 22327 15997 22339 16000
rect 22281 15991 22339 15997
rect 22554 15960 22560 15972
rect 22066 15932 22560 15960
rect 21913 15923 21971 15929
rect 22554 15920 22560 15932
rect 22612 15920 22618 15972
rect 20993 15895 21051 15901
rect 20993 15892 21005 15895
rect 20640 15864 21005 15892
rect 20993 15861 21005 15864
rect 21039 15892 21051 15895
rect 21174 15892 21180 15904
rect 21039 15864 21180 15892
rect 21039 15861 21051 15864
rect 20993 15855 21051 15861
rect 21174 15852 21180 15864
rect 21232 15852 21238 15904
rect 22664 15892 22692 16000
rect 22738 15988 22744 16040
rect 22796 16028 22802 16040
rect 22796 16000 22841 16028
rect 22796 15988 22802 16000
rect 24026 15988 24032 16040
rect 24084 16028 24090 16040
rect 29181 16031 29239 16037
rect 29181 16028 29193 16031
rect 24084 16000 29193 16028
rect 24084 15988 24090 16000
rect 29181 15997 29193 16000
rect 29227 15997 29239 16031
rect 29181 15991 29239 15997
rect 22925 15963 22983 15969
rect 22925 15929 22937 15963
rect 22971 15960 22983 15963
rect 23750 15960 23756 15972
rect 22971 15932 23756 15960
rect 22971 15929 22983 15932
rect 22925 15923 22983 15929
rect 23750 15920 23756 15932
rect 23808 15920 23814 15972
rect 24302 15960 24308 15972
rect 24263 15932 24308 15960
rect 24302 15920 24308 15932
rect 24360 15920 24366 15972
rect 24854 15960 24860 15972
rect 24412 15932 24860 15960
rect 24412 15892 24440 15932
rect 24854 15920 24860 15932
rect 24912 15960 24918 15972
rect 29733 15963 29791 15969
rect 29733 15960 29745 15963
rect 24912 15932 29745 15960
rect 24912 15920 24918 15932
rect 29733 15929 29745 15932
rect 29779 15929 29791 15963
rect 29733 15923 29791 15929
rect 22664 15864 24440 15892
rect 24670 15852 24676 15904
rect 24728 15892 24734 15904
rect 26602 15892 26608 15904
rect 24728 15864 26608 15892
rect 24728 15852 24734 15864
rect 26602 15852 26608 15864
rect 26660 15892 26666 15904
rect 28077 15895 28135 15901
rect 28077 15892 28089 15895
rect 26660 15864 28089 15892
rect 26660 15852 26666 15864
rect 28077 15861 28089 15864
rect 28123 15861 28135 15895
rect 28626 15892 28632 15904
rect 28587 15864 28632 15892
rect 28077 15855 28135 15861
rect 28626 15852 28632 15864
rect 28684 15852 28690 15904
rect 1104 15802 44896 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 44896 15802
rect 1104 15728 44896 15750
rect 1762 15688 1768 15700
rect 1675 15660 1768 15688
rect 1762 15648 1768 15660
rect 1820 15688 1826 15700
rect 2130 15688 2136 15700
rect 1820 15660 2136 15688
rect 1820 15648 1826 15660
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 3878 15648 3884 15700
rect 3936 15688 3942 15700
rect 3936 15660 9260 15688
rect 3936 15648 3942 15660
rect 750 15580 756 15632
rect 808 15620 814 15632
rect 1949 15623 2007 15629
rect 808 15592 1900 15620
rect 808 15580 814 15592
rect 1394 15512 1400 15564
rect 1452 15552 1458 15564
rect 1581 15555 1639 15561
rect 1581 15552 1593 15555
rect 1452 15524 1593 15552
rect 1452 15512 1458 15524
rect 1581 15521 1593 15524
rect 1627 15521 1639 15555
rect 1872 15552 1900 15592
rect 1949 15589 1961 15623
rect 1995 15620 2007 15623
rect 4982 15620 4988 15632
rect 1995 15592 4988 15620
rect 1995 15589 2007 15592
rect 1949 15583 2007 15589
rect 4982 15580 4988 15592
rect 5040 15580 5046 15632
rect 8297 15623 8355 15629
rect 8297 15589 8309 15623
rect 8343 15620 8355 15623
rect 8754 15620 8760 15632
rect 8343 15592 8760 15620
rect 8343 15589 8355 15592
rect 8297 15583 8355 15589
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 2409 15555 2467 15561
rect 2409 15552 2421 15555
rect 1872 15524 2421 15552
rect 1581 15515 1639 15521
rect 2409 15521 2421 15524
rect 2455 15521 2467 15555
rect 4614 15552 4620 15564
rect 4575 15524 4620 15552
rect 2409 15515 2467 15521
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 9232 15561 9260 15660
rect 13630 15648 13636 15700
rect 13688 15688 13694 15700
rect 14185 15691 14243 15697
rect 14185 15688 14197 15691
rect 13688 15660 14197 15688
rect 13688 15648 13694 15660
rect 14185 15657 14197 15660
rect 14231 15688 14243 15691
rect 14458 15688 14464 15700
rect 14231 15660 14464 15688
rect 14231 15657 14243 15660
rect 14185 15651 14243 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 14884 15660 17172 15688
rect 14884 15648 14890 15660
rect 9217 15555 9275 15561
rect 9217 15521 9229 15555
rect 9263 15521 9275 15555
rect 10870 15552 10876 15564
rect 10831 15524 10876 15552
rect 9217 15515 9275 15521
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15552 11115 15555
rect 11606 15552 11612 15564
rect 11103 15524 11612 15552
rect 11103 15521 11115 15524
rect 11057 15515 11115 15521
rect 11606 15512 11612 15524
rect 11664 15512 11670 15564
rect 13265 15555 13323 15561
rect 13265 15521 13277 15555
rect 13311 15552 13323 15555
rect 13722 15552 13728 15564
rect 13311 15524 13728 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 13722 15512 13728 15524
rect 13780 15512 13786 15564
rect 17144 15552 17172 15660
rect 18138 15648 18144 15700
rect 18196 15688 18202 15700
rect 19705 15691 19763 15697
rect 18196 15660 19656 15688
rect 18196 15648 18202 15660
rect 17218 15580 17224 15632
rect 17276 15620 17282 15632
rect 19242 15620 19248 15632
rect 17276 15592 18000 15620
rect 19203 15592 19248 15620
rect 17276 15580 17282 15592
rect 17865 15555 17923 15561
rect 17865 15552 17877 15555
rect 17144 15524 17877 15552
rect 17865 15521 17877 15524
rect 17911 15521 17923 15555
rect 17972 15552 18000 15592
rect 19242 15580 19248 15592
rect 19300 15580 19306 15632
rect 19628 15620 19656 15660
rect 19705 15657 19717 15691
rect 19751 15688 19763 15691
rect 20530 15688 20536 15700
rect 19751 15660 20536 15688
rect 19751 15657 19763 15660
rect 19705 15651 19763 15657
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 20625 15691 20683 15697
rect 20625 15657 20637 15691
rect 20671 15657 20683 15691
rect 20625 15651 20683 15657
rect 21361 15691 21419 15697
rect 21361 15657 21373 15691
rect 21407 15688 21419 15691
rect 21542 15688 21548 15700
rect 21407 15660 21441 15688
rect 21503 15660 21548 15688
rect 21407 15657 21419 15660
rect 21361 15651 21419 15657
rect 20640 15620 20668 15651
rect 20898 15620 20904 15632
rect 19628 15592 20208 15620
rect 20640 15592 20904 15620
rect 20180 15564 20208 15592
rect 20898 15580 20904 15592
rect 20956 15620 20962 15632
rect 21376 15620 21404 15651
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 23661 15691 23719 15697
rect 23661 15688 23673 15691
rect 21652 15660 23673 15688
rect 21652 15632 21680 15660
rect 23661 15657 23673 15660
rect 23707 15688 23719 15691
rect 24946 15688 24952 15700
rect 23707 15660 24952 15688
rect 23707 15657 23719 15660
rect 23661 15651 23719 15657
rect 24946 15648 24952 15660
rect 25004 15648 25010 15700
rect 25777 15691 25835 15697
rect 25777 15657 25789 15691
rect 25823 15688 25835 15691
rect 26142 15688 26148 15700
rect 25823 15660 26148 15688
rect 25823 15657 25835 15660
rect 25777 15651 25835 15657
rect 26142 15648 26148 15660
rect 26200 15648 26206 15700
rect 26326 15688 26332 15700
rect 26287 15660 26332 15688
rect 26326 15648 26332 15660
rect 26384 15648 26390 15700
rect 26786 15688 26792 15700
rect 26747 15660 26792 15688
rect 26786 15648 26792 15660
rect 26844 15648 26850 15700
rect 26970 15648 26976 15700
rect 27028 15688 27034 15700
rect 27341 15691 27399 15697
rect 27341 15688 27353 15691
rect 27028 15660 27353 15688
rect 27028 15648 27034 15660
rect 27341 15657 27353 15660
rect 27387 15657 27399 15691
rect 27341 15651 27399 15657
rect 29362 15648 29368 15700
rect 29420 15688 29426 15700
rect 29549 15691 29607 15697
rect 29549 15688 29561 15691
rect 29420 15660 29561 15688
rect 29420 15648 29426 15660
rect 29549 15657 29561 15660
rect 29595 15657 29607 15691
rect 29549 15651 29607 15657
rect 29638 15648 29644 15700
rect 29696 15688 29702 15700
rect 30101 15691 30159 15697
rect 30101 15688 30113 15691
rect 29696 15660 30113 15688
rect 29696 15648 29702 15660
rect 30101 15657 30113 15660
rect 30147 15657 30159 15691
rect 30101 15651 30159 15657
rect 21634 15620 21640 15632
rect 20956 15592 21640 15620
rect 20956 15580 20962 15592
rect 21634 15580 21640 15592
rect 21692 15580 21698 15632
rect 22278 15620 22284 15632
rect 22239 15592 22284 15620
rect 22278 15580 22284 15592
rect 22336 15580 22342 15632
rect 22922 15620 22928 15632
rect 22883 15592 22928 15620
rect 22922 15580 22928 15592
rect 22980 15580 22986 15632
rect 24210 15580 24216 15632
rect 24268 15620 24274 15632
rect 24397 15623 24455 15629
rect 24397 15620 24409 15623
rect 24268 15592 24409 15620
rect 24268 15580 24274 15592
rect 24397 15589 24409 15592
rect 24443 15589 24455 15623
rect 24397 15583 24455 15589
rect 24578 15580 24584 15632
rect 24636 15620 24642 15632
rect 25866 15620 25872 15632
rect 24636 15592 25872 15620
rect 24636 15580 24642 15592
rect 25866 15580 25872 15592
rect 25924 15580 25930 15632
rect 26050 15580 26056 15632
rect 26108 15620 26114 15632
rect 26344 15620 26372 15648
rect 26108 15592 26372 15620
rect 26108 15580 26114 15592
rect 27430 15580 27436 15632
rect 27488 15620 27494 15632
rect 29656 15620 29684 15648
rect 27488 15592 29684 15620
rect 27488 15580 27494 15592
rect 19150 15552 19156 15564
rect 17972 15524 19156 15552
rect 17865 15515 17923 15521
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 19610 15552 19616 15564
rect 19571 15524 19616 15552
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 20162 15512 20168 15564
rect 20220 15552 20226 15564
rect 20714 15552 20720 15564
rect 20220 15524 20720 15552
rect 20220 15512 20226 15524
rect 1762 15484 1768 15496
rect 1723 15456 1768 15484
rect 1762 15444 1768 15456
rect 1820 15444 1826 15496
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15484 2743 15487
rect 3234 15484 3240 15496
rect 2731 15456 3240 15484
rect 2731 15453 2743 15456
rect 2685 15447 2743 15453
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15453 4399 15487
rect 4341 15447 4399 15453
rect 1489 15419 1547 15425
rect 1489 15385 1501 15419
rect 1535 15416 1547 15419
rect 3326 15416 3332 15428
rect 1535 15388 3332 15416
rect 1535 15385 1547 15388
rect 1489 15379 1547 15385
rect 3326 15376 3332 15388
rect 3384 15376 3390 15428
rect 4356 15416 4384 15447
rect 4522 15444 4528 15496
rect 4580 15484 4586 15496
rect 5077 15487 5135 15493
rect 5077 15484 5089 15487
rect 4580 15456 5089 15484
rect 4580 15444 4586 15456
rect 5077 15453 5089 15456
rect 5123 15453 5135 15487
rect 6638 15484 6644 15496
rect 5077 15447 5135 15453
rect 5276 15456 6644 15484
rect 5276 15416 5304 15456
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 6822 15444 6828 15496
rect 6880 15484 6886 15496
rect 7190 15493 7196 15496
rect 6917 15487 6975 15493
rect 6917 15484 6929 15487
rect 6880 15456 6929 15484
rect 6880 15444 6886 15456
rect 6917 15453 6929 15456
rect 6963 15453 6975 15487
rect 6917 15447 6975 15453
rect 7184 15447 7196 15493
rect 7248 15484 7254 15496
rect 7248 15456 7284 15484
rect 7190 15444 7196 15447
rect 7248 15444 7254 15456
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11517 15487 11575 15493
rect 11517 15484 11529 15487
rect 11204 15456 11529 15484
rect 11204 15444 11210 15456
rect 11517 15453 11529 15456
rect 11563 15453 11575 15487
rect 11517 15447 11575 15453
rect 12342 15444 12348 15496
rect 12400 15484 12406 15496
rect 13814 15484 13820 15496
rect 12400 15456 13820 15484
rect 12400 15444 12406 15456
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 15565 15487 15623 15493
rect 15565 15484 15577 15487
rect 14792 15456 15577 15484
rect 14792 15444 14798 15456
rect 15565 15453 15577 15456
rect 15611 15484 15623 15487
rect 16025 15487 16083 15493
rect 16025 15484 16037 15487
rect 15611 15456 16037 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 16025 15453 16037 15456
rect 16071 15484 16083 15487
rect 16666 15484 16672 15496
rect 16071 15456 16672 15484
rect 16071 15453 16083 15456
rect 16025 15447 16083 15453
rect 16666 15444 16672 15456
rect 16724 15484 16730 15496
rect 17954 15484 17960 15496
rect 16724 15456 17960 15484
rect 16724 15444 16730 15456
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 18141 15487 18199 15493
rect 18141 15453 18153 15487
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15484 19487 15487
rect 19518 15484 19524 15496
rect 19475 15456 19524 15484
rect 19475 15453 19487 15456
rect 19429 15447 19487 15453
rect 4356 15388 5304 15416
rect 5344 15419 5402 15425
rect 5344 15385 5356 15419
rect 5390 15416 5402 15419
rect 6546 15416 6552 15428
rect 5390 15388 6552 15416
rect 5390 15385 5402 15388
rect 5344 15379 5402 15385
rect 6546 15376 6552 15388
rect 6604 15376 6610 15428
rect 11422 15376 11428 15428
rect 11480 15416 11486 15428
rect 15320 15419 15378 15425
rect 11480 15388 14320 15416
rect 11480 15376 11486 15388
rect 2130 15308 2136 15360
rect 2188 15348 2194 15360
rect 5626 15348 5632 15360
rect 2188 15320 5632 15348
rect 2188 15308 2194 15320
rect 5626 15308 5632 15320
rect 5684 15308 5690 15360
rect 6457 15351 6515 15357
rect 6457 15317 6469 15351
rect 6503 15348 6515 15351
rect 9950 15348 9956 15360
rect 6503 15320 9956 15348
rect 6503 15317 6515 15320
rect 6457 15311 6515 15317
rect 9950 15308 9956 15320
rect 10008 15308 10014 15360
rect 14292 15348 14320 15388
rect 15320 15385 15332 15419
rect 15366 15416 15378 15419
rect 15470 15416 15476 15428
rect 15366 15388 15476 15416
rect 15366 15385 15378 15388
rect 15320 15379 15378 15385
rect 15470 15376 15476 15388
rect 15528 15376 15534 15428
rect 15746 15376 15752 15428
rect 15804 15416 15810 15428
rect 16270 15419 16328 15425
rect 16270 15416 16282 15419
rect 15804 15388 16282 15416
rect 15804 15376 15810 15388
rect 16270 15385 16282 15388
rect 16316 15385 16328 15419
rect 18156 15416 18184 15447
rect 19518 15444 19524 15456
rect 19576 15444 19582 15496
rect 20070 15484 20076 15496
rect 19628 15456 20076 15484
rect 19628 15416 19656 15456
rect 20070 15444 20076 15456
rect 20128 15444 20134 15496
rect 20364 15493 20392 15524
rect 20714 15512 20720 15524
rect 20772 15512 20778 15564
rect 21266 15552 21272 15564
rect 21227 15524 21272 15552
rect 21266 15512 21272 15524
rect 21324 15512 21330 15564
rect 22370 15512 22376 15564
rect 22428 15552 22434 15564
rect 22465 15555 22523 15561
rect 22465 15552 22477 15555
rect 22428 15524 22477 15552
rect 22428 15512 22434 15524
rect 22465 15521 22477 15524
rect 22511 15521 22523 15555
rect 26326 15552 26332 15564
rect 22465 15515 22523 15521
rect 22572 15524 23336 15552
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15453 20407 15487
rect 20349 15447 20407 15453
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15484 20499 15487
rect 21284 15484 21312 15512
rect 20487 15456 21312 15484
rect 21361 15487 21419 15493
rect 20487 15453 20499 15456
rect 20441 15447 20499 15453
rect 21361 15453 21373 15487
rect 21407 15484 21419 15487
rect 21542 15484 21548 15496
rect 21407 15456 21548 15484
rect 21407 15453 21419 15456
rect 21361 15447 21419 15453
rect 21542 15444 21548 15456
rect 21600 15444 21606 15496
rect 22572 15484 22600 15524
rect 22020 15456 22600 15484
rect 22020 15428 22048 15456
rect 22738 15444 22744 15496
rect 22796 15484 22802 15496
rect 23201 15487 23259 15493
rect 23201 15484 23213 15487
rect 22796 15456 23213 15484
rect 22796 15444 22802 15456
rect 23201 15453 23213 15456
rect 23247 15453 23259 15487
rect 23308 15484 23336 15524
rect 23860 15524 26332 15552
rect 23860 15496 23888 15524
rect 26326 15512 26332 15524
rect 26384 15512 26390 15564
rect 26418 15512 26424 15564
rect 26476 15552 26482 15564
rect 27893 15555 27951 15561
rect 27893 15552 27905 15555
rect 26476 15524 27905 15552
rect 26476 15512 26482 15524
rect 27893 15521 27905 15524
rect 27939 15521 27951 15555
rect 27893 15515 27951 15521
rect 23842 15484 23848 15496
rect 23308 15456 23428 15484
rect 23803 15456 23848 15484
rect 23201 15447 23259 15453
rect 16270 15379 16328 15385
rect 16408 15388 18184 15416
rect 18248 15388 19656 15416
rect 19705 15419 19763 15425
rect 16408 15348 16436 15388
rect 14292 15320 16436 15348
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 17218 15348 17224 15360
rect 16632 15320 17224 15348
rect 16632 15308 16638 15320
rect 17218 15308 17224 15320
rect 17276 15308 17282 15360
rect 17402 15348 17408 15360
rect 17363 15320 17408 15348
rect 17402 15308 17408 15320
rect 17460 15308 17466 15360
rect 17862 15308 17868 15360
rect 17920 15348 17926 15360
rect 18248 15348 18276 15388
rect 19705 15385 19717 15419
rect 19751 15416 19763 15419
rect 19978 15416 19984 15428
rect 19751 15388 19984 15416
rect 19751 15385 19763 15388
rect 19705 15379 19763 15385
rect 19978 15376 19984 15388
rect 20036 15376 20042 15428
rect 20622 15416 20628 15428
rect 20088 15388 20484 15416
rect 20535 15388 20628 15416
rect 17920 15320 18276 15348
rect 17920 15308 17926 15320
rect 18322 15308 18328 15360
rect 18380 15348 18386 15360
rect 20088 15348 20116 15388
rect 18380 15320 20116 15348
rect 18380 15308 18386 15320
rect 20162 15308 20168 15360
rect 20220 15348 20226 15360
rect 20456 15348 20484 15388
rect 20622 15376 20628 15388
rect 20680 15416 20686 15428
rect 21085 15419 21143 15425
rect 21085 15416 21097 15419
rect 20680 15388 21097 15416
rect 20680 15376 20686 15388
rect 21085 15385 21097 15388
rect 21131 15416 21143 15419
rect 21266 15416 21272 15428
rect 21131 15388 21272 15416
rect 21131 15385 21143 15388
rect 21085 15379 21143 15385
rect 21266 15376 21272 15388
rect 21324 15376 21330 15428
rect 22002 15416 22008 15428
rect 21963 15388 22008 15416
rect 22002 15376 22008 15388
rect 22060 15376 22066 15428
rect 22925 15419 22983 15425
rect 22925 15416 22937 15419
rect 22112 15388 22937 15416
rect 22112 15348 22140 15388
rect 22925 15385 22937 15388
rect 22971 15385 22983 15419
rect 22925 15379 22983 15385
rect 23109 15419 23167 15425
rect 23109 15385 23121 15419
rect 23155 15416 23167 15419
rect 23290 15416 23296 15428
rect 23155 15388 23296 15416
rect 23155 15385 23167 15388
rect 23109 15379 23167 15385
rect 23290 15376 23296 15388
rect 23348 15376 23354 15428
rect 20220 15320 20265 15348
rect 20456 15320 22140 15348
rect 23400 15348 23428 15456
rect 23842 15444 23848 15456
rect 23900 15444 23906 15496
rect 24394 15444 24400 15496
rect 24452 15484 24458 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 24452 15456 24593 15484
rect 24452 15444 24458 15456
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 24581 15447 24639 15453
rect 25225 15487 25283 15493
rect 25225 15453 25237 15487
rect 25271 15484 25283 15487
rect 29362 15484 29368 15496
rect 25271 15456 29368 15484
rect 25271 15453 25283 15456
rect 25225 15447 25283 15453
rect 24596 15416 24624 15447
rect 29362 15444 29368 15456
rect 29420 15444 29426 15496
rect 25682 15416 25688 15428
rect 24596 15388 25688 15416
rect 25682 15376 25688 15388
rect 25740 15376 25746 15428
rect 25041 15351 25099 15357
rect 25041 15348 25053 15351
rect 23400 15320 25053 15348
rect 20220 15308 20226 15320
rect 25041 15317 25053 15320
rect 25087 15348 25099 15351
rect 27430 15348 27436 15360
rect 25087 15320 27436 15348
rect 25087 15317 25099 15320
rect 25041 15311 25099 15317
rect 27430 15308 27436 15320
rect 27488 15308 27494 15360
rect 27522 15308 27528 15360
rect 27580 15348 27586 15360
rect 28445 15351 28503 15357
rect 28445 15348 28457 15351
rect 27580 15320 28457 15348
rect 27580 15308 27586 15320
rect 28445 15317 28457 15320
rect 28491 15348 28503 15351
rect 28626 15348 28632 15360
rect 28491 15320 28632 15348
rect 28491 15317 28503 15320
rect 28445 15311 28503 15317
rect 28626 15308 28632 15320
rect 28684 15308 28690 15360
rect 1104 15258 44896 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 44896 15258
rect 1104 15184 44896 15206
rect 8478 15144 8484 15156
rect 3436 15116 8484 15144
rect 2130 14968 2136 15020
rect 2188 15008 2194 15020
rect 3436 15017 3464 15116
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 8846 15104 8852 15156
rect 8904 15144 8910 15156
rect 11238 15144 11244 15156
rect 8904 15116 11244 15144
rect 8904 15104 8910 15116
rect 11238 15104 11244 15116
rect 11296 15144 11302 15156
rect 13354 15144 13360 15156
rect 11296 15116 13360 15144
rect 11296 15104 11302 15116
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 18598 15144 18604 15156
rect 15344 15116 18604 15144
rect 15344 15104 15350 15116
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 20165 15147 20223 15153
rect 18748 15116 20024 15144
rect 18748 15104 18754 15116
rect 8202 15076 8208 15088
rect 6288 15048 8208 15076
rect 3145 15011 3203 15017
rect 3145 15008 3157 15011
rect 2188 14980 3157 15008
rect 2188 14968 2194 14980
rect 3145 14977 3157 14980
rect 3191 14977 3203 15011
rect 3145 14971 3203 14977
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 4433 15011 4491 15017
rect 4433 14977 4445 15011
rect 4479 15008 4491 15011
rect 4522 15008 4528 15020
rect 4479 14980 4528 15008
rect 4479 14977 4491 14980
rect 4433 14971 4491 14977
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 4700 15011 4758 15017
rect 4700 14977 4712 15011
rect 4746 15008 4758 15011
rect 6288 15008 6316 15048
rect 8202 15036 8208 15048
rect 8260 15036 8266 15088
rect 12250 15076 12256 15088
rect 8312 15048 12256 15076
rect 4746 14980 6316 15008
rect 6365 15011 6423 15017
rect 4746 14977 4758 14980
rect 4700 14971 4758 14977
rect 6365 14977 6377 15011
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 15008 7067 15011
rect 7098 15008 7104 15020
rect 7055 14980 7104 15008
rect 7055 14977 7067 14980
rect 7009 14971 7067 14977
rect 2406 14940 2412 14952
rect 2367 14912 2412 14940
rect 2406 14900 2412 14912
rect 2464 14900 2470 14952
rect 2685 14943 2743 14949
rect 2685 14909 2697 14943
rect 2731 14909 2743 14943
rect 2685 14903 2743 14909
rect 750 14832 756 14884
rect 808 14872 814 14884
rect 2700 14872 2728 14903
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 6380 14940 6408 14971
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 7276 15011 7334 15017
rect 7276 14977 7288 15011
rect 7322 15008 7334 15011
rect 7558 15008 7564 15020
rect 7322 14980 7564 15008
rect 7322 14977 7334 14980
rect 7276 14971 7334 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 7742 14968 7748 15020
rect 7800 15008 7806 15020
rect 8312 15008 8340 15048
rect 12250 15036 12256 15048
rect 12308 15036 12314 15088
rect 12744 15079 12802 15085
rect 12744 15045 12756 15079
rect 12790 15076 12802 15079
rect 12894 15076 12900 15088
rect 12790 15048 12900 15076
rect 12790 15045 12802 15048
rect 12744 15039 12802 15045
rect 12894 15036 12900 15048
rect 12952 15036 12958 15088
rect 15010 15036 15016 15088
rect 15068 15076 15074 15088
rect 16936 15079 16994 15085
rect 15068 15048 16896 15076
rect 15068 15036 15074 15048
rect 12986 15008 12992 15020
rect 7800 14980 8340 15008
rect 12947 14980 12992 15008
rect 7800 14968 7806 14980
rect 12986 14968 12992 14980
rect 13044 14968 13050 15020
rect 14084 15011 14142 15017
rect 14084 14977 14096 15011
rect 14130 15008 14142 15011
rect 14550 15008 14556 15020
rect 14130 14980 14556 15008
rect 14130 14977 14142 14980
rect 14084 14971 14142 14977
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 15838 15008 15844 15020
rect 15799 14980 15844 15008
rect 15838 14968 15844 14980
rect 15896 14968 15902 15020
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 14977 15991 15011
rect 16666 15008 16672 15020
rect 16627 14980 16672 15008
rect 15933 14971 15991 14977
rect 8938 14940 8944 14952
rect 5684 14912 6408 14940
rect 8899 14912 8944 14940
rect 5684 14900 5690 14912
rect 8938 14900 8944 14912
rect 8996 14900 9002 14952
rect 10597 14943 10655 14949
rect 10597 14909 10609 14943
rect 10643 14909 10655 14943
rect 10597 14903 10655 14909
rect 10781 14943 10839 14949
rect 10781 14909 10793 14943
rect 10827 14940 10839 14943
rect 13817 14943 13875 14949
rect 10827 14912 11652 14940
rect 10827 14909 10839 14912
rect 10781 14903 10839 14909
rect 808 14844 2728 14872
rect 808 14832 814 14844
rect 8018 14832 8024 14884
rect 8076 14872 8082 14884
rect 10612 14872 10640 14903
rect 11624 14884 11652 14912
rect 13817 14909 13829 14943
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 11606 14872 11612 14884
rect 8076 14844 10640 14872
rect 11567 14844 11612 14872
rect 8076 14832 8082 14844
rect 11606 14832 11612 14844
rect 11664 14832 11670 14884
rect 5810 14804 5816 14816
rect 5771 14776 5816 14804
rect 5810 14764 5816 14776
rect 5868 14764 5874 14816
rect 5902 14764 5908 14816
rect 5960 14804 5966 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 5960 14776 6561 14804
rect 5960 14764 5966 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6549 14767 6607 14773
rect 6730 14764 6736 14816
rect 6788 14804 6794 14816
rect 7650 14804 7656 14816
rect 6788 14776 7656 14804
rect 6788 14764 6794 14776
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 8389 14807 8447 14813
rect 8389 14773 8401 14807
rect 8435 14804 8447 14807
rect 9490 14804 9496 14816
rect 8435 14776 9496 14804
rect 8435 14773 8447 14776
rect 8389 14767 8447 14773
rect 9490 14764 9496 14776
rect 9548 14764 9554 14816
rect 13832 14804 13860 14903
rect 15562 14900 15568 14952
rect 15620 14940 15626 14952
rect 15948 14940 15976 14971
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 16868 15008 16896 15048
rect 16936 15045 16948 15079
rect 16982 15076 16994 15079
rect 19797 15079 19855 15085
rect 16982 15048 19755 15076
rect 16982 15045 16994 15048
rect 16936 15039 16994 15045
rect 16868 14980 18000 15008
rect 16574 14940 16580 14952
rect 15620 14912 16580 14940
rect 15620 14900 15626 14912
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 17972 14940 18000 14980
rect 18046 14968 18052 15020
rect 18104 15008 18110 15020
rect 18509 15011 18567 15017
rect 18509 15008 18521 15011
rect 18104 14980 18521 15008
rect 18104 14968 18110 14980
rect 18509 14977 18521 14980
rect 18555 15008 18567 15011
rect 18874 15008 18880 15020
rect 18555 14980 18880 15008
rect 18555 14977 18567 14980
rect 18509 14971 18567 14977
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 19610 14940 19616 14952
rect 17972 14912 19616 14940
rect 19610 14900 19616 14912
rect 19668 14900 19674 14952
rect 19727 14940 19755 15048
rect 19797 15045 19809 15079
rect 19843 15076 19855 15079
rect 19886 15076 19892 15088
rect 19843 15048 19892 15076
rect 19843 15045 19855 15048
rect 19797 15039 19855 15045
rect 19886 15036 19892 15048
rect 19944 15036 19950 15088
rect 19996 15020 20024 15116
rect 20165 15113 20177 15147
rect 20211 15144 20223 15147
rect 20530 15144 20536 15156
rect 20211 15116 20536 15144
rect 20211 15113 20223 15116
rect 20165 15107 20223 15113
rect 20530 15104 20536 15116
rect 20588 15144 20594 15156
rect 20806 15144 20812 15156
rect 20588 15116 20812 15144
rect 20588 15104 20594 15116
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 21174 15144 21180 15156
rect 21135 15116 21180 15144
rect 21174 15104 21180 15116
rect 21232 15144 21238 15156
rect 21232 15116 22324 15144
rect 21232 15104 21238 15116
rect 21821 15079 21879 15085
rect 21821 15076 21833 15079
rect 20364 15048 21833 15076
rect 19978 15008 19984 15020
rect 19939 14980 19984 15008
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20073 15011 20131 15017
rect 20073 14977 20085 15011
rect 20119 15008 20131 15011
rect 20162 15008 20168 15020
rect 20119 14980 20168 15008
rect 20119 14977 20131 14980
rect 20073 14971 20131 14977
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 20364 15008 20392 15048
rect 21821 15045 21833 15048
rect 21867 15045 21879 15079
rect 22296 15076 22324 15116
rect 22370 15104 22376 15156
rect 22428 15144 22434 15156
rect 24670 15144 24676 15156
rect 22428 15116 24676 15144
rect 22428 15104 22434 15116
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 25590 15104 25596 15156
rect 25648 15144 25654 15156
rect 25685 15147 25743 15153
rect 25685 15144 25697 15147
rect 25648 15116 25697 15144
rect 25648 15104 25654 15116
rect 25685 15113 25697 15116
rect 25731 15113 25743 15147
rect 26326 15144 26332 15156
rect 26287 15116 26332 15144
rect 25685 15107 25743 15113
rect 26326 15104 26332 15116
rect 26384 15104 26390 15156
rect 26418 15104 26424 15156
rect 26476 15144 26482 15156
rect 26973 15147 27031 15153
rect 26973 15144 26985 15147
rect 26476 15116 26985 15144
rect 26476 15104 26482 15116
rect 26973 15113 26985 15116
rect 27019 15113 27031 15147
rect 26973 15107 27031 15113
rect 28258 15104 28264 15156
rect 28316 15144 28322 15156
rect 28442 15144 28448 15156
rect 28316 15116 28448 15144
rect 28316 15104 28322 15116
rect 28442 15104 28448 15116
rect 28500 15144 28506 15156
rect 30377 15147 30435 15153
rect 30377 15144 30389 15147
rect 28500 15116 30389 15144
rect 28500 15104 28506 15116
rect 30377 15113 30389 15116
rect 30423 15113 30435 15147
rect 30377 15107 30435 15113
rect 23198 15076 23204 15088
rect 22296 15048 23204 15076
rect 21821 15039 21879 15045
rect 23198 15036 23204 15048
rect 23256 15036 23262 15088
rect 25225 15079 25283 15085
rect 25225 15045 25237 15079
rect 25271 15076 25283 15079
rect 25498 15076 25504 15088
rect 25271 15048 25504 15076
rect 25271 15045 25283 15048
rect 25225 15039 25283 15045
rect 25498 15036 25504 15048
rect 25556 15036 25562 15088
rect 27246 15036 27252 15088
rect 27304 15076 27310 15088
rect 29733 15079 29791 15085
rect 29733 15076 29745 15079
rect 27304 15048 29745 15076
rect 27304 15036 27310 15048
rect 29733 15045 29745 15048
rect 29779 15045 29791 15079
rect 29733 15039 29791 15045
rect 20990 15008 20996 15020
rect 20272 14980 20392 15008
rect 20951 14980 20996 15008
rect 20272 14940 20300 14980
rect 20990 14968 20996 14980
rect 21048 14968 21054 15020
rect 21266 15008 21272 15020
rect 21179 14980 21272 15008
rect 21266 14968 21272 14980
rect 21324 15008 21330 15020
rect 21324 14980 21404 15008
rect 21324 14968 21330 14980
rect 19727 14912 20300 14940
rect 20349 14943 20407 14949
rect 20349 14909 20361 14943
rect 20395 14940 20407 14943
rect 20806 14940 20812 14952
rect 20395 14912 20812 14940
rect 20395 14909 20407 14912
rect 20349 14903 20407 14909
rect 18049 14875 18107 14881
rect 18049 14841 18061 14875
rect 18095 14872 18107 14875
rect 18966 14872 18972 14884
rect 18095 14844 18972 14872
rect 18095 14841 18107 14844
rect 18049 14835 18107 14841
rect 18966 14832 18972 14844
rect 19024 14832 19030 14884
rect 19426 14832 19432 14884
rect 19484 14872 19490 14884
rect 20364 14872 20392 14903
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 21376 14940 21404 14980
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21968 14980 22017 15008
rect 21968 14968 21974 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22186 14968 22192 15020
rect 22244 15008 22250 15020
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 22244 14980 22293 15008
rect 22244 14968 22250 14980
rect 22281 14977 22293 14980
rect 22327 14977 22339 15011
rect 22281 14971 22339 14977
rect 22738 14968 22744 15020
rect 22796 15008 22802 15020
rect 23385 15011 23443 15017
rect 23385 15008 23397 15011
rect 22796 14980 23397 15008
rect 22796 14968 22802 14980
rect 23385 14977 23397 14980
rect 23431 14977 23443 15011
rect 23385 14971 23443 14977
rect 25038 14968 25044 15020
rect 25096 15008 25102 15020
rect 25869 15011 25927 15017
rect 25869 15008 25881 15011
rect 25096 14980 25881 15008
rect 25096 14968 25102 14980
rect 25869 14977 25881 14980
rect 25915 14977 25927 15011
rect 25869 14971 25927 14977
rect 26418 14968 26424 15020
rect 26476 15008 26482 15020
rect 26694 15008 26700 15020
rect 26476 14980 26700 15008
rect 26476 14968 26482 14980
rect 26694 14968 26700 14980
rect 26752 14968 26758 15020
rect 27617 15011 27675 15017
rect 27617 14977 27629 15011
rect 27663 15008 27675 15011
rect 27706 15008 27712 15020
rect 27663 14980 27712 15008
rect 27663 14977 27675 14980
rect 27617 14971 27675 14977
rect 27706 14968 27712 14980
rect 27764 15008 27770 15020
rect 28442 15008 28448 15020
rect 27764 14980 28448 15008
rect 27764 14968 27770 14980
rect 28442 14968 28448 14980
rect 28500 15008 28506 15020
rect 28810 15008 28816 15020
rect 28500 14980 28816 15008
rect 28500 14968 28506 14980
rect 28810 14968 28816 14980
rect 28868 14968 28874 15020
rect 22830 14940 22836 14952
rect 21376 14912 22836 14940
rect 22830 14900 22836 14912
rect 22888 14900 22894 14952
rect 23290 14940 23296 14952
rect 23124 14912 23296 14940
rect 19484 14844 20392 14872
rect 19484 14832 19490 14844
rect 20438 14832 20444 14884
rect 20496 14872 20502 14884
rect 21358 14872 21364 14884
rect 20496 14844 21364 14872
rect 20496 14832 20502 14844
rect 21358 14832 21364 14844
rect 21416 14872 21422 14884
rect 23124 14881 23152 14912
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 23566 14900 23572 14952
rect 23624 14940 23630 14952
rect 24305 14943 24363 14949
rect 24305 14940 24317 14943
rect 23624 14912 24317 14940
rect 23624 14900 23630 14912
rect 24305 14909 24317 14912
rect 24351 14940 24363 14943
rect 24394 14940 24400 14952
rect 24351 14912 24400 14940
rect 24351 14909 24363 14912
rect 24305 14903 24363 14909
rect 24394 14900 24400 14912
rect 24452 14940 24458 14952
rect 28077 14943 28135 14949
rect 28077 14940 28089 14943
rect 24452 14912 28089 14940
rect 24452 14900 24458 14912
rect 28077 14909 28089 14912
rect 28123 14909 28135 14943
rect 28077 14903 28135 14909
rect 22189 14875 22247 14881
rect 22189 14872 22201 14875
rect 21416 14844 22201 14872
rect 21416 14832 21422 14844
rect 22189 14841 22201 14844
rect 22235 14841 22247 14875
rect 22189 14835 22247 14841
rect 23109 14875 23167 14881
rect 23109 14841 23121 14875
rect 23155 14841 23167 14875
rect 24026 14872 24032 14884
rect 23987 14844 24032 14872
rect 23109 14835 23167 14841
rect 24026 14832 24032 14844
rect 24084 14872 24090 14884
rect 24670 14872 24676 14884
rect 24084 14844 24676 14872
rect 24084 14832 24090 14844
rect 24670 14832 24676 14844
rect 24728 14832 24734 14884
rect 24857 14875 24915 14881
rect 24857 14841 24869 14875
rect 24903 14841 24915 14875
rect 24857 14835 24915 14841
rect 14090 14804 14096 14816
rect 13832 14776 14096 14804
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 15102 14764 15108 14816
rect 15160 14804 15166 14816
rect 15197 14807 15255 14813
rect 15197 14804 15209 14807
rect 15160 14776 15209 14804
rect 15160 14764 15166 14776
rect 15197 14773 15209 14776
rect 15243 14773 15255 14807
rect 15197 14767 15255 14773
rect 16117 14807 16175 14813
rect 16117 14773 16129 14807
rect 16163 14804 16175 14807
rect 16574 14804 16580 14816
rect 16163 14776 16580 14804
rect 16163 14773 16175 14776
rect 16117 14767 16175 14773
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 18739 14807 18797 14813
rect 18739 14804 18751 14807
rect 18472 14776 18751 14804
rect 18472 14764 18478 14776
rect 18739 14773 18751 14776
rect 18785 14773 18797 14807
rect 18739 14767 18797 14773
rect 19702 14764 19708 14816
rect 19760 14804 19766 14816
rect 20809 14807 20867 14813
rect 20809 14804 20821 14807
rect 19760 14776 20821 14804
rect 19760 14764 19766 14776
rect 20809 14773 20821 14776
rect 20855 14773 20867 14807
rect 20809 14767 20867 14773
rect 20990 14764 20996 14816
rect 21048 14804 21054 14816
rect 22830 14804 22836 14816
rect 21048 14776 22836 14804
rect 21048 14764 21054 14776
rect 22830 14764 22836 14776
rect 22888 14764 22894 14816
rect 22925 14807 22983 14813
rect 22925 14773 22937 14807
rect 22971 14804 22983 14807
rect 23290 14804 23296 14816
rect 22971 14776 23296 14804
rect 22971 14773 22983 14776
rect 22925 14767 22983 14773
rect 23290 14764 23296 14776
rect 23348 14764 23354 14816
rect 23842 14804 23848 14816
rect 23803 14776 23848 14804
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 24578 14764 24584 14816
rect 24636 14804 24642 14816
rect 24765 14807 24823 14813
rect 24765 14804 24777 14807
rect 24636 14776 24777 14804
rect 24636 14764 24642 14776
rect 24765 14773 24777 14776
rect 24811 14773 24823 14807
rect 24872 14804 24900 14835
rect 24946 14832 24952 14884
rect 25004 14872 25010 14884
rect 29181 14875 29239 14881
rect 29181 14872 29193 14875
rect 25004 14844 29193 14872
rect 25004 14832 25010 14844
rect 29181 14841 29193 14844
rect 29227 14841 29239 14875
rect 29181 14835 29239 14841
rect 27430 14804 27436 14816
rect 24872 14776 27436 14804
rect 24765 14767 24823 14773
rect 27430 14764 27436 14776
rect 27488 14764 27494 14816
rect 27798 14764 27804 14816
rect 27856 14804 27862 14816
rect 28258 14804 28264 14816
rect 27856 14776 28264 14804
rect 27856 14764 27862 14776
rect 28258 14764 28264 14776
rect 28316 14764 28322 14816
rect 28626 14804 28632 14816
rect 28587 14776 28632 14804
rect 28626 14764 28632 14776
rect 28684 14764 28690 14816
rect 1104 14714 44896 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 44896 14714
rect 1104 14640 44896 14662
rect 934 14560 940 14612
rect 992 14600 998 14612
rect 1489 14603 1547 14609
rect 1489 14600 1501 14603
rect 992 14572 1501 14600
rect 992 14560 998 14572
rect 1489 14569 1501 14572
rect 1535 14569 1547 14603
rect 1489 14563 1547 14569
rect 1949 14603 2007 14609
rect 1949 14569 1961 14603
rect 1995 14600 2007 14603
rect 3970 14600 3976 14612
rect 1995 14572 3976 14600
rect 1995 14569 2007 14572
rect 1949 14563 2007 14569
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 8938 14600 8944 14612
rect 4120 14572 8944 14600
rect 4120 14560 4126 14572
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 12986 14600 12992 14612
rect 9916 14572 12992 14600
rect 9916 14560 9922 14572
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 13170 14600 13176 14612
rect 13131 14572 13176 14600
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 13320 14572 19012 14600
rect 13320 14560 13326 14572
rect 3007 14535 3065 14541
rect 3007 14501 3019 14535
rect 3053 14532 3065 14535
rect 4338 14532 4344 14544
rect 3053 14504 4344 14532
rect 3053 14501 3065 14504
rect 3007 14495 3065 14501
rect 4338 14492 4344 14504
rect 4396 14492 4402 14544
rect 4798 14532 4804 14544
rect 4448 14504 4804 14532
rect 1857 14467 1915 14473
rect 1857 14433 1869 14467
rect 1903 14464 1915 14467
rect 3786 14464 3792 14476
rect 1903 14436 3792 14464
rect 1903 14433 1915 14436
rect 1857 14427 1915 14433
rect 3786 14424 3792 14436
rect 3844 14424 3850 14476
rect 4448 14473 4476 14504
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 6270 14492 6276 14544
rect 6328 14532 6334 14544
rect 6549 14535 6607 14541
rect 6549 14532 6561 14535
rect 6328 14504 6561 14532
rect 6328 14492 6334 14504
rect 6549 14501 6561 14504
rect 6595 14501 6607 14535
rect 6549 14495 6607 14501
rect 8294 14492 8300 14544
rect 8352 14532 8358 14544
rect 11146 14532 11152 14544
rect 8352 14504 11152 14532
rect 8352 14492 8358 14504
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 12618 14532 12624 14544
rect 12579 14504 12624 14532
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 12710 14492 12716 14544
rect 12768 14532 12774 14544
rect 15473 14535 15531 14541
rect 12768 14504 14136 14532
rect 12768 14492 12774 14504
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14433 4491 14467
rect 4706 14464 4712 14476
rect 4667 14436 4712 14464
rect 4433 14427 4491 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 7009 14467 7067 14473
rect 7009 14464 7021 14467
rect 6880 14436 7021 14464
rect 6880 14424 6886 14436
rect 7009 14433 7021 14436
rect 7055 14433 7067 14467
rect 14108 14464 14136 14504
rect 15473 14501 15485 14535
rect 15519 14532 15531 14535
rect 15654 14532 15660 14544
rect 15519 14504 15660 14532
rect 15519 14501 15531 14504
rect 15473 14495 15531 14501
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 17402 14532 17408 14544
rect 17363 14504 17408 14532
rect 17402 14492 17408 14504
rect 17460 14492 17466 14544
rect 18417 14467 18475 14473
rect 14108 14436 14228 14464
rect 7009 14427 7067 14433
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 3234 14396 3240 14408
rect 3195 14368 3240 14396
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3602 14356 3608 14408
rect 3660 14396 3666 14408
rect 3660 14368 4568 14396
rect 3660 14356 3666 14368
rect 1949 14331 2007 14337
rect 1949 14297 1961 14331
rect 1995 14328 2007 14331
rect 3694 14328 3700 14340
rect 1995 14300 3700 14328
rect 1995 14297 2007 14300
rect 1949 14291 2007 14297
rect 3694 14288 3700 14300
rect 3752 14288 3758 14340
rect 4540 14328 4568 14368
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 4672 14368 5181 14396
rect 4672 14356 4678 14368
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5433 14396 5439 14408
rect 5394 14368 5439 14396
rect 5169 14359 5227 14365
rect 5433 14356 5439 14368
rect 5491 14356 5497 14408
rect 6270 14356 6276 14408
rect 6328 14396 6334 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 6328 14368 8953 14396
rect 6328 14356 6334 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 11238 14396 11244 14408
rect 10836 14368 10881 14396
rect 11199 14368 11244 14396
rect 10836 14356 10842 14368
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 11514 14405 11520 14408
rect 11508 14359 11520 14405
rect 11572 14396 11578 14408
rect 13906 14396 13912 14408
rect 11572 14368 11608 14396
rect 12406 14368 13912 14396
rect 11514 14356 11520 14359
rect 11572 14356 11578 14368
rect 6178 14328 6184 14340
rect 4540 14300 6184 14328
rect 6178 14288 6184 14300
rect 6236 14288 6242 14340
rect 6362 14288 6368 14340
rect 6420 14328 6426 14340
rect 7276 14331 7334 14337
rect 6420 14300 6684 14328
rect 6420 14288 6426 14300
rect 3234 14220 3240 14272
rect 3292 14260 3298 14272
rect 3878 14260 3884 14272
rect 3292 14232 3884 14260
rect 3292 14220 3298 14232
rect 3878 14220 3884 14232
rect 3936 14260 3942 14272
rect 6454 14260 6460 14272
rect 3936 14232 6460 14260
rect 3936 14220 3942 14232
rect 6454 14220 6460 14232
rect 6512 14220 6518 14272
rect 6656 14260 6684 14300
rect 7276 14297 7288 14331
rect 7322 14328 7334 14331
rect 7834 14328 7840 14340
rect 7322 14300 7840 14328
rect 7322 14297 7334 14300
rect 7276 14291 7334 14297
rect 7834 14288 7840 14300
rect 7892 14288 7898 14340
rect 7926 14288 7932 14340
rect 7984 14328 7990 14340
rect 8570 14328 8576 14340
rect 7984 14300 8576 14328
rect 7984 14288 7990 14300
rect 8570 14288 8576 14300
rect 8628 14288 8634 14340
rect 10042 14288 10048 14340
rect 10100 14328 10106 14340
rect 10597 14331 10655 14337
rect 10597 14328 10609 14331
rect 10100 14300 10609 14328
rect 10100 14288 10106 14300
rect 10597 14297 10609 14300
rect 10643 14297 10655 14331
rect 10597 14291 10655 14297
rect 11146 14288 11152 14340
rect 11204 14328 11210 14340
rect 11974 14328 11980 14340
rect 11204 14300 11980 14328
rect 11204 14288 11210 14300
rect 11974 14288 11980 14300
rect 12032 14288 12038 14340
rect 8018 14260 8024 14272
rect 6656 14232 8024 14260
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 8389 14263 8447 14269
rect 8389 14229 8401 14263
rect 8435 14260 8447 14263
rect 12406 14260 12434 14368
rect 13906 14356 13912 14368
rect 13964 14356 13970 14408
rect 14090 14396 14096 14408
rect 14051 14368 14096 14396
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 14200 14396 14228 14436
rect 18417 14433 18429 14467
rect 18463 14433 18475 14467
rect 18984 14464 19012 14572
rect 19610 14560 19616 14612
rect 19668 14600 19674 14612
rect 19889 14603 19947 14609
rect 19889 14600 19901 14603
rect 19668 14572 19901 14600
rect 19668 14560 19674 14572
rect 19889 14569 19901 14572
rect 19935 14569 19947 14603
rect 19889 14563 19947 14569
rect 19978 14560 19984 14612
rect 20036 14600 20042 14612
rect 20438 14600 20444 14612
rect 20036 14572 20444 14600
rect 20036 14560 20042 14572
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 21726 14560 21732 14612
rect 21784 14600 21790 14612
rect 22002 14600 22008 14612
rect 21784 14572 22008 14600
rect 21784 14560 21790 14572
rect 22002 14560 22008 14572
rect 22060 14600 22066 14612
rect 22373 14603 22431 14609
rect 22373 14600 22385 14603
rect 22060 14572 22385 14600
rect 22060 14560 22066 14572
rect 22373 14569 22385 14572
rect 22419 14600 22431 14603
rect 24397 14603 24455 14609
rect 24397 14600 24409 14603
rect 22419 14572 24409 14600
rect 22419 14569 22431 14572
rect 22373 14563 22431 14569
rect 24397 14569 24409 14572
rect 24443 14569 24455 14603
rect 24397 14563 24455 14569
rect 25777 14603 25835 14609
rect 25777 14569 25789 14603
rect 25823 14600 25835 14603
rect 26050 14600 26056 14612
rect 25823 14572 26056 14600
rect 25823 14569 25835 14572
rect 25777 14563 25835 14569
rect 26050 14560 26056 14572
rect 26108 14560 26114 14612
rect 26881 14603 26939 14609
rect 26881 14569 26893 14603
rect 26927 14600 26939 14603
rect 26970 14600 26976 14612
rect 26927 14572 26976 14600
rect 26927 14569 26939 14572
rect 26881 14563 26939 14569
rect 26970 14560 26976 14572
rect 27028 14560 27034 14612
rect 27430 14600 27436 14612
rect 27391 14572 27436 14600
rect 27430 14560 27436 14572
rect 27488 14560 27494 14612
rect 27614 14560 27620 14612
rect 27672 14600 27678 14612
rect 28445 14603 28503 14609
rect 28445 14600 28457 14603
rect 27672 14572 28457 14600
rect 27672 14560 27678 14572
rect 28445 14569 28457 14572
rect 28491 14569 28503 14603
rect 28445 14563 28503 14569
rect 29641 14603 29699 14609
rect 29641 14569 29653 14603
rect 29687 14600 29699 14603
rect 30006 14600 30012 14612
rect 29687 14572 30012 14600
rect 29687 14569 29699 14572
rect 29641 14563 29699 14569
rect 20070 14492 20076 14544
rect 20128 14532 20134 14544
rect 20128 14504 20300 14532
rect 20128 14492 20134 14504
rect 20272 14464 20300 14504
rect 20346 14492 20352 14544
rect 20404 14532 20410 14544
rect 20717 14535 20775 14541
rect 20404 14504 20449 14532
rect 20404 14492 20410 14504
rect 20717 14501 20729 14535
rect 20763 14532 20775 14535
rect 22186 14532 22192 14544
rect 20763 14504 22192 14532
rect 20763 14501 20775 14504
rect 20717 14495 20775 14501
rect 22186 14492 22192 14504
rect 22244 14492 22250 14544
rect 22830 14492 22836 14544
rect 22888 14532 22894 14544
rect 23017 14535 23075 14541
rect 23017 14532 23029 14535
rect 22888 14504 23029 14532
rect 22888 14492 22894 14504
rect 23017 14501 23029 14504
rect 23063 14501 23075 14535
rect 23382 14532 23388 14544
rect 23017 14495 23075 14501
rect 23124 14504 23388 14532
rect 21637 14467 21695 14473
rect 18984 14436 19196 14464
rect 20272 14436 21588 14464
rect 18417 14427 18475 14433
rect 15562 14396 15568 14408
rect 14200 14368 15568 14396
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14396 16083 14399
rect 16666 14396 16672 14408
rect 16071 14368 16672 14396
rect 16071 14365 16083 14368
rect 16025 14359 16083 14365
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 16758 14356 16764 14408
rect 16816 14396 16822 14408
rect 18432 14396 18460 14427
rect 18690 14396 18696 14408
rect 16816 14368 18460 14396
rect 18651 14368 18696 14396
rect 16816 14356 16822 14368
rect 18690 14356 18696 14368
rect 18748 14356 18754 14408
rect 19168 14392 19196 14436
rect 19242 14392 19248 14408
rect 19168 14364 19248 14392
rect 19300 14396 19306 14408
rect 19300 14368 19393 14396
rect 19242 14356 19248 14364
rect 19300 14356 19306 14368
rect 19426 14356 19432 14408
rect 19484 14405 19490 14408
rect 19484 14399 19533 14405
rect 19484 14365 19487 14399
rect 19521 14365 19533 14399
rect 19484 14359 19533 14365
rect 19484 14356 19490 14359
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 20533 14399 20591 14405
rect 19760 14368 19805 14396
rect 19760 14356 19766 14368
rect 20533 14365 20545 14399
rect 20579 14365 20591 14399
rect 20806 14396 20812 14408
rect 20767 14368 20812 14396
rect 20533 14359 20591 14365
rect 13354 14328 13360 14340
rect 13315 14300 13360 14328
rect 13354 14288 13360 14300
rect 13412 14288 13418 14340
rect 13538 14328 13544 14340
rect 13499 14300 13544 14328
rect 13538 14288 13544 14300
rect 13596 14288 13602 14340
rect 13998 14288 14004 14340
rect 14056 14328 14062 14340
rect 16298 14337 16304 14340
rect 14338 14331 14396 14337
rect 14338 14328 14350 14331
rect 14056 14300 14350 14328
rect 14056 14288 14062 14300
rect 14338 14297 14350 14300
rect 14384 14297 14396 14331
rect 14338 14291 14396 14297
rect 16292 14291 16304 14337
rect 16356 14328 16362 14340
rect 20548 14328 20576 14359
rect 20806 14356 20812 14368
rect 20864 14356 20870 14408
rect 21450 14396 21456 14408
rect 21411 14368 21456 14396
rect 21450 14356 21456 14368
rect 21508 14356 21514 14408
rect 21082 14328 21088 14340
rect 16356 14300 16392 14328
rect 16500 14300 20392 14328
rect 20548 14300 21088 14328
rect 16298 14288 16304 14291
rect 16356 14288 16362 14300
rect 8435 14232 12434 14260
rect 8435 14229 8447 14232
rect 8389 14223 8447 14229
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 16500 14260 16528 14300
rect 13688 14232 16528 14260
rect 13688 14220 13694 14232
rect 16574 14220 16580 14272
rect 16632 14260 16638 14272
rect 18414 14260 18420 14272
rect 16632 14232 18420 14260
rect 16632 14220 16638 14232
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 19242 14220 19248 14272
rect 19300 14260 19306 14272
rect 20162 14260 20168 14272
rect 19300 14232 20168 14260
rect 19300 14220 19306 14232
rect 20162 14220 20168 14232
rect 20220 14220 20226 14272
rect 20364 14260 20392 14300
rect 21082 14288 21088 14300
rect 21140 14288 21146 14340
rect 21266 14328 21272 14340
rect 21227 14300 21272 14328
rect 21266 14288 21272 14300
rect 21324 14288 21330 14340
rect 21560 14328 21588 14436
rect 21637 14433 21649 14467
rect 21683 14464 21695 14467
rect 22370 14464 22376 14476
rect 21683 14436 22376 14464
rect 21683 14433 21695 14436
rect 21637 14427 21695 14433
rect 22370 14424 22376 14436
rect 22428 14424 22434 14476
rect 23124 14464 23152 14504
rect 23382 14492 23388 14504
rect 23440 14532 23446 14544
rect 27062 14532 27068 14544
rect 23440 14504 27068 14532
rect 23440 14492 23446 14504
rect 27062 14492 27068 14504
rect 27120 14492 27126 14544
rect 22572 14436 23152 14464
rect 21726 14396 21732 14408
rect 21687 14368 21732 14396
rect 21726 14356 21732 14368
rect 21784 14356 21790 14408
rect 22462 14328 22468 14340
rect 21560 14300 22468 14328
rect 22462 14288 22468 14300
rect 22520 14288 22526 14340
rect 22572 14337 22600 14436
rect 23566 14424 23572 14476
rect 23624 14464 23630 14476
rect 25133 14467 25191 14473
rect 25133 14464 25145 14467
rect 23624 14436 25145 14464
rect 23624 14424 23630 14436
rect 25133 14433 25145 14436
rect 25179 14433 25191 14467
rect 25133 14427 25191 14433
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14396 23259 14399
rect 23385 14399 23443 14405
rect 23247 14368 23336 14396
rect 23247 14365 23259 14368
rect 23201 14359 23259 14365
rect 22557 14331 22615 14337
rect 22557 14297 22569 14331
rect 22603 14297 22615 14331
rect 22557 14291 22615 14297
rect 22094 14260 22100 14272
rect 20364 14232 22100 14260
rect 22094 14220 22100 14232
rect 22152 14260 22158 14272
rect 22347 14263 22405 14269
rect 22347 14260 22359 14263
rect 22152 14232 22359 14260
rect 22152 14220 22158 14232
rect 22347 14229 22359 14232
rect 22393 14229 22405 14263
rect 23308 14260 23336 14368
rect 23385 14365 23397 14399
rect 23431 14396 23443 14399
rect 24026 14396 24032 14408
rect 23431 14368 24032 14396
rect 23431 14365 23443 14368
rect 23385 14359 23443 14365
rect 24026 14356 24032 14368
rect 24084 14356 24090 14408
rect 24581 14399 24639 14405
rect 24581 14365 24593 14399
rect 24627 14396 24639 14399
rect 24670 14396 24676 14408
rect 24627 14368 24676 14396
rect 24627 14365 24639 14368
rect 24581 14359 24639 14365
rect 24670 14356 24676 14368
rect 24728 14356 24734 14408
rect 24854 14356 24860 14408
rect 24912 14396 24918 14408
rect 25041 14399 25099 14405
rect 25041 14396 25053 14399
rect 24912 14368 25053 14396
rect 24912 14356 24918 14368
rect 25041 14365 25053 14368
rect 25087 14365 25099 14399
rect 25041 14359 25099 14365
rect 25225 14399 25283 14405
rect 25225 14365 25237 14399
rect 25271 14396 25283 14399
rect 29656 14396 29684 14563
rect 30006 14560 30012 14572
rect 30064 14560 30070 14612
rect 25271 14368 29684 14396
rect 25271 14365 25283 14368
rect 25225 14359 25283 14365
rect 24044 14328 24072 14356
rect 24946 14328 24952 14340
rect 24044 14300 24952 14328
rect 24946 14288 24952 14300
rect 25004 14288 25010 14340
rect 26786 14328 26792 14340
rect 26160 14300 26792 14328
rect 26160 14260 26188 14300
rect 26786 14288 26792 14300
rect 26844 14328 26850 14340
rect 30101 14331 30159 14337
rect 30101 14328 30113 14331
rect 26844 14300 30113 14328
rect 26844 14288 26850 14300
rect 30101 14297 30113 14300
rect 30147 14297 30159 14331
rect 30101 14291 30159 14297
rect 26326 14260 26332 14272
rect 23308 14232 26188 14260
rect 26287 14232 26332 14260
rect 22347 14223 22405 14229
rect 26326 14220 26332 14232
rect 26384 14220 26390 14272
rect 27890 14260 27896 14272
rect 27851 14232 27896 14260
rect 27890 14220 27896 14232
rect 27948 14220 27954 14272
rect 30650 14260 30656 14272
rect 30611 14232 30656 14260
rect 30650 14220 30656 14232
rect 30708 14260 30714 14272
rect 33502 14260 33508 14272
rect 30708 14232 33508 14260
rect 30708 14220 30714 14232
rect 33502 14220 33508 14232
rect 33560 14220 33566 14272
rect 1104 14170 44896 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 44896 14170
rect 1104 14096 44896 14118
rect 382 14016 388 14068
rect 440 14056 446 14068
rect 2501 14059 2559 14065
rect 2501 14056 2513 14059
rect 440 14028 2513 14056
rect 440 14016 446 14028
rect 2501 14025 2513 14028
rect 2547 14025 2559 14059
rect 2501 14019 2559 14025
rect 2682 14016 2688 14068
rect 2740 14016 2746 14068
rect 5813 14059 5871 14065
rect 5813 14025 5825 14059
rect 5859 14056 5871 14059
rect 7466 14056 7472 14068
rect 5859 14028 7472 14056
rect 5859 14025 5871 14028
rect 5813 14019 5871 14025
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 7745 14059 7803 14065
rect 7745 14025 7757 14059
rect 7791 14056 7803 14059
rect 7926 14056 7932 14068
rect 7791 14028 7932 14056
rect 7791 14025 7803 14028
rect 7745 14019 7803 14025
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 8260 14028 11928 14056
rect 8260 14016 8266 14028
rect 2700 13988 2728 14016
rect 5626 13988 5632 14000
rect 1412 13960 2728 13988
rect 4356 13960 5632 13988
rect 1412 13929 1440 13960
rect 1397 13923 1455 13929
rect 1397 13889 1409 13923
rect 1443 13889 1455 13923
rect 1397 13883 1455 13889
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13889 2191 13923
rect 2314 13920 2320 13932
rect 2275 13892 2320 13920
rect 2133 13883 2191 13889
rect 2148 13852 2176 13883
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 3510 13920 3516 13932
rect 2731 13892 3516 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 3510 13880 3516 13892
rect 3568 13920 3574 13932
rect 4356 13920 4384 13960
rect 5626 13948 5632 13960
rect 5684 13948 5690 14000
rect 6454 13988 6460 14000
rect 6367 13960 6460 13988
rect 3568 13892 4384 13920
rect 4433 13923 4491 13929
rect 3568 13880 3574 13892
rect 4433 13889 4445 13923
rect 4479 13920 4491 13923
rect 4522 13920 4528 13932
rect 4479 13892 4528 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4700 13923 4758 13929
rect 4700 13889 4712 13923
rect 4746 13920 4758 13923
rect 4982 13920 4988 13932
rect 4746 13892 4988 13920
rect 4746 13889 4758 13892
rect 4700 13883 4758 13889
rect 4982 13880 4988 13892
rect 5040 13880 5046 13932
rect 5258 13880 5264 13932
rect 5316 13920 5322 13932
rect 6270 13920 6276 13932
rect 5316 13892 6276 13920
rect 5316 13880 5322 13892
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 6380 13929 6408 13960
rect 6454 13948 6460 13960
rect 6512 13988 6518 14000
rect 6822 13988 6828 14000
rect 6512 13960 6828 13988
rect 6512 13948 6518 13960
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 8389 13991 8447 13997
rect 8389 13988 8401 13991
rect 8076 13960 8401 13988
rect 8076 13948 8082 13960
rect 8389 13957 8401 13960
rect 8435 13957 8447 13991
rect 8389 13951 8447 13957
rect 9306 13948 9312 14000
rect 9364 13988 9370 14000
rect 9364 13960 9628 13988
rect 9364 13948 9370 13960
rect 6638 13929 6644 13932
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 6632 13883 6644 13929
rect 6696 13920 6702 13932
rect 8205 13923 8263 13929
rect 8205 13920 8217 13923
rect 6696 13892 6732 13920
rect 8128 13892 8217 13920
rect 6638 13880 6644 13883
rect 6696 13880 6702 13892
rect 2590 13852 2596 13864
rect 2148 13824 2596 13852
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 3602 13852 3608 13864
rect 2700 13824 3608 13852
rect 1578 13784 1584 13796
rect 1491 13756 1584 13784
rect 1578 13744 1584 13756
rect 1636 13784 1642 13796
rect 2700 13784 2728 13824
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13821 3755 13855
rect 3970 13852 3976 13864
rect 3931 13824 3976 13852
rect 3697 13815 3755 13821
rect 1636 13756 2728 13784
rect 1636 13744 1642 13756
rect 2222 13716 2228 13728
rect 2183 13688 2228 13716
rect 2222 13676 2228 13688
rect 2280 13716 2286 13728
rect 3234 13716 3240 13728
rect 2280 13688 3240 13716
rect 2280 13676 2286 13688
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 3712 13716 3740 13815
rect 3970 13812 3976 13824
rect 4028 13812 4034 13864
rect 7926 13744 7932 13796
rect 7984 13784 7990 13796
rect 8128 13784 8156 13892
rect 8205 13889 8217 13892
rect 8251 13889 8263 13923
rect 9600 13920 9628 13960
rect 10502 13948 10508 14000
rect 10560 13988 10566 14000
rect 10560 13960 10824 13988
rect 10560 13948 10566 13960
rect 10796 13929 10824 13960
rect 11054 13948 11060 14000
rect 11112 13988 11118 14000
rect 11762 13991 11820 13997
rect 11762 13988 11774 13991
rect 11112 13960 11774 13988
rect 11112 13948 11118 13960
rect 11762 13957 11774 13960
rect 11808 13957 11820 13991
rect 11762 13951 11820 13957
rect 10689 13923 10747 13929
rect 10689 13920 10701 13923
rect 9600 13892 10701 13920
rect 8205 13883 8263 13889
rect 10689 13889 10701 13892
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13889 11023 13923
rect 11900 13920 11928 14028
rect 12250 14016 12256 14068
rect 12308 14056 12314 14068
rect 18046 14056 18052 14068
rect 12308 14028 18052 14056
rect 12308 14016 12314 14028
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 19242 14056 19248 14068
rect 18432 14028 19248 14056
rect 11974 13948 11980 14000
rect 12032 13988 12038 14000
rect 13817 13991 13875 13997
rect 13817 13988 13829 13991
rect 12032 13960 13829 13988
rect 12032 13948 12038 13960
rect 13817 13957 13829 13960
rect 13863 13957 13875 13991
rect 13817 13951 13875 13957
rect 14090 13948 14096 14000
rect 14148 13988 14154 14000
rect 16936 13991 16994 13997
rect 14148 13960 16712 13988
rect 14148 13948 14154 13960
rect 14458 13920 14464 13932
rect 11900 13892 12940 13920
rect 10965 13883 11023 13889
rect 8570 13812 8576 13864
rect 8628 13852 8634 13864
rect 9858 13852 9864 13864
rect 8628 13824 9864 13852
rect 8628 13812 8634 13824
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 7984 13756 9260 13784
rect 7984 13744 7990 13756
rect 9122 13716 9128 13728
rect 3712 13688 9128 13716
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9232 13716 9260 13756
rect 9674 13744 9680 13796
rect 9732 13784 9738 13796
rect 10060 13784 10088 13815
rect 10410 13812 10416 13864
rect 10468 13852 10474 13864
rect 10468 13824 10548 13852
rect 10468 13812 10474 13824
rect 10520 13793 10548 13824
rect 10594 13812 10600 13864
rect 10652 13852 10658 13864
rect 10980 13852 11008 13883
rect 10652 13824 11008 13852
rect 10652 13812 10658 13824
rect 11238 13812 11244 13864
rect 11296 13852 11302 13864
rect 11517 13855 11575 13861
rect 11517 13852 11529 13855
rect 11296 13824 11529 13852
rect 11296 13812 11302 13824
rect 11517 13821 11529 13824
rect 11563 13821 11575 13855
rect 11517 13815 11575 13821
rect 12912 13852 12940 13892
rect 13924 13892 14464 13920
rect 13814 13852 13820 13864
rect 12912 13824 13820 13852
rect 9732 13756 10088 13784
rect 10505 13787 10563 13793
rect 9732 13744 9738 13756
rect 10505 13753 10517 13787
rect 10551 13753 10563 13787
rect 11146 13784 11152 13796
rect 10505 13747 10563 13753
rect 10612 13756 11152 13784
rect 10612 13716 10640 13756
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 12912 13793 12940 13824
rect 13814 13812 13820 13824
rect 13872 13852 13878 13864
rect 13924 13861 13952 13892
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 14660 13929 14688 13960
rect 16684 13932 16712 13960
rect 16936 13957 16948 13991
rect 16982 13988 16994 13991
rect 17034 13988 17040 14000
rect 16982 13960 17040 13988
rect 16982 13957 16994 13960
rect 16936 13951 16994 13957
rect 17034 13948 17040 13960
rect 17092 13948 17098 14000
rect 18432 13988 18460 14028
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 22649 14059 22707 14065
rect 20404 14028 22140 14056
rect 20404 14016 20410 14028
rect 17797 13960 18460 13988
rect 14918 13929 14924 13932
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14912 13920 14924 13929
rect 14879 13892 14924 13920
rect 14645 13883 14703 13889
rect 14912 13883 14924 13892
rect 14918 13880 14924 13883
rect 14976 13880 14982 13932
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 16666 13920 16672 13932
rect 15712 13892 16528 13920
rect 16627 13892 16672 13920
rect 15712 13880 15718 13892
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13872 13824 13921 13852
rect 13872 13812 13878 13824
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 13909 13815 13967 13821
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 14056 13824 14101 13852
rect 14056 13812 14062 13824
rect 15746 13812 15752 13864
rect 15804 13852 15810 13864
rect 16500 13852 16528 13892
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 17797 13920 17825 13960
rect 18506 13948 18512 14000
rect 18564 13988 18570 14000
rect 18564 13960 21036 13988
rect 18564 13948 18570 13960
rect 16776 13892 17825 13920
rect 16776 13852 16804 13892
rect 18046 13880 18052 13932
rect 18104 13920 18110 13932
rect 18598 13920 18604 13932
rect 18104 13892 18604 13920
rect 18104 13880 18110 13892
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 18877 13923 18935 13929
rect 18877 13889 18889 13923
rect 18923 13920 18935 13923
rect 19705 13923 19763 13929
rect 18923 13892 19012 13920
rect 18923 13889 18935 13892
rect 18877 13883 18935 13889
rect 15804 13824 16068 13852
rect 16500 13824 16804 13852
rect 15804 13812 15810 13824
rect 12897 13787 12955 13793
rect 12897 13753 12909 13787
rect 12943 13753 12955 13787
rect 12897 13747 12955 13753
rect 14458 13744 14464 13796
rect 14516 13784 14522 13796
rect 14642 13784 14648 13796
rect 14516 13756 14648 13784
rect 14516 13744 14522 13756
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 16040 13793 16068 13824
rect 18322 13812 18328 13864
rect 18380 13852 18386 13864
rect 18693 13855 18751 13861
rect 18693 13852 18705 13855
rect 18380 13824 18705 13852
rect 18380 13812 18386 13824
rect 18693 13821 18705 13824
rect 18739 13821 18751 13855
rect 18693 13815 18751 13821
rect 18785 13855 18843 13861
rect 18785 13821 18797 13855
rect 18831 13821 18843 13855
rect 18984 13852 19012 13892
rect 19705 13889 19717 13923
rect 19751 13910 19763 13923
rect 20070 13920 20076 13932
rect 19812 13910 20076 13920
rect 19751 13892 20076 13910
rect 19751 13889 19840 13892
rect 19705 13883 19840 13889
rect 19720 13882 19840 13883
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 20162 13880 20168 13932
rect 20220 13920 20226 13932
rect 20441 13923 20499 13929
rect 20441 13920 20453 13923
rect 20220 13892 20453 13920
rect 20220 13880 20226 13892
rect 20441 13889 20453 13892
rect 20487 13889 20499 13923
rect 20441 13883 20499 13889
rect 20530 13880 20536 13932
rect 20588 13920 20594 13932
rect 20717 13926 20775 13929
rect 20898 13926 20904 13932
rect 20717 13923 20904 13926
rect 20588 13892 20681 13920
rect 20588 13880 20594 13892
rect 20717 13889 20729 13923
rect 20763 13898 20904 13923
rect 20763 13889 20775 13898
rect 20717 13883 20775 13889
rect 20898 13880 20904 13898
rect 20956 13880 20962 13932
rect 21008 13920 21036 13960
rect 21082 13948 21088 14000
rect 21140 13988 21146 14000
rect 21821 13991 21879 13997
rect 21821 13988 21833 13991
rect 21140 13960 21833 13988
rect 21140 13948 21146 13960
rect 21821 13957 21833 13960
rect 21867 13957 21879 13991
rect 22021 13991 22079 13997
rect 22021 13988 22033 13991
rect 21821 13951 21879 13957
rect 21928 13960 22033 13988
rect 21928 13920 21956 13960
rect 22021 13957 22033 13960
rect 22067 13957 22079 13991
rect 22112 13988 22140 14028
rect 22649 14025 22661 14059
rect 22695 14056 22707 14059
rect 22695 14028 23336 14056
rect 22695 14025 22707 14028
rect 22649 14019 22707 14025
rect 22925 13991 22983 13997
rect 22925 13988 22937 13991
rect 22112 13960 22937 13988
rect 22021 13951 22079 13957
rect 22925 13957 22937 13960
rect 22971 13988 22983 13991
rect 23308 13988 23336 14028
rect 23382 14016 23388 14068
rect 23440 14056 23446 14068
rect 23483 14059 23541 14065
rect 23483 14056 23495 14059
rect 23440 14028 23495 14056
rect 23440 14016 23446 14028
rect 23483 14025 23495 14028
rect 23529 14025 23541 14059
rect 23483 14019 23541 14025
rect 23569 14059 23627 14065
rect 23569 14025 23581 14059
rect 23615 14056 23627 14059
rect 23750 14056 23756 14068
rect 23615 14028 23756 14056
rect 23615 14025 23627 14028
rect 23569 14019 23627 14025
rect 23750 14016 23756 14028
rect 23808 14056 23814 14068
rect 23808 14028 24624 14056
rect 23808 14016 23814 14028
rect 23934 13988 23940 14000
rect 22971 13960 23060 13988
rect 23308 13960 23940 13988
rect 22971 13957 22983 13960
rect 22925 13951 22983 13957
rect 21008 13892 21956 13920
rect 22646 13880 22652 13932
rect 22704 13929 22710 13932
rect 22704 13923 22729 13929
rect 22717 13889 22729 13923
rect 22704 13883 22729 13889
rect 22704 13880 22710 13883
rect 19426 13852 19432 13864
rect 18984 13824 19432 13852
rect 18785 13815 18843 13821
rect 16025 13787 16083 13793
rect 16025 13753 16037 13787
rect 16071 13753 16083 13787
rect 16025 13747 16083 13753
rect 18049 13787 18107 13793
rect 18049 13753 18061 13787
rect 18095 13784 18107 13787
rect 18598 13784 18604 13796
rect 18095 13756 18604 13784
rect 18095 13753 18107 13756
rect 18049 13747 18107 13753
rect 18598 13744 18604 13756
rect 18656 13744 18662 13796
rect 18800 13784 18828 13815
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 19981 13855 20039 13861
rect 19981 13852 19993 13855
rect 19812 13824 19993 13852
rect 18874 13784 18880 13796
rect 18800 13756 18880 13784
rect 18874 13744 18880 13756
rect 18932 13744 18938 13796
rect 19518 13744 19524 13796
rect 19576 13784 19582 13796
rect 19576 13756 19621 13784
rect 19576 13744 19582 13756
rect 19702 13744 19708 13796
rect 19760 13784 19766 13796
rect 19812 13784 19840 13824
rect 19981 13821 19993 13824
rect 20027 13821 20039 13855
rect 19981 13815 20039 13821
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 20548 13852 20576 13880
rect 20312 13824 20576 13852
rect 20312 13812 20318 13824
rect 21818 13812 21824 13864
rect 21876 13852 21882 13864
rect 21876 13824 22876 13852
rect 21876 13812 21882 13824
rect 19760 13756 19840 13784
rect 19889 13787 19947 13793
rect 19760 13744 19766 13756
rect 19889 13753 19901 13787
rect 19935 13784 19947 13787
rect 20162 13784 20168 13796
rect 19935 13756 20168 13784
rect 19935 13753 19947 13756
rect 19889 13747 19947 13753
rect 20162 13744 20168 13756
rect 20220 13744 20226 13796
rect 22094 13744 22100 13796
rect 22152 13784 22158 13796
rect 22741 13787 22799 13793
rect 22741 13784 22753 13787
rect 22152 13756 22753 13784
rect 22152 13744 22158 13756
rect 22741 13753 22753 13756
rect 22787 13753 22799 13787
rect 22741 13747 22799 13753
rect 10870 13716 10876 13728
rect 9232 13688 10640 13716
rect 10831 13688 10876 13716
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 13449 13719 13507 13725
rect 13449 13716 13461 13719
rect 12768 13688 13461 13716
rect 12768 13676 12774 13688
rect 13449 13685 13461 13688
rect 13495 13685 13507 13719
rect 13449 13679 13507 13685
rect 13538 13676 13544 13728
rect 13596 13716 13602 13728
rect 18138 13716 18144 13728
rect 13596 13688 18144 13716
rect 13596 13676 13602 13688
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 19058 13716 19064 13728
rect 19019 13688 19064 13716
rect 19058 13676 19064 13688
rect 19116 13676 19122 13728
rect 19150 13676 19156 13728
rect 19208 13716 19214 13728
rect 20901 13719 20959 13725
rect 20901 13716 20913 13719
rect 19208 13688 20913 13716
rect 19208 13676 19214 13688
rect 20901 13685 20913 13688
rect 20947 13685 20959 13719
rect 20901 13679 20959 13685
rect 21910 13676 21916 13728
rect 21968 13716 21974 13728
rect 22005 13719 22063 13725
rect 22005 13716 22017 13719
rect 21968 13688 22017 13716
rect 21968 13676 21974 13688
rect 22005 13685 22017 13688
rect 22051 13685 22063 13719
rect 22005 13679 22063 13685
rect 22189 13719 22247 13725
rect 22189 13685 22201 13719
rect 22235 13716 22247 13719
rect 22370 13716 22376 13728
rect 22235 13688 22376 13716
rect 22235 13685 22247 13688
rect 22189 13679 22247 13685
rect 22370 13676 22376 13688
rect 22428 13676 22434 13728
rect 22848 13716 22876 13824
rect 23032 13784 23060 13960
rect 23934 13948 23940 13960
rect 23992 13948 23998 14000
rect 23385 13923 23443 13929
rect 23385 13889 23397 13923
rect 23431 13889 23443 13923
rect 24121 13923 24179 13929
rect 23385 13883 23443 13889
rect 23670 13913 23728 13919
rect 23400 13852 23428 13883
rect 23670 13879 23682 13913
rect 23716 13910 23728 13913
rect 23716 13882 23796 13910
rect 24121 13889 24133 13923
rect 24167 13889 24179 13923
rect 24302 13920 24308 13932
rect 24263 13892 24308 13920
rect 24121 13883 24179 13889
rect 23716 13879 23728 13882
rect 23670 13873 23728 13879
rect 23400 13824 23520 13852
rect 23382 13784 23388 13796
rect 23032 13756 23388 13784
rect 23382 13744 23388 13756
rect 23440 13744 23446 13796
rect 23492 13716 23520 13824
rect 23566 13744 23572 13796
rect 23624 13784 23630 13796
rect 23768 13784 23796 13882
rect 23624 13756 23796 13784
rect 24136 13784 24164 13883
rect 24302 13880 24308 13892
rect 24360 13880 24366 13932
rect 24596 13852 24624 14028
rect 24670 14016 24676 14068
rect 24728 14056 24734 14068
rect 28077 14059 28135 14065
rect 28077 14056 28089 14059
rect 24728 14028 28089 14056
rect 24728 14016 24734 14028
rect 28077 14025 28089 14028
rect 28123 14025 28135 14059
rect 28077 14019 28135 14025
rect 28534 14016 28540 14068
rect 28592 14056 28598 14068
rect 28629 14059 28687 14065
rect 28629 14056 28641 14059
rect 28592 14028 28641 14056
rect 28592 14016 28598 14028
rect 28629 14025 28641 14028
rect 28675 14025 28687 14059
rect 29270 14056 29276 14068
rect 29231 14028 29276 14056
rect 28629 14019 28687 14025
rect 29270 14016 29276 14028
rect 29328 14016 29334 14068
rect 30834 14056 30840 14068
rect 30795 14028 30840 14056
rect 30834 14016 30840 14028
rect 30892 14016 30898 14068
rect 25314 13988 25320 14000
rect 25275 13960 25320 13988
rect 25314 13948 25320 13960
rect 25372 13948 25378 14000
rect 25682 13948 25688 14000
rect 25740 13988 25746 14000
rect 25869 13991 25927 13997
rect 25869 13988 25881 13991
rect 25740 13960 25881 13988
rect 25740 13948 25746 13960
rect 25869 13957 25881 13960
rect 25915 13957 25927 13991
rect 27522 13988 27528 14000
rect 27483 13960 27528 13988
rect 25869 13951 25927 13957
rect 27522 13948 27528 13960
rect 27580 13988 27586 14000
rect 28350 13988 28356 14000
rect 27580 13960 28356 13988
rect 27580 13948 27586 13960
rect 28350 13948 28356 13960
rect 28408 13948 28414 14000
rect 24857 13923 24915 13929
rect 24857 13889 24869 13923
rect 24903 13920 24915 13923
rect 26142 13920 26148 13932
rect 24903 13892 26148 13920
rect 24903 13889 24915 13892
rect 24857 13883 24915 13889
rect 26142 13880 26148 13892
rect 26200 13880 26206 13932
rect 30285 13923 30343 13929
rect 30285 13920 30297 13923
rect 26988 13892 30297 13920
rect 26988 13864 27016 13892
rect 30285 13889 30297 13892
rect 30331 13889 30343 13923
rect 30285 13883 30343 13889
rect 26970 13852 26976 13864
rect 24596 13824 26976 13852
rect 26970 13812 26976 13824
rect 27028 13812 27034 13864
rect 28994 13812 29000 13864
rect 29052 13852 29058 13864
rect 29733 13855 29791 13861
rect 29733 13852 29745 13855
rect 29052 13824 29745 13852
rect 29052 13812 29058 13824
rect 29733 13821 29745 13824
rect 29779 13821 29791 13855
rect 29733 13815 29791 13821
rect 28534 13784 28540 13796
rect 24136 13756 28540 13784
rect 23624 13744 23630 13756
rect 28534 13744 28540 13756
rect 28592 13744 28598 13796
rect 22848 13688 23520 13716
rect 23658 13676 23664 13728
rect 23716 13716 23722 13728
rect 24121 13719 24179 13725
rect 24121 13716 24133 13719
rect 23716 13688 24133 13716
rect 23716 13676 23722 13688
rect 24121 13685 24133 13688
rect 24167 13685 24179 13719
rect 24121 13679 24179 13685
rect 25222 13676 25228 13728
rect 25280 13716 25286 13728
rect 25958 13716 25964 13728
rect 25280 13688 25964 13716
rect 25280 13676 25286 13688
rect 25958 13676 25964 13688
rect 26016 13676 26022 13728
rect 1104 13626 44896 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 44896 13626
rect 1104 13552 44896 13574
rect 1673 13515 1731 13521
rect 1673 13481 1685 13515
rect 1719 13512 1731 13515
rect 1762 13512 1768 13524
rect 1719 13484 1768 13512
rect 1719 13481 1731 13484
rect 1673 13475 1731 13481
rect 1762 13472 1768 13484
rect 1820 13472 1826 13524
rect 1872 13484 3740 13512
rect 842 13404 848 13456
rect 900 13444 906 13456
rect 1872 13444 1900 13484
rect 900 13416 1900 13444
rect 900 13404 906 13416
rect 2038 13404 2044 13456
rect 2096 13444 2102 13456
rect 2222 13444 2228 13456
rect 2096 13416 2228 13444
rect 2096 13404 2102 13416
rect 2222 13404 2228 13416
rect 2280 13404 2286 13456
rect 2314 13404 2320 13456
rect 2372 13444 2378 13456
rect 2498 13444 2504 13456
rect 2372 13416 2504 13444
rect 2372 13404 2378 13416
rect 2498 13404 2504 13416
rect 2556 13404 2562 13456
rect 3326 13444 3332 13456
rect 2700 13416 3332 13444
rect 1486 13376 1492 13388
rect 1447 13348 1492 13376
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 2700 13385 2728 13416
rect 3326 13404 3332 13416
rect 3384 13404 3390 13456
rect 3712 13444 3740 13484
rect 3878 13472 3884 13524
rect 3936 13512 3942 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 3936 13484 4077 13512
rect 3936 13472 3942 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 4249 13515 4307 13521
rect 4249 13481 4261 13515
rect 4295 13512 4307 13515
rect 5350 13512 5356 13524
rect 4295 13484 5356 13512
rect 4295 13481 4307 13484
rect 4249 13475 4307 13481
rect 4080 13444 4108 13475
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 9674 13512 9680 13524
rect 6236 13484 9680 13512
rect 6236 13472 6242 13484
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 13998 13512 14004 13524
rect 9784 13484 14004 13512
rect 4154 13444 4160 13456
rect 3712 13416 4016 13444
rect 4080 13416 4160 13444
rect 2685 13379 2743 13385
rect 1596 13348 2544 13376
rect 1210 13268 1216 13320
rect 1268 13308 1274 13320
rect 1596 13308 1624 13348
rect 1268 13280 1624 13308
rect 1673 13311 1731 13317
rect 1268 13268 1274 13280
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 2038 13308 2044 13320
rect 1719 13280 2044 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 1394 13240 1400 13252
rect 1355 13212 1400 13240
rect 1394 13200 1400 13212
rect 1452 13200 1458 13252
rect 1486 13200 1492 13252
rect 1544 13240 1550 13252
rect 2314 13240 2320 13252
rect 1544 13212 2320 13240
rect 1544 13200 1550 13212
rect 2314 13200 2320 13212
rect 2372 13200 2378 13252
rect 2516 13240 2544 13348
rect 2685 13345 2697 13379
rect 2731 13345 2743 13379
rect 2685 13339 2743 13345
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 3878 13376 3884 13388
rect 2832 13348 2877 13376
rect 3839 13348 3884 13376
rect 2832 13336 2838 13348
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 2866 13308 2872 13320
rect 2827 13280 2872 13308
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 3786 13308 3792 13320
rect 3747 13280 3792 13308
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 3988 13240 4016 13416
rect 4154 13404 4160 13416
rect 4212 13404 4218 13456
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 9490 13444 9496 13456
rect 6972 13416 9496 13444
rect 6972 13404 6978 13416
rect 9490 13404 9496 13416
rect 9548 13404 9554 13456
rect 6549 13379 6607 13385
rect 6549 13345 6561 13379
rect 6595 13376 6607 13379
rect 8202 13376 8208 13388
rect 6595 13348 8208 13376
rect 6595 13345 6607 13348
rect 6549 13339 6607 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 8846 13336 8852 13388
rect 8904 13376 8910 13388
rect 9784 13376 9812 13484
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 16298 13472 16304 13524
rect 16356 13512 16362 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 16356 13484 19257 13512
rect 16356 13472 16362 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 19426 13472 19432 13524
rect 19484 13512 19490 13524
rect 21266 13512 21272 13524
rect 19484 13484 21272 13512
rect 19484 13472 19490 13484
rect 21266 13472 21272 13484
rect 21324 13472 21330 13524
rect 22094 13472 22100 13524
rect 22152 13512 22158 13524
rect 22370 13512 22376 13524
rect 22152 13484 22376 13512
rect 22152 13472 22158 13484
rect 22370 13472 22376 13484
rect 22428 13472 22434 13524
rect 22554 13472 22560 13524
rect 22612 13512 22618 13524
rect 22649 13515 22707 13521
rect 22649 13512 22661 13515
rect 22612 13484 22661 13512
rect 22612 13472 22618 13484
rect 22649 13481 22661 13484
rect 22695 13481 22707 13515
rect 22649 13475 22707 13481
rect 23385 13515 23443 13521
rect 23385 13481 23397 13515
rect 23431 13512 23443 13515
rect 23842 13512 23848 13524
rect 23431 13484 23848 13512
rect 23431 13481 23443 13484
rect 23385 13475 23443 13481
rect 23842 13472 23848 13484
rect 23900 13472 23906 13524
rect 25041 13515 25099 13521
rect 25041 13481 25053 13515
rect 25087 13512 25099 13515
rect 25314 13512 25320 13524
rect 25087 13484 25320 13512
rect 25087 13481 25099 13484
rect 25041 13475 25099 13481
rect 25314 13472 25320 13484
rect 25372 13472 25378 13524
rect 25498 13472 25504 13524
rect 25556 13512 25562 13524
rect 26053 13515 26111 13521
rect 26053 13512 26065 13515
rect 25556 13484 26065 13512
rect 25556 13472 25562 13484
rect 26053 13481 26065 13484
rect 26099 13481 26111 13515
rect 26053 13475 26111 13481
rect 27249 13515 27307 13521
rect 27249 13481 27261 13515
rect 27295 13512 27307 13515
rect 27614 13512 27620 13524
rect 27295 13484 27620 13512
rect 27295 13481 27307 13484
rect 27249 13475 27307 13481
rect 27614 13472 27620 13484
rect 27672 13472 27678 13524
rect 28258 13512 28264 13524
rect 28219 13484 28264 13512
rect 28258 13472 28264 13484
rect 28316 13472 28322 13524
rect 28350 13472 28356 13524
rect 28408 13512 28414 13524
rect 30101 13515 30159 13521
rect 30101 13512 30113 13515
rect 28408 13484 30113 13512
rect 28408 13472 28414 13484
rect 30101 13481 30113 13484
rect 30147 13481 30159 13515
rect 30101 13475 30159 13481
rect 12250 13404 12256 13456
rect 12308 13444 12314 13456
rect 13541 13447 13599 13453
rect 13541 13444 13553 13447
rect 12308 13416 13553 13444
rect 12308 13404 12314 13416
rect 13541 13413 13553 13416
rect 13587 13413 13599 13447
rect 13541 13407 13599 13413
rect 17402 13404 17408 13456
rect 17460 13444 17466 13456
rect 18325 13447 18383 13453
rect 18325 13444 18337 13447
rect 17460 13416 18337 13444
rect 17460 13404 17466 13416
rect 18325 13413 18337 13416
rect 18371 13444 18383 13447
rect 19518 13444 19524 13456
rect 18371 13416 19524 13444
rect 18371 13413 18383 13416
rect 18325 13407 18383 13413
rect 19518 13404 19524 13416
rect 19576 13404 19582 13456
rect 20622 13444 20628 13456
rect 19628 13416 20628 13444
rect 8904 13348 9812 13376
rect 8904 13336 8910 13348
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 12710 13376 12716 13388
rect 12400 13348 12716 13376
rect 12400 13336 12406 13348
rect 12710 13336 12716 13348
rect 12768 13336 12774 13388
rect 17862 13336 17868 13388
rect 17920 13376 17926 13388
rect 18874 13376 18880 13388
rect 17920 13348 18460 13376
rect 17920 13336 17926 13348
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4120 13280 4165 13308
rect 4120 13268 4126 13280
rect 4614 13268 4620 13320
rect 4672 13308 4678 13320
rect 4709 13311 4767 13317
rect 4709 13308 4721 13311
rect 4672 13280 4721 13308
rect 4672 13268 4678 13280
rect 4709 13277 4721 13280
rect 4755 13277 4767 13311
rect 4709 13271 4767 13277
rect 10778 13268 10784 13320
rect 10836 13308 10842 13320
rect 11238 13308 11244 13320
rect 10836 13280 10881 13308
rect 11199 13280 11244 13308
rect 10836 13268 10842 13280
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 12406 13280 13369 13308
rect 4954 13243 5012 13249
rect 4954 13240 4966 13243
rect 2516 13212 3280 13240
rect 3988 13212 4966 13240
rect 1857 13175 1915 13181
rect 1857 13141 1869 13175
rect 1903 13172 1915 13175
rect 2498 13172 2504 13184
rect 1903 13144 2504 13172
rect 1903 13141 1915 13144
rect 1857 13135 1915 13141
rect 2498 13132 2504 13144
rect 2556 13132 2562 13184
rect 3252 13181 3280 13212
rect 4954 13209 4966 13212
rect 5000 13209 5012 13243
rect 4954 13203 5012 13209
rect 6546 13200 6552 13252
rect 6604 13240 6610 13252
rect 6733 13243 6791 13249
rect 6733 13240 6745 13243
rect 6604 13212 6745 13240
rect 6604 13200 6610 13212
rect 6733 13209 6745 13212
rect 6779 13209 6791 13243
rect 6733 13203 6791 13209
rect 8389 13243 8447 13249
rect 8389 13209 8401 13243
rect 8435 13209 8447 13243
rect 8389 13203 8447 13209
rect 3237 13175 3295 13181
rect 3237 13141 3249 13175
rect 3283 13141 3295 13175
rect 3237 13135 3295 13141
rect 3786 13132 3792 13184
rect 3844 13172 3850 13184
rect 8294 13172 8300 13184
rect 3844 13144 8300 13172
rect 3844 13132 3850 13144
rect 8294 13132 8300 13144
rect 8352 13172 8358 13184
rect 8404 13172 8432 13203
rect 8570 13200 8576 13252
rect 8628 13240 8634 13252
rect 8941 13243 8999 13249
rect 8941 13240 8953 13243
rect 8628 13212 8953 13240
rect 8628 13200 8634 13212
rect 8941 13209 8953 13212
rect 8987 13209 8999 13243
rect 8941 13203 8999 13209
rect 10410 13200 10416 13252
rect 10468 13240 10474 13252
rect 10597 13243 10655 13249
rect 10597 13240 10609 13243
rect 10468 13212 10609 13240
rect 10468 13200 10474 13212
rect 10597 13209 10609 13212
rect 10643 13209 10655 13243
rect 10597 13203 10655 13209
rect 10870 13200 10876 13252
rect 10928 13240 10934 13252
rect 11486 13243 11544 13249
rect 11486 13240 11498 13243
rect 10928 13212 11498 13240
rect 10928 13200 10934 13212
rect 11486 13209 11498 13212
rect 11532 13209 11544 13243
rect 11486 13203 11544 13209
rect 8352 13144 8432 13172
rect 8352 13132 8358 13144
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 11698 13172 11704 13184
rect 8812 13144 11704 13172
rect 8812 13132 8818 13144
rect 11698 13132 11704 13144
rect 11756 13172 11762 13184
rect 12406 13172 12434 13280
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 14090 13308 14096 13320
rect 14003 13280 14096 13308
rect 13357 13271 13415 13277
rect 14090 13268 14096 13280
rect 14148 13308 14154 13320
rect 14826 13308 14832 13320
rect 14148 13280 14832 13308
rect 14148 13268 14154 13280
rect 14826 13268 14832 13280
rect 14884 13308 14890 13320
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 14884 13280 15945 13308
rect 14884 13268 14890 13280
rect 15933 13277 15945 13280
rect 15979 13308 15991 13311
rect 16666 13308 16672 13320
rect 15979 13280 16672 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18156 13308 18276 13310
rect 18322 13308 18328 13320
rect 18003 13282 18328 13308
rect 18003 13280 18184 13282
rect 18248 13280 18328 13282
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 12710 13200 12716 13252
rect 12768 13240 12774 13252
rect 13173 13243 13231 13249
rect 13173 13240 13185 13243
rect 12768 13212 13185 13240
rect 12768 13200 12774 13212
rect 13173 13209 13185 13212
rect 13219 13209 13231 13243
rect 13173 13203 13231 13209
rect 14360 13243 14418 13249
rect 14360 13209 14372 13243
rect 14406 13240 14418 13243
rect 15102 13240 15108 13252
rect 14406 13212 15108 13240
rect 14406 13209 14418 13212
rect 14360 13203 14418 13209
rect 15102 13200 15108 13212
rect 15160 13200 15166 13252
rect 15194 13200 15200 13252
rect 15252 13240 15258 13252
rect 16178 13243 16236 13249
rect 16178 13240 16190 13243
rect 15252 13212 16190 13240
rect 15252 13200 15258 13212
rect 16178 13209 16190 13212
rect 16224 13209 16236 13243
rect 16178 13203 16236 13209
rect 18049 13243 18107 13249
rect 18049 13209 18061 13243
rect 18095 13240 18107 13243
rect 18432 13240 18460 13348
rect 18524 13348 18880 13376
rect 18524 13320 18552 13348
rect 18874 13336 18880 13348
rect 18932 13376 18938 13388
rect 19628 13376 19656 13416
rect 20622 13404 20628 13416
rect 20680 13404 20686 13456
rect 21910 13444 21916 13456
rect 21284 13416 21916 13444
rect 18932 13348 19656 13376
rect 18932 13336 18938 13348
rect 19702 13336 19708 13388
rect 19760 13376 19766 13388
rect 21082 13376 21088 13388
rect 19760 13348 21088 13376
rect 19760 13336 19766 13348
rect 21082 13336 21088 13348
rect 21140 13336 21146 13388
rect 18506 13268 18512 13320
rect 18564 13268 18570 13320
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 18892 13280 19441 13308
rect 18892 13252 18920 13280
rect 19429 13277 19441 13280
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 18095 13212 18828 13240
rect 18095 13209 18107 13212
rect 18049 13203 18107 13209
rect 11756 13144 12434 13172
rect 12621 13175 12679 13181
rect 11756 13132 11762 13144
rect 12621 13141 12633 13175
rect 12667 13172 12679 13175
rect 12986 13172 12992 13184
rect 12667 13144 12992 13172
rect 12667 13141 12679 13144
rect 12621 13135 12679 13141
rect 12986 13132 12992 13144
rect 13044 13172 13050 13184
rect 13446 13172 13452 13184
rect 13044 13144 13452 13172
rect 13044 13132 13050 13144
rect 13446 13132 13452 13144
rect 13504 13172 13510 13184
rect 14274 13172 14280 13184
rect 13504 13144 14280 13172
rect 13504 13132 13510 13144
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 15473 13175 15531 13181
rect 15473 13141 15485 13175
rect 15519 13172 15531 13175
rect 16298 13172 16304 13184
rect 15519 13144 16304 13172
rect 15519 13141 15531 13144
rect 15473 13135 15531 13141
rect 16298 13132 16304 13144
rect 16356 13132 16362 13184
rect 17218 13132 17224 13184
rect 17276 13172 17282 13184
rect 17313 13175 17371 13181
rect 17313 13172 17325 13175
rect 17276 13144 17325 13172
rect 17276 13132 17282 13144
rect 17313 13141 17325 13144
rect 17359 13141 17371 13175
rect 17313 13135 17371 13141
rect 17402 13132 17408 13184
rect 17460 13172 17466 13184
rect 17773 13175 17831 13181
rect 17773 13172 17785 13175
rect 17460 13144 17785 13172
rect 17460 13132 17466 13144
rect 17773 13141 17785 13144
rect 17819 13141 17831 13175
rect 17773 13135 17831 13141
rect 18138 13132 18144 13184
rect 18196 13172 18202 13184
rect 18800 13172 18828 13212
rect 18874 13200 18880 13252
rect 18932 13200 18938 13252
rect 19628 13240 19656 13271
rect 20254 13268 20260 13320
rect 20312 13308 20318 13320
rect 20349 13311 20407 13317
rect 20349 13308 20361 13311
rect 20312 13280 20361 13308
rect 20312 13268 20318 13280
rect 20349 13277 20361 13280
rect 20395 13277 20407 13311
rect 20622 13308 20628 13320
rect 20583 13280 20628 13308
rect 20349 13271 20407 13277
rect 20622 13268 20628 13280
rect 20680 13268 20686 13320
rect 21284 13317 21312 13416
rect 21910 13404 21916 13416
rect 21968 13444 21974 13456
rect 26697 13447 26755 13453
rect 26697 13444 26709 13447
rect 21968 13416 26709 13444
rect 21968 13404 21974 13416
rect 26697 13413 26709 13416
rect 26743 13444 26755 13447
rect 28905 13447 28963 13453
rect 28905 13444 28917 13447
rect 26743 13416 28917 13444
rect 26743 13413 26755 13416
rect 26697 13407 26755 13413
rect 28905 13413 28917 13416
rect 28951 13444 28963 13447
rect 28994 13444 29000 13456
rect 28951 13416 29000 13444
rect 28951 13413 28963 13416
rect 28905 13407 28963 13413
rect 28994 13404 29000 13416
rect 29052 13404 29058 13456
rect 21358 13336 21364 13388
rect 21416 13376 21422 13388
rect 21416 13348 23612 13376
rect 21416 13336 21422 13348
rect 21269 13311 21327 13317
rect 21269 13277 21281 13311
rect 21315 13277 21327 13311
rect 22925 13311 22983 13317
rect 21269 13271 21327 13277
rect 22296 13280 22876 13308
rect 21284 13240 21312 13271
rect 21450 13240 21456 13252
rect 19628 13212 21312 13240
rect 21411 13212 21456 13240
rect 19628 13172 19656 13212
rect 21450 13200 21456 13212
rect 21508 13200 21514 13252
rect 21726 13200 21732 13252
rect 21784 13240 21790 13252
rect 21910 13240 21916 13252
rect 21784 13212 21916 13240
rect 21784 13200 21790 13212
rect 21910 13200 21916 13212
rect 21968 13240 21974 13252
rect 22005 13243 22063 13249
rect 22005 13240 22017 13243
rect 21968 13212 22017 13240
rect 21968 13200 21974 13212
rect 22005 13209 22017 13212
rect 22051 13209 22063 13243
rect 22005 13203 22063 13209
rect 18196 13144 18241 13172
rect 18800 13144 19656 13172
rect 18196 13132 18202 13144
rect 20070 13132 20076 13184
rect 20128 13172 20134 13184
rect 20165 13175 20223 13181
rect 20165 13172 20177 13175
rect 20128 13144 20177 13172
rect 20128 13132 20134 13144
rect 20165 13141 20177 13144
rect 20211 13141 20223 13175
rect 20165 13135 20223 13141
rect 20533 13175 20591 13181
rect 20533 13141 20545 13175
rect 20579 13172 20591 13175
rect 20714 13172 20720 13184
rect 20579 13144 20720 13172
rect 20579 13141 20591 13144
rect 20533 13135 20591 13141
rect 20714 13132 20720 13144
rect 20772 13172 20778 13184
rect 22296 13172 22324 13280
rect 22554 13200 22560 13252
rect 22612 13240 22618 13252
rect 22848 13249 22876 13280
rect 22925 13277 22937 13311
rect 22971 13308 22983 13311
rect 23198 13308 23204 13320
rect 22971 13280 23204 13308
rect 22971 13277 22983 13280
rect 22925 13271 22983 13277
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 23584 13317 23612 13348
rect 24762 13336 24768 13388
rect 24820 13376 24826 13388
rect 25501 13379 25559 13385
rect 25501 13376 25513 13379
rect 24820 13348 25513 13376
rect 24820 13336 24826 13348
rect 25501 13345 25513 13348
rect 25547 13376 25559 13379
rect 26050 13376 26056 13388
rect 25547 13348 26056 13376
rect 25547 13345 25559 13348
rect 25501 13339 25559 13345
rect 26050 13336 26056 13348
rect 26108 13336 26114 13388
rect 27890 13336 27896 13388
rect 27948 13376 27954 13388
rect 28258 13376 28264 13388
rect 27948 13348 28264 13376
rect 27948 13336 27954 13348
rect 28258 13336 28264 13348
rect 28316 13336 28322 13388
rect 23569 13311 23627 13317
rect 23569 13277 23581 13311
rect 23615 13277 23627 13311
rect 24486 13308 24492 13320
rect 24399 13280 24492 13308
rect 23569 13271 23627 13277
rect 24486 13268 24492 13280
rect 24544 13308 24550 13320
rect 26326 13308 26332 13320
rect 24544 13280 26332 13308
rect 24544 13268 24550 13280
rect 26326 13268 26332 13280
rect 26384 13268 26390 13320
rect 22649 13243 22707 13249
rect 22649 13240 22661 13243
rect 22612 13212 22661 13240
rect 22612 13200 22618 13212
rect 22649 13209 22661 13212
rect 22695 13209 22707 13243
rect 22649 13203 22707 13209
rect 22833 13243 22891 13249
rect 22833 13209 22845 13243
rect 22879 13240 22891 13243
rect 26142 13240 26148 13252
rect 22879 13212 26148 13240
rect 22879 13209 22891 13212
rect 22833 13203 22891 13209
rect 20772 13144 22324 13172
rect 22664 13172 22692 13203
rect 26142 13200 26148 13212
rect 26200 13200 26206 13252
rect 26694 13200 26700 13252
rect 26752 13240 26758 13252
rect 27709 13243 27767 13249
rect 27709 13240 27721 13243
rect 26752 13212 27721 13240
rect 26752 13200 26758 13212
rect 27709 13209 27721 13212
rect 27755 13209 27767 13243
rect 27709 13203 27767 13209
rect 24302 13172 24308 13184
rect 22664 13144 24308 13172
rect 20772 13132 20778 13144
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 27522 13132 27528 13184
rect 27580 13172 27586 13184
rect 29549 13175 29607 13181
rect 29549 13172 29561 13175
rect 27580 13144 29561 13172
rect 27580 13132 27586 13144
rect 29549 13141 29561 13144
rect 29595 13141 29607 13175
rect 29549 13135 29607 13141
rect 29638 13132 29644 13184
rect 29696 13172 29702 13184
rect 30653 13175 30711 13181
rect 30653 13172 30665 13175
rect 29696 13144 30665 13172
rect 29696 13132 29702 13144
rect 30653 13141 30665 13144
rect 30699 13141 30711 13175
rect 30653 13135 30711 13141
rect 1104 13082 44896 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 44896 13082
rect 1104 13008 44896 13030
rect 1857 12971 1915 12977
rect 1857 12937 1869 12971
rect 1903 12968 1915 12971
rect 2130 12968 2136 12980
rect 1903 12940 2136 12968
rect 1903 12937 1915 12940
rect 1857 12931 1915 12937
rect 2130 12928 2136 12940
rect 2188 12928 2194 12980
rect 3510 12968 3516 12980
rect 3471 12940 3516 12968
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 6086 12928 6092 12980
rect 6144 12968 6150 12980
rect 7837 12971 7895 12977
rect 6144 12940 7236 12968
rect 6144 12928 6150 12940
rect 2222 12900 2228 12912
rect 1596 12872 2228 12900
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12832 1455 12835
rect 1486 12832 1492 12844
rect 1443 12804 1492 12832
rect 1443 12801 1455 12804
rect 1397 12795 1455 12801
rect 1486 12792 1492 12804
rect 1544 12792 1550 12844
rect 1596 12841 1624 12872
rect 2222 12860 2228 12872
rect 2280 12900 2286 12912
rect 2866 12900 2872 12912
rect 2280 12872 2872 12900
rect 2280 12860 2286 12872
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 3602 12900 3608 12912
rect 3563 12872 3608 12900
rect 3602 12860 3608 12872
rect 3660 12900 3666 12912
rect 6178 12900 6184 12912
rect 3660 12872 6184 12900
rect 3660 12860 3666 12872
rect 6178 12860 6184 12872
rect 6236 12860 6242 12912
rect 6822 12900 6828 12912
rect 6472 12872 6828 12900
rect 6472 12844 6500 12872
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12801 1639 12835
rect 1581 12795 1639 12801
rect 1670 12792 1676 12844
rect 1728 12832 1734 12844
rect 2501 12835 2559 12841
rect 1728 12804 1773 12832
rect 1728 12792 1734 12804
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 2590 12832 2596 12844
rect 2547 12804 2596 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 2590 12792 2596 12804
rect 2648 12792 2654 12844
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 4062 12832 4068 12844
rect 2823 12804 4068 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12832 4491 12835
rect 4522 12832 4528 12844
rect 4479 12804 4528 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 4706 12841 4712 12844
rect 4700 12795 4712 12841
rect 4764 12832 4770 12844
rect 6454 12832 6460 12844
rect 4764 12804 4800 12832
rect 6415 12804 6460 12832
rect 4706 12792 4712 12795
rect 4764 12792 4770 12804
rect 6454 12792 6460 12804
rect 6512 12792 6518 12844
rect 6730 12841 6736 12844
rect 6724 12832 6736 12841
rect 6691 12804 6736 12832
rect 6724 12795 6736 12804
rect 6730 12792 6736 12795
rect 6788 12792 6794 12844
rect 7208 12832 7236 12940
rect 7837 12937 7849 12971
rect 7883 12968 7895 12971
rect 9674 12968 9680 12980
rect 7883 12940 9680 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 10318 12928 10324 12980
rect 10376 12968 10382 12980
rect 15519 12971 15577 12977
rect 15519 12968 15531 12971
rect 10376 12940 15531 12968
rect 10376 12928 10382 12940
rect 15519 12937 15531 12940
rect 15565 12937 15577 12971
rect 15519 12931 15577 12937
rect 15930 12928 15936 12980
rect 15988 12968 15994 12980
rect 16206 12968 16212 12980
rect 15988 12940 16212 12968
rect 15988 12928 15994 12940
rect 16206 12928 16212 12940
rect 16264 12928 16270 12980
rect 16574 12928 16580 12980
rect 16632 12968 16638 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 16632 12940 16681 12968
rect 16632 12928 16638 12940
rect 16669 12937 16681 12940
rect 16715 12968 16727 12971
rect 18322 12968 18328 12980
rect 16715 12940 18328 12968
rect 16715 12937 16727 12940
rect 16669 12931 16727 12937
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 19150 12968 19156 12980
rect 18748 12940 19156 12968
rect 18748 12928 18754 12940
rect 19150 12928 19156 12940
rect 19208 12928 19214 12980
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19587 12971 19645 12977
rect 19587 12968 19599 12971
rect 19392 12940 19599 12968
rect 19392 12928 19398 12940
rect 19587 12937 19599 12940
rect 19633 12937 19645 12971
rect 20714 12968 20720 12980
rect 19587 12931 19645 12937
rect 19812 12940 20720 12968
rect 8478 12900 8484 12912
rect 8439 12872 8484 12900
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 14584 12903 14642 12909
rect 14584 12869 14596 12903
rect 14630 12900 14642 12903
rect 18509 12903 18567 12909
rect 18509 12900 18521 12903
rect 14630 12872 18521 12900
rect 14630 12869 14642 12872
rect 14584 12863 14642 12869
rect 18509 12869 18521 12872
rect 18555 12869 18567 12903
rect 19242 12900 19248 12912
rect 18509 12863 18567 12869
rect 18984 12872 19248 12900
rect 7926 12832 7932 12844
rect 7208 12804 7932 12832
rect 7926 12792 7932 12804
rect 7984 12832 7990 12844
rect 8297 12835 8355 12841
rect 8297 12832 8309 12835
rect 7984 12804 8309 12832
rect 7984 12792 7990 12804
rect 8297 12801 8309 12804
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 9950 12792 9956 12844
rect 10008 12832 10014 12844
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10008 12804 10793 12832
rect 10008 12792 10014 12804
rect 10781 12801 10793 12804
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 12722 12835 12780 12841
rect 12722 12832 12734 12835
rect 11112 12804 12734 12832
rect 11112 12792 11118 12804
rect 12722 12801 12734 12804
rect 12768 12801 12780 12835
rect 12722 12795 12780 12801
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 14090 12832 14096 12844
rect 13035 12804 14096 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 15286 12832 15292 12844
rect 14884 12804 14929 12832
rect 15247 12804 15292 12832
rect 14884 12792 14890 12804
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 15470 12792 15476 12844
rect 15528 12832 15534 12844
rect 17402 12832 17408 12844
rect 15528 12804 17408 12832
rect 15528 12792 15534 12804
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 17782 12835 17840 12841
rect 17782 12832 17794 12835
rect 17552 12804 17794 12832
rect 17552 12792 17558 12804
rect 17782 12801 17794 12804
rect 17828 12801 17840 12835
rect 17782 12795 17840 12801
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18984 12841 19012 12872
rect 19242 12860 19248 12872
rect 19300 12860 19306 12912
rect 19702 12860 19708 12912
rect 19760 12900 19766 12912
rect 19812 12909 19840 12940
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 23017 12971 23075 12977
rect 23017 12937 23029 12971
rect 23063 12968 23075 12971
rect 23474 12968 23480 12980
rect 23063 12940 23480 12968
rect 23063 12937 23075 12940
rect 23017 12931 23075 12937
rect 23474 12928 23480 12940
rect 23532 12928 23538 12980
rect 23658 12928 23664 12980
rect 23716 12968 23722 12980
rect 24762 12968 24768 12980
rect 23716 12940 24768 12968
rect 23716 12928 23722 12940
rect 24762 12928 24768 12940
rect 24820 12968 24826 12980
rect 25958 12968 25964 12980
rect 24820 12940 25544 12968
rect 25919 12940 25964 12968
rect 24820 12928 24826 12940
rect 19797 12903 19855 12909
rect 19797 12900 19809 12903
rect 19760 12872 19809 12900
rect 19760 12860 19766 12872
rect 19797 12869 19809 12872
rect 19843 12869 19855 12903
rect 19797 12863 19855 12869
rect 19978 12860 19984 12912
rect 20036 12900 20042 12912
rect 20257 12903 20315 12909
rect 20257 12900 20269 12903
rect 20036 12872 20269 12900
rect 20036 12860 20042 12872
rect 20257 12869 20269 12872
rect 20303 12869 20315 12903
rect 20257 12863 20315 12869
rect 20473 12903 20531 12909
rect 20473 12869 20485 12903
rect 20519 12900 20531 12903
rect 20622 12900 20628 12912
rect 20519 12872 20628 12900
rect 20519 12869 20531 12872
rect 20473 12863 20531 12869
rect 20622 12860 20628 12872
rect 20680 12860 20686 12912
rect 21174 12900 21180 12912
rect 21135 12872 21180 12900
rect 21174 12860 21180 12872
rect 21232 12860 21238 12912
rect 22373 12903 22431 12909
rect 22373 12869 22385 12903
rect 22419 12900 22431 12903
rect 22554 12900 22560 12912
rect 22419 12872 22560 12900
rect 22419 12869 22431 12872
rect 22373 12863 22431 12869
rect 22554 12860 22560 12872
rect 22612 12900 22618 12912
rect 24486 12900 24492 12912
rect 22612 12872 24492 12900
rect 22612 12860 22618 12872
rect 24486 12860 24492 12872
rect 24544 12860 24550 12912
rect 25516 12909 25544 12940
rect 25958 12928 25964 12940
rect 26016 12928 26022 12980
rect 26142 12928 26148 12980
rect 26200 12968 26206 12980
rect 28166 12968 28172 12980
rect 26200 12940 27936 12968
rect 28127 12940 28172 12968
rect 26200 12928 26206 12940
rect 25501 12903 25559 12909
rect 25501 12869 25513 12903
rect 25547 12900 25559 12903
rect 26510 12900 26516 12912
rect 25547 12872 26516 12900
rect 25547 12869 25559 12872
rect 25501 12863 25559 12869
rect 26510 12860 26516 12872
rect 26568 12860 26574 12912
rect 27614 12860 27620 12912
rect 27672 12900 27678 12912
rect 27798 12900 27804 12912
rect 27672 12872 27804 12900
rect 27672 12860 27678 12872
rect 27798 12860 27804 12872
rect 27856 12860 27862 12912
rect 27908 12900 27936 12940
rect 28166 12928 28172 12940
rect 28224 12928 28230 12980
rect 28721 12971 28779 12977
rect 28721 12937 28733 12971
rect 28767 12968 28779 12971
rect 28994 12968 29000 12980
rect 28767 12940 29000 12968
rect 28767 12937 28779 12940
rect 28721 12931 28779 12937
rect 28994 12928 29000 12940
rect 29052 12928 29058 12980
rect 29273 12971 29331 12977
rect 29273 12937 29285 12971
rect 29319 12968 29331 12971
rect 29638 12968 29644 12980
rect 29319 12940 29644 12968
rect 29319 12937 29331 12940
rect 29273 12931 29331 12937
rect 28902 12900 28908 12912
rect 27908 12872 28908 12900
rect 28902 12860 28908 12872
rect 28960 12900 28966 12912
rect 29288 12900 29316 12931
rect 29638 12928 29644 12940
rect 29696 12928 29702 12980
rect 28960 12872 29316 12900
rect 28960 12860 28966 12872
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 18012 12804 18705 12832
rect 18012 12792 18018 12804
rect 18693 12801 18705 12804
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 18969 12835 19027 12841
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 19058 12792 19064 12844
rect 19116 12832 19122 12844
rect 21085 12835 21143 12841
rect 21085 12832 21097 12835
rect 19116 12804 21097 12832
rect 19116 12792 19122 12804
rect 21085 12801 21097 12804
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 21269 12835 21327 12841
rect 21269 12801 21281 12835
rect 21315 12801 21327 12835
rect 22186 12832 22192 12844
rect 22147 12804 22192 12832
rect 21269 12795 21327 12801
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12764 2743 12767
rect 2958 12764 2964 12776
rect 2731 12736 2964 12764
rect 2731 12733 2743 12736
rect 2685 12727 2743 12733
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 3326 12764 3332 12776
rect 3287 12736 3332 12764
rect 3326 12724 3332 12736
rect 3384 12724 3390 12776
rect 8757 12767 8815 12773
rect 8757 12733 8769 12767
rect 8803 12733 8815 12767
rect 10594 12764 10600 12776
rect 10555 12736 10600 12764
rect 8757 12727 8815 12733
rect 1118 12656 1124 12708
rect 1176 12696 1182 12708
rect 2317 12699 2375 12705
rect 2317 12696 2329 12699
rect 1176 12668 2329 12696
rect 1176 12656 1182 12668
rect 2317 12665 2329 12668
rect 2363 12665 2375 12699
rect 2317 12659 2375 12665
rect 2516 12668 4108 12696
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 2516 12637 2544 12668
rect 2501 12631 2559 12637
rect 2501 12597 2513 12631
rect 2547 12597 2559 12631
rect 2501 12591 2559 12597
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 3694 12628 3700 12640
rect 2648 12600 3700 12628
rect 2648 12588 2654 12600
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 3878 12588 3884 12640
rect 3936 12628 3942 12640
rect 3973 12631 4031 12637
rect 3973 12628 3985 12631
rect 3936 12600 3985 12628
rect 3936 12588 3942 12600
rect 3973 12597 3985 12600
rect 4019 12597 4031 12631
rect 4080 12628 4108 12668
rect 7742 12656 7748 12708
rect 7800 12696 7806 12708
rect 8772 12696 8800 12727
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 18095 12736 19104 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 7800 12668 8800 12696
rect 7800 12656 7806 12668
rect 11146 12656 11152 12708
rect 11204 12696 11210 12708
rect 11609 12699 11667 12705
rect 11609 12696 11621 12699
rect 11204 12668 11621 12696
rect 11204 12656 11210 12668
rect 11609 12665 11621 12668
rect 11655 12696 11667 12699
rect 11974 12696 11980 12708
rect 11655 12668 11980 12696
rect 11655 12665 11667 12668
rect 11609 12659 11667 12665
rect 11974 12656 11980 12668
rect 12032 12656 12038 12708
rect 15010 12656 15016 12708
rect 15068 12696 15074 12708
rect 16942 12696 16948 12708
rect 15068 12668 16948 12696
rect 15068 12656 15074 12668
rect 16942 12656 16948 12668
rect 17000 12656 17006 12708
rect 4706 12628 4712 12640
rect 4080 12600 4712 12628
rect 3973 12591 4031 12597
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 5813 12631 5871 12637
rect 5813 12597 5825 12631
rect 5859 12628 5871 12631
rect 5902 12628 5908 12640
rect 5859 12600 5908 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 6730 12628 6736 12640
rect 6420 12600 6736 12628
rect 6420 12588 6426 12600
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 9214 12588 9220 12640
rect 9272 12628 9278 12640
rect 10965 12631 11023 12637
rect 10965 12628 10977 12631
rect 9272 12600 10977 12628
rect 9272 12588 9278 12600
rect 10965 12597 10977 12600
rect 11011 12597 11023 12631
rect 10965 12591 11023 12597
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 13449 12631 13507 12637
rect 13449 12628 13461 12631
rect 11388 12600 13461 12628
rect 11388 12588 11394 12600
rect 13449 12597 13461 12600
rect 13495 12628 13507 12631
rect 14642 12628 14648 12640
rect 13495 12600 14648 12628
rect 13495 12597 13507 12600
rect 13449 12591 13507 12597
rect 14642 12588 14648 12600
rect 14700 12588 14706 12640
rect 16390 12588 16396 12640
rect 16448 12628 16454 12640
rect 16574 12628 16580 12640
rect 16448 12600 16580 12628
rect 16448 12588 16454 12600
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 16666 12588 16672 12640
rect 16724 12628 16730 12640
rect 18064 12628 18092 12727
rect 18322 12656 18328 12708
rect 18380 12696 18386 12708
rect 19076 12696 19104 12736
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 20438 12764 20444 12776
rect 19392 12736 20444 12764
rect 19392 12724 19398 12736
rect 20438 12724 20444 12736
rect 20496 12724 20502 12776
rect 21082 12696 21088 12708
rect 18380 12668 19012 12696
rect 19076 12668 21088 12696
rect 18380 12656 18386 12668
rect 18984 12640 19012 12668
rect 21082 12656 21088 12668
rect 21140 12656 21146 12708
rect 21284 12696 21312 12795
rect 22186 12792 22192 12804
rect 22244 12832 22250 12844
rect 23014 12832 23020 12844
rect 22244 12804 23020 12832
rect 22244 12792 22250 12804
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 23658 12832 23664 12844
rect 23619 12804 23664 12832
rect 23658 12792 23664 12804
rect 23716 12792 23722 12844
rect 23842 12832 23848 12844
rect 23803 12804 23848 12832
rect 23842 12792 23848 12804
rect 23900 12792 23906 12844
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12832 24455 12835
rect 29822 12832 29828 12844
rect 24443 12804 29828 12832
rect 24443 12801 24455 12804
rect 24397 12795 24455 12801
rect 29822 12792 29828 12804
rect 29880 12792 29886 12844
rect 22922 12764 22928 12776
rect 22066 12736 22928 12764
rect 22066 12696 22094 12736
rect 22922 12724 22928 12736
rect 22980 12724 22986 12776
rect 24949 12767 25007 12773
rect 24949 12733 24961 12767
rect 24995 12764 25007 12767
rect 25222 12764 25228 12776
rect 24995 12736 25228 12764
rect 24995 12733 25007 12736
rect 24949 12727 25007 12733
rect 25222 12724 25228 12736
rect 25280 12724 25286 12776
rect 29733 12767 29791 12773
rect 29733 12764 29745 12767
rect 27540 12736 29745 12764
rect 23474 12696 23480 12708
rect 21284 12668 22094 12696
rect 23435 12668 23480 12696
rect 23474 12656 23480 12668
rect 23532 12656 23538 12708
rect 24302 12656 24308 12708
rect 24360 12696 24366 12708
rect 27540 12705 27568 12736
rect 29733 12733 29745 12736
rect 29779 12733 29791 12767
rect 29733 12727 29791 12733
rect 27525 12699 27583 12705
rect 27525 12696 27537 12699
rect 24360 12668 27537 12696
rect 24360 12656 24366 12668
rect 27525 12665 27537 12668
rect 27571 12665 27583 12699
rect 27525 12659 27583 12665
rect 28442 12656 28448 12708
rect 28500 12696 28506 12708
rect 28500 12668 31754 12696
rect 28500 12656 28506 12668
rect 16724 12600 18092 12628
rect 16724 12588 16730 12600
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 18877 12631 18935 12637
rect 18877 12628 18889 12631
rect 18656 12600 18889 12628
rect 18656 12588 18662 12600
rect 18877 12597 18889 12600
rect 18923 12597 18935 12631
rect 18877 12591 18935 12597
rect 18966 12588 18972 12640
rect 19024 12588 19030 12640
rect 19426 12628 19432 12640
rect 19387 12600 19432 12628
rect 19426 12588 19432 12600
rect 19484 12588 19490 12640
rect 19610 12628 19616 12640
rect 19571 12600 19616 12628
rect 19610 12588 19616 12600
rect 19668 12628 19674 12640
rect 20254 12628 20260 12640
rect 19668 12600 20260 12628
rect 19668 12588 19674 12600
rect 20254 12588 20260 12600
rect 20312 12588 20318 12640
rect 20438 12628 20444 12640
rect 20399 12600 20444 12628
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 20625 12631 20683 12637
rect 20625 12597 20637 12631
rect 20671 12628 20683 12631
rect 20714 12628 20720 12640
rect 20671 12600 20720 12628
rect 20671 12597 20683 12600
rect 20625 12591 20683 12597
rect 20714 12588 20720 12600
rect 20772 12628 20778 12640
rect 24854 12628 24860 12640
rect 20772 12600 24860 12628
rect 20772 12588 20778 12600
rect 24854 12588 24860 12600
rect 24912 12588 24918 12640
rect 27062 12628 27068 12640
rect 26975 12600 27068 12628
rect 27062 12588 27068 12600
rect 27120 12628 27126 12640
rect 27246 12628 27252 12640
rect 27120 12600 27252 12628
rect 27120 12588 27126 12600
rect 27246 12588 27252 12600
rect 27304 12588 27310 12640
rect 31726 12628 31754 12668
rect 34606 12628 34612 12640
rect 31726 12600 34612 12628
rect 34606 12588 34612 12600
rect 34664 12588 34670 12640
rect 1104 12538 44896 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 44896 12538
rect 1104 12464 44896 12486
rect 2590 12424 2596 12436
rect 2551 12396 2596 12424
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 5902 12384 5908 12436
rect 5960 12424 5966 12436
rect 6270 12424 6276 12436
rect 5960 12396 6276 12424
rect 5960 12384 5966 12396
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 6420 12396 10456 12424
rect 6420 12384 6426 12396
rect 1854 12356 1860 12368
rect 1815 12328 1860 12356
rect 1854 12316 1860 12328
rect 1912 12316 1918 12368
rect 5258 12356 5264 12368
rect 4724 12328 5264 12356
rect 2498 12288 2504 12300
rect 2459 12260 2504 12288
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 3694 12248 3700 12300
rect 3752 12288 3758 12300
rect 4246 12288 4252 12300
rect 3752 12260 4252 12288
rect 3752 12248 3758 12260
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 4522 12248 4528 12300
rect 4580 12288 4586 12300
rect 4724 12297 4752 12328
rect 5258 12316 5264 12328
rect 5316 12316 5322 12368
rect 5442 12316 5448 12368
rect 5500 12356 5506 12368
rect 7190 12356 7196 12368
rect 5500 12328 7196 12356
rect 5500 12316 5506 12328
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 8110 12356 8116 12368
rect 7524 12328 8116 12356
rect 7524 12316 7530 12328
rect 8110 12316 8116 12328
rect 8168 12316 8174 12368
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 8352 12328 9444 12356
rect 8352 12316 8358 12328
rect 4709 12291 4767 12297
rect 4580 12260 4625 12288
rect 4580 12248 4586 12260
rect 4709 12257 4721 12291
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 4816 12260 5120 12288
rect 1946 12180 1952 12232
rect 2004 12220 2010 12232
rect 2409 12223 2467 12229
rect 2409 12220 2421 12223
rect 2004 12192 2421 12220
rect 2004 12180 2010 12192
rect 2409 12189 2421 12192
rect 2455 12189 2467 12223
rect 2682 12220 2688 12232
rect 2643 12192 2688 12220
rect 2409 12183 2467 12189
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 2866 12180 2872 12232
rect 2924 12220 2930 12232
rect 3418 12220 3424 12232
rect 2924 12192 3424 12220
rect 2924 12180 2930 12192
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3786 12180 3792 12232
rect 3844 12220 3850 12232
rect 4816 12220 4844 12260
rect 3844 12192 4844 12220
rect 5092 12220 5120 12260
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 8938 12288 8944 12300
rect 5592 12260 8432 12288
rect 8899 12260 8944 12288
rect 5592 12248 5598 12260
rect 8404 12232 8432 12260
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 9122 12288 9128 12300
rect 9083 12260 9128 12288
rect 9122 12248 9128 12260
rect 9180 12248 9186 12300
rect 9416 12288 9444 12328
rect 10428 12297 10456 12396
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12710 12424 12716 12436
rect 12584 12396 12716 12424
rect 12584 12384 12590 12396
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 12820 12396 15056 12424
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 11882 12356 11888 12368
rect 11020 12328 11888 12356
rect 11020 12316 11026 12328
rect 11882 12316 11888 12328
rect 11940 12316 11946 12368
rect 12820 12356 12848 12396
rect 12406 12328 12848 12356
rect 15028 12356 15056 12396
rect 15102 12384 15108 12436
rect 15160 12424 15166 12436
rect 15286 12424 15292 12436
rect 15160 12396 15292 12424
rect 15160 12384 15166 12396
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 15473 12427 15531 12433
rect 15473 12393 15485 12427
rect 15519 12424 15531 12427
rect 15654 12424 15660 12436
rect 15519 12396 15660 12424
rect 15519 12393 15531 12396
rect 15473 12387 15531 12393
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 16390 12424 16396 12436
rect 15764 12396 16396 12424
rect 15764 12356 15792 12396
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 16592 12396 17877 12424
rect 16482 12356 16488 12368
rect 15028 12328 15792 12356
rect 16443 12328 16488 12356
rect 10413 12291 10471 12297
rect 9416 12260 10364 12288
rect 5810 12220 5816 12232
rect 5092 12192 5488 12220
rect 5771 12192 5816 12220
rect 3844 12180 3850 12192
rect 5460 12164 5488 12192
rect 5810 12180 5816 12192
rect 5868 12180 5874 12232
rect 6086 12220 6092 12232
rect 6047 12192 6092 12220
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 8444 12192 8489 12220
rect 8444 12180 8450 12192
rect 1489 12155 1547 12161
rect 1489 12121 1501 12155
rect 1535 12152 1547 12155
rect 2498 12152 2504 12164
rect 1535 12124 2504 12152
rect 1535 12121 1547 12124
rect 1489 12115 1547 12121
rect 2498 12112 2504 12124
rect 2556 12112 2562 12164
rect 3878 12112 3884 12164
rect 3936 12152 3942 12164
rect 5074 12152 5080 12164
rect 3936 12124 5080 12152
rect 3936 12112 3942 12124
rect 5074 12112 5080 12124
rect 5132 12112 5138 12164
rect 5442 12112 5448 12164
rect 5500 12152 5506 12164
rect 6549 12155 6607 12161
rect 6549 12152 6561 12155
rect 5500 12124 6561 12152
rect 5500 12112 5506 12124
rect 6549 12121 6561 12124
rect 6595 12121 6607 12155
rect 6549 12115 6607 12121
rect 7466 12112 7472 12164
rect 7524 12152 7530 12164
rect 7742 12152 7748 12164
rect 7524 12124 7748 12152
rect 7524 12112 7530 12124
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 8202 12152 8208 12164
rect 8163 12124 8208 12152
rect 8202 12112 8208 12124
rect 8260 12112 8266 12164
rect 9306 12152 9312 12164
rect 8312 12124 9312 12152
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 2314 12044 2320 12096
rect 2372 12084 2378 12096
rect 2774 12084 2780 12096
rect 2372 12056 2780 12084
rect 2372 12044 2378 12056
rect 2774 12044 2780 12056
rect 2832 12084 2838 12096
rect 2869 12087 2927 12093
rect 2869 12084 2881 12087
rect 2832 12056 2881 12084
rect 2832 12044 2838 12056
rect 2869 12053 2881 12056
rect 2915 12084 2927 12087
rect 3050 12084 3056 12096
rect 2915 12056 3056 12084
rect 2915 12053 2927 12056
rect 2869 12047 2927 12053
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 4062 12084 4068 12096
rect 4023 12056 4068 12084
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 4433 12087 4491 12093
rect 4433 12053 4445 12087
rect 4479 12084 4491 12087
rect 4890 12084 4896 12096
rect 4479 12056 4896 12084
rect 4479 12053 4491 12056
rect 4433 12047 4491 12053
rect 4890 12044 4896 12056
rect 4948 12084 4954 12096
rect 8312 12084 8340 12124
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 10336 12152 10364 12260
rect 10413 12257 10425 12291
rect 10459 12257 10471 12291
rect 11241 12291 11299 12297
rect 11241 12288 11253 12291
rect 10413 12251 10471 12257
rect 10888 12260 11253 12288
rect 10888 12152 10916 12260
rect 11241 12257 11253 12260
rect 11287 12288 11299 12291
rect 12406 12288 12434 12328
rect 16482 12316 16488 12328
rect 16540 12316 16546 12368
rect 12710 12288 12716 12300
rect 11287 12260 12434 12288
rect 12671 12260 12716 12288
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 15102 12248 15108 12300
rect 15160 12288 15166 12300
rect 16592 12288 16620 12396
rect 17865 12393 17877 12396
rect 17911 12393 17923 12427
rect 18690 12424 18696 12436
rect 17865 12387 17923 12393
rect 17972 12396 18696 12424
rect 17310 12356 17316 12368
rect 17271 12328 17316 12356
rect 17310 12316 17316 12328
rect 17368 12316 17374 12368
rect 15160 12260 16620 12288
rect 15160 12248 15166 12260
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 17972 12288 18000 12396
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 19058 12384 19064 12436
rect 19116 12424 19122 12436
rect 19426 12424 19432 12436
rect 19116 12396 19432 12424
rect 19116 12384 19122 12396
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 19518 12384 19524 12436
rect 19576 12424 19582 12436
rect 21545 12427 21603 12433
rect 21545 12424 21557 12427
rect 19576 12396 21557 12424
rect 19576 12384 19582 12396
rect 21545 12393 21557 12396
rect 21591 12393 21603 12427
rect 24118 12424 24124 12436
rect 21545 12387 21603 12393
rect 21652 12396 24124 12424
rect 18046 12316 18052 12368
rect 18104 12356 18110 12368
rect 20257 12359 20315 12365
rect 18104 12328 20116 12356
rect 18104 12316 18110 12328
rect 16724 12260 18000 12288
rect 18233 12291 18291 12297
rect 16724 12248 16730 12260
rect 18233 12257 18245 12291
rect 18279 12288 18291 12291
rect 19334 12288 19340 12300
rect 18279 12260 19340 12288
rect 18279 12257 18291 12260
rect 18233 12251 18291 12257
rect 19334 12248 19340 12260
rect 19392 12248 19398 12300
rect 19613 12291 19671 12297
rect 19613 12257 19625 12291
rect 19659 12288 19671 12291
rect 19702 12288 19708 12300
rect 19659 12260 19708 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12220 14151 12223
rect 14826 12220 14832 12232
rect 14139 12192 14832 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 16114 12220 16120 12232
rect 16075 12192 16120 12220
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 16298 12220 16304 12232
rect 16259 12192 16304 12220
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 17129 12223 17187 12229
rect 17129 12189 17141 12223
rect 17175 12220 17187 12223
rect 17310 12220 17316 12232
rect 17175 12192 17316 12220
rect 17175 12189 17187 12192
rect 17129 12183 17187 12189
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12220 17463 12223
rect 17494 12220 17500 12232
rect 17451 12192 17500 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 17586 12180 17592 12232
rect 17644 12220 17650 12232
rect 18049 12223 18107 12229
rect 18049 12220 18061 12223
rect 17644 12192 18061 12220
rect 17644 12180 17650 12192
rect 18049 12189 18061 12192
rect 18095 12189 18107 12223
rect 18322 12220 18328 12232
rect 18283 12192 18328 12220
rect 18049 12183 18107 12189
rect 18322 12180 18328 12192
rect 18380 12220 18386 12232
rect 19150 12220 19156 12232
rect 18380 12192 19156 12220
rect 18380 12180 18386 12192
rect 19150 12180 19156 12192
rect 19208 12180 19214 12232
rect 19426 12220 19432 12232
rect 19387 12192 19432 12220
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 20088 12229 20116 12328
rect 20257 12325 20269 12359
rect 20303 12356 20315 12359
rect 20346 12356 20352 12368
rect 20303 12328 20352 12356
rect 20303 12325 20315 12328
rect 20257 12319 20315 12325
rect 20346 12316 20352 12328
rect 20404 12316 20410 12368
rect 20898 12316 20904 12368
rect 20956 12356 20962 12368
rect 20993 12359 21051 12365
rect 20993 12356 21005 12359
rect 20956 12328 21005 12356
rect 20956 12316 20962 12328
rect 20993 12325 21005 12328
rect 21039 12356 21051 12359
rect 21652 12356 21680 12396
rect 24118 12384 24124 12396
rect 24176 12384 24182 12436
rect 25593 12427 25651 12433
rect 25593 12393 25605 12427
rect 25639 12424 25651 12427
rect 25682 12424 25688 12436
rect 25639 12396 25688 12424
rect 25639 12393 25651 12396
rect 25593 12387 25651 12393
rect 25682 12384 25688 12396
rect 25740 12384 25746 12436
rect 26142 12424 26148 12436
rect 26103 12396 26148 12424
rect 26142 12384 26148 12396
rect 26200 12384 26206 12436
rect 26970 12384 26976 12436
rect 27028 12424 27034 12436
rect 28261 12427 28319 12433
rect 28261 12424 28273 12427
rect 27028 12396 28273 12424
rect 27028 12384 27034 12396
rect 28261 12393 28273 12396
rect 28307 12393 28319 12427
rect 28261 12387 28319 12393
rect 21039 12328 21680 12356
rect 21039 12325 21051 12328
rect 20993 12319 21051 12325
rect 21726 12316 21732 12368
rect 21784 12356 21790 12368
rect 27801 12359 27859 12365
rect 21784 12328 23428 12356
rect 21784 12316 21790 12328
rect 20824 12260 23336 12288
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20438 12180 20444 12232
rect 20496 12220 20502 12232
rect 20824 12229 20852 12260
rect 20809 12223 20867 12229
rect 20496 12192 20668 12220
rect 20496 12180 20502 12192
rect 10336 12124 10916 12152
rect 11146 12112 11152 12164
rect 11204 12152 11210 12164
rect 11425 12155 11483 12161
rect 11425 12152 11437 12155
rect 11204 12124 11437 12152
rect 11204 12112 11210 12124
rect 11425 12121 11437 12124
rect 11471 12121 11483 12155
rect 11425 12115 11483 12121
rect 14360 12155 14418 12161
rect 14360 12121 14372 12155
rect 14406 12152 14418 12155
rect 16666 12152 16672 12164
rect 14406 12124 16672 12152
rect 14406 12121 14418 12124
rect 14360 12115 14418 12121
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 16942 12152 16948 12164
rect 16903 12124 16948 12152
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 19242 12152 19248 12164
rect 17052 12124 17954 12152
rect 19203 12124 19248 12152
rect 4948 12056 8340 12084
rect 4948 12044 4954 12056
rect 9030 12044 9036 12096
rect 9088 12084 9094 12096
rect 15102 12084 15108 12096
rect 9088 12056 15108 12084
rect 9088 12044 9094 12056
rect 15102 12044 15108 12056
rect 15160 12044 15166 12096
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 15654 12084 15660 12096
rect 15344 12056 15660 12084
rect 15344 12044 15350 12056
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 15933 12087 15991 12093
rect 15933 12053 15945 12087
rect 15979 12084 15991 12087
rect 16114 12084 16120 12096
rect 15979 12056 16120 12084
rect 15979 12053 15991 12056
rect 15933 12047 15991 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16209 12087 16267 12093
rect 16209 12053 16221 12087
rect 16255 12084 16267 12087
rect 16390 12084 16396 12096
rect 16255 12056 16396 12084
rect 16255 12053 16267 12056
rect 16209 12047 16267 12053
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 16482 12044 16488 12096
rect 16540 12084 16546 12096
rect 17052 12084 17080 12124
rect 16540 12056 17080 12084
rect 16540 12044 16546 12056
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 17586 12084 17592 12096
rect 17368 12056 17592 12084
rect 17368 12044 17374 12056
rect 17586 12044 17592 12056
rect 17644 12044 17650 12096
rect 17926 12084 17954 12124
rect 19242 12112 19248 12124
rect 19300 12112 19306 12164
rect 19334 12112 19340 12164
rect 19392 12152 19398 12164
rect 20640 12152 20668 12192
rect 20809 12189 20821 12223
rect 20855 12189 20867 12223
rect 21545 12223 21603 12229
rect 21545 12220 21557 12223
rect 20809 12183 20867 12189
rect 21100 12192 21557 12220
rect 21100 12152 21128 12192
rect 21545 12189 21557 12192
rect 21591 12189 21603 12223
rect 21545 12183 21603 12189
rect 21726 12180 21732 12232
rect 21784 12220 21790 12232
rect 21784 12192 21877 12220
rect 21784 12180 21790 12192
rect 22462 12180 22468 12232
rect 22520 12220 22526 12232
rect 22557 12223 22615 12229
rect 22557 12220 22569 12223
rect 22520 12192 22569 12220
rect 22520 12180 22526 12192
rect 22557 12189 22569 12192
rect 22603 12189 22615 12223
rect 23198 12220 23204 12232
rect 23159 12192 23204 12220
rect 22557 12183 22615 12189
rect 23198 12180 23204 12192
rect 23256 12180 23262 12232
rect 19392 12124 20576 12152
rect 20640 12124 21128 12152
rect 19392 12112 19398 12124
rect 20438 12084 20444 12096
rect 17926 12056 20444 12084
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 20548 12084 20576 12124
rect 21174 12112 21180 12164
rect 21232 12152 21238 12164
rect 21744 12152 21772 12180
rect 23216 12152 23244 12180
rect 21232 12124 21772 12152
rect 22756 12124 23244 12152
rect 23308 12152 23336 12260
rect 23400 12229 23428 12328
rect 27801 12325 27813 12359
rect 27847 12356 27859 12359
rect 28534 12356 28540 12368
rect 27847 12328 28540 12356
rect 27847 12325 27859 12328
rect 27801 12319 27859 12325
rect 28534 12316 28540 12328
rect 28592 12316 28598 12368
rect 25222 12248 25228 12300
rect 25280 12288 25286 12300
rect 27982 12288 27988 12300
rect 25280 12260 27988 12288
rect 25280 12248 25286 12260
rect 27982 12248 27988 12260
rect 28040 12248 28046 12300
rect 29546 12288 29552 12300
rect 29507 12260 29552 12288
rect 29546 12248 29552 12260
rect 29604 12248 29610 12300
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12220 23443 12223
rect 27798 12220 27804 12232
rect 23431 12192 27804 12220
rect 23431 12189 23443 12192
rect 23385 12183 23443 12189
rect 27798 12180 27804 12192
rect 27856 12220 27862 12232
rect 28813 12223 28871 12229
rect 28813 12220 28825 12223
rect 27856 12192 28825 12220
rect 27856 12180 27862 12192
rect 28813 12189 28825 12192
rect 28859 12189 28871 12223
rect 28813 12183 28871 12189
rect 24394 12152 24400 12164
rect 23308 12124 24400 12152
rect 21232 12112 21238 12124
rect 22756 12093 22784 12124
rect 24394 12112 24400 12124
rect 24452 12112 24458 12164
rect 24486 12112 24492 12164
rect 24544 12152 24550 12164
rect 25041 12155 25099 12161
rect 25041 12152 25053 12155
rect 24544 12124 25053 12152
rect 24544 12112 24550 12124
rect 25041 12121 25053 12124
rect 25087 12152 25099 12155
rect 30101 12155 30159 12161
rect 30101 12152 30113 12155
rect 25087 12124 30113 12152
rect 25087 12121 25099 12124
rect 25041 12115 25099 12121
rect 30101 12121 30113 12124
rect 30147 12121 30159 12155
rect 30101 12115 30159 12121
rect 22741 12087 22799 12093
rect 22741 12084 22753 12087
rect 20548 12056 22753 12084
rect 22741 12053 22753 12056
rect 22787 12053 22799 12087
rect 23290 12084 23296 12096
rect 23251 12056 23296 12084
rect 22741 12047 22799 12053
rect 23290 12044 23296 12056
rect 23348 12044 23354 12096
rect 23382 12044 23388 12096
rect 23440 12084 23446 12096
rect 26605 12087 26663 12093
rect 26605 12084 26617 12087
rect 23440 12056 26617 12084
rect 23440 12044 23446 12056
rect 26605 12053 26617 12056
rect 26651 12084 26663 12087
rect 26694 12084 26700 12096
rect 26651 12056 26700 12084
rect 26651 12053 26663 12056
rect 26605 12047 26663 12053
rect 26694 12044 26700 12056
rect 26752 12044 26758 12096
rect 27249 12087 27307 12093
rect 27249 12053 27261 12087
rect 27295 12084 27307 12087
rect 27430 12084 27436 12096
rect 27295 12056 27436 12084
rect 27295 12053 27307 12056
rect 27249 12047 27307 12053
rect 27430 12044 27436 12056
rect 27488 12044 27494 12096
rect 1104 11994 44896 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 44896 11994
rect 1104 11920 44896 11942
rect 1854 11840 1860 11892
rect 1912 11880 1918 11892
rect 3602 11880 3608 11892
rect 1912 11852 3608 11880
rect 1912 11840 1918 11852
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 3697 11883 3755 11889
rect 3697 11849 3709 11883
rect 3743 11880 3755 11883
rect 3970 11880 3976 11892
rect 3743 11852 3976 11880
rect 3743 11849 3755 11852
rect 3697 11843 3755 11849
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 4154 11880 4160 11892
rect 4080 11852 4160 11880
rect 1302 11772 1308 11824
rect 1360 11812 1366 11824
rect 1673 11815 1731 11821
rect 1673 11812 1685 11815
rect 1360 11784 1685 11812
rect 1360 11772 1366 11784
rect 1673 11781 1685 11784
rect 1719 11781 1731 11815
rect 1673 11775 1731 11781
rect 2958 11704 2964 11756
rect 3016 11744 3022 11756
rect 3237 11747 3295 11753
rect 3237 11744 3249 11747
rect 3016 11716 3249 11744
rect 3016 11704 3022 11716
rect 3237 11713 3249 11716
rect 3283 11713 3295 11747
rect 3418 11744 3424 11756
rect 3379 11716 3424 11744
rect 3237 11707 3295 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 3510 11704 3516 11756
rect 3568 11744 3574 11756
rect 3878 11744 3884 11756
rect 3568 11716 3884 11744
rect 3568 11704 3574 11716
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 3970 11704 3976 11756
rect 4028 11744 4034 11756
rect 4080 11744 4108 11852
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5353 11883 5411 11889
rect 5353 11849 5365 11883
rect 5399 11880 5411 11883
rect 5718 11880 5724 11892
rect 5399 11852 5724 11880
rect 5399 11849 5411 11852
rect 5353 11843 5411 11849
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 8110 11840 8116 11892
rect 8168 11840 8174 11892
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 12894 11880 12900 11892
rect 8444 11852 12900 11880
rect 8444 11840 8450 11852
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 13354 11880 13360 11892
rect 13315 11852 13360 11880
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 15286 11880 15292 11892
rect 14384 11852 15292 11880
rect 6178 11812 6184 11824
rect 4816 11784 6184 11812
rect 4157 11747 4215 11753
rect 4157 11744 4169 11747
rect 4028 11716 4169 11744
rect 4028 11704 4034 11716
rect 4157 11713 4169 11716
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 4246 11704 4252 11756
rect 4304 11744 4310 11756
rect 4426 11747 4484 11753
rect 4426 11744 4438 11747
rect 4304 11716 4438 11744
rect 4304 11704 4310 11716
rect 4426 11713 4438 11716
rect 4472 11713 4484 11747
rect 4426 11707 4484 11713
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 4816 11744 4844 11784
rect 6178 11772 6184 11784
rect 6236 11772 6242 11824
rect 7742 11812 7748 11824
rect 6472 11784 7748 11812
rect 4764 11716 4844 11744
rect 4764 11704 4770 11716
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11676 2375 11679
rect 2498 11676 2504 11688
rect 2363 11648 2504 11676
rect 2363 11645 2375 11648
rect 2317 11639 2375 11645
rect 2498 11636 2504 11648
rect 2556 11636 2562 11688
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 2866 11676 2872 11688
rect 2823 11648 2872 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 4341 11679 4399 11685
rect 4341 11645 4353 11679
rect 4387 11645 4399 11679
rect 4341 11639 4399 11645
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11608 1915 11611
rect 2222 11608 2228 11620
rect 1903 11580 2228 11608
rect 1903 11577 1915 11580
rect 1857 11571 1915 11577
rect 2222 11568 2228 11580
rect 2280 11568 2286 11620
rect 2685 11611 2743 11617
rect 2685 11577 2697 11611
rect 2731 11608 2743 11611
rect 4062 11608 4068 11620
rect 2731 11580 4068 11608
rect 2731 11577 2743 11580
rect 2685 11571 2743 11577
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 3050 11540 3056 11552
rect 1636 11512 3056 11540
rect 1636 11500 1642 11512
rect 3050 11500 3056 11512
rect 3108 11540 3114 11552
rect 3237 11543 3295 11549
rect 3237 11540 3249 11543
rect 3108 11512 3249 11540
rect 3108 11500 3114 11512
rect 3237 11509 3249 11512
rect 3283 11509 3295 11543
rect 3237 11503 3295 11509
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 4356 11540 4384 11639
rect 4816 11608 4844 11716
rect 5445 11747 5503 11753
rect 5445 11713 5457 11747
rect 5491 11744 5503 11747
rect 6362 11744 6368 11756
rect 5491 11716 6368 11744
rect 5491 11713 5503 11716
rect 5445 11707 5503 11713
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 5258 11676 5264 11688
rect 5171 11648 5264 11676
rect 5258 11636 5264 11648
rect 5316 11676 5322 11688
rect 6472 11676 6500 11784
rect 7742 11772 7748 11784
rect 7800 11772 7806 11824
rect 8128 11812 8156 11840
rect 10318 11812 10324 11824
rect 8128 11784 9168 11812
rect 10279 11784 10324 11812
rect 7092 11747 7150 11753
rect 7092 11713 7104 11747
rect 7138 11744 7150 11747
rect 7138 11716 8892 11744
rect 7138 11713 7150 11716
rect 7092 11707 7150 11713
rect 8864 11688 8892 11716
rect 6822 11676 6828 11688
rect 5316 11648 6500 11676
rect 6783 11648 6828 11676
rect 5316 11636 5322 11648
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 8846 11636 8852 11688
rect 8904 11636 8910 11688
rect 9030 11676 9036 11688
rect 8991 11648 9036 11676
rect 9030 11636 9036 11648
rect 9088 11636 9094 11688
rect 9140 11676 9168 11784
rect 10318 11772 10324 11784
rect 10376 11772 10382 11824
rect 11790 11821 11796 11824
rect 11784 11812 11796 11821
rect 11751 11784 11796 11812
rect 11784 11775 11796 11784
rect 11790 11772 11796 11775
rect 11848 11772 11854 11824
rect 14384 11812 14412 11852
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 15746 11880 15752 11892
rect 15707 11852 15752 11880
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 16298 11840 16304 11892
rect 16356 11880 16362 11892
rect 17494 11880 17500 11892
rect 16356 11852 17500 11880
rect 16356 11840 16362 11852
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 18509 11883 18567 11889
rect 18509 11849 18521 11883
rect 18555 11880 18567 11883
rect 18598 11880 18604 11892
rect 18555 11852 18604 11880
rect 18555 11849 18567 11852
rect 18509 11843 18567 11849
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 20254 11840 20260 11892
rect 20312 11880 20318 11892
rect 20312 11852 20357 11880
rect 20312 11840 20318 11852
rect 20714 11840 20720 11892
rect 20772 11840 20778 11892
rect 21818 11880 21824 11892
rect 21779 11852 21824 11880
rect 21818 11840 21824 11852
rect 21876 11840 21882 11892
rect 22646 11880 22652 11892
rect 22607 11852 22652 11880
rect 22646 11840 22652 11852
rect 22704 11840 22710 11892
rect 23474 11840 23480 11892
rect 23532 11880 23538 11892
rect 24118 11880 24124 11892
rect 23532 11852 24124 11880
rect 23532 11840 23538 11852
rect 24118 11840 24124 11852
rect 24176 11840 24182 11892
rect 25314 11840 25320 11892
rect 25372 11880 25378 11892
rect 27522 11880 27528 11892
rect 25372 11852 27528 11880
rect 25372 11840 25378 11852
rect 27522 11840 27528 11852
rect 27580 11840 27586 11892
rect 27798 11840 27804 11892
rect 27856 11880 27862 11892
rect 28077 11883 28135 11889
rect 28077 11880 28089 11883
rect 27856 11852 28089 11880
rect 27856 11840 27862 11852
rect 28077 11849 28089 11852
rect 28123 11849 28135 11883
rect 28626 11880 28632 11892
rect 28587 11852 28632 11880
rect 28077 11843 28135 11849
rect 28626 11840 28632 11852
rect 28684 11840 28690 11892
rect 12176 11784 14412 11812
rect 14492 11815 14550 11821
rect 12176 11756 12204 11784
rect 14492 11781 14504 11815
rect 14538 11812 14550 11815
rect 15010 11812 15016 11824
rect 14538 11784 15016 11812
rect 14538 11781 14550 11784
rect 14492 11775 14550 11781
rect 15010 11772 15016 11784
rect 15068 11772 15074 11824
rect 15470 11812 15476 11824
rect 15431 11784 15476 11812
rect 15470 11772 15476 11784
rect 15528 11772 15534 11824
rect 15930 11772 15936 11824
rect 15988 11812 15994 11824
rect 15988 11784 17724 11812
rect 15988 11772 15994 11784
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 12158 11744 12164 11756
rect 10560 11716 10605 11744
rect 11164 11716 12164 11744
rect 10560 11704 10566 11716
rect 9140 11648 9996 11676
rect 4448 11580 4844 11608
rect 4448 11549 4476 11580
rect 4982 11568 4988 11620
rect 5040 11608 5046 11620
rect 6454 11608 6460 11620
rect 5040 11580 6460 11608
rect 5040 11568 5046 11580
rect 6454 11568 6460 11580
rect 6512 11568 6518 11620
rect 8205 11611 8263 11617
rect 8205 11577 8217 11611
rect 8251 11608 8263 11611
rect 8386 11608 8392 11620
rect 8251 11580 8392 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 8386 11568 8392 11580
rect 8444 11608 8450 11620
rect 9968 11608 9996 11648
rect 11164 11608 11192 11716
rect 12158 11704 12164 11716
rect 12216 11704 12222 11756
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 13280 11716 15393 11744
rect 13280 11688 13308 11716
rect 15381 11713 15393 11716
rect 15427 11713 15439 11747
rect 15562 11744 15568 11756
rect 15523 11716 15568 11744
rect 15381 11707 15439 11713
rect 11238 11636 11244 11688
rect 11296 11676 11302 11688
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11296 11648 11529 11676
rect 11296 11636 11302 11648
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 13262 11636 13268 11688
rect 13320 11636 13326 11688
rect 14734 11676 14740 11688
rect 14695 11648 14740 11676
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 15197 11679 15255 11685
rect 15197 11645 15209 11679
rect 15243 11676 15255 11679
rect 15286 11676 15292 11688
rect 15243 11648 15292 11676
rect 15243 11645 15255 11648
rect 15197 11639 15255 11645
rect 15286 11636 15292 11648
rect 15344 11636 15350 11688
rect 15396 11676 15424 11707
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 15746 11704 15752 11756
rect 15804 11744 15810 11756
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 15804 11716 16681 11744
rect 15804 11704 15810 11716
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 16669 11707 16727 11713
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11744 16911 11747
rect 16899 11716 16988 11744
rect 16899 11713 16911 11716
rect 16853 11707 16911 11713
rect 16022 11676 16028 11688
rect 15396 11648 16028 11676
rect 16022 11636 16028 11648
rect 16080 11636 16086 11688
rect 8444 11580 9904 11608
rect 9968 11580 11192 11608
rect 12897 11611 12955 11617
rect 8444 11568 8450 11580
rect 4028 11512 4384 11540
rect 4433 11543 4491 11549
rect 4028 11500 4034 11512
rect 4433 11509 4445 11543
rect 4479 11509 4491 11543
rect 4433 11503 4491 11509
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11540 4675 11543
rect 5626 11540 5632 11552
rect 4663 11512 5632 11540
rect 4663 11509 4675 11512
rect 4617 11503 4675 11509
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 5813 11543 5871 11549
rect 5813 11509 5825 11543
rect 5859 11540 5871 11543
rect 7098 11540 7104 11552
rect 5859 11512 7104 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 7098 11500 7104 11512
rect 7156 11500 7162 11552
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 9766 11540 9772 11552
rect 7616 11512 9772 11540
rect 7616 11500 7622 11512
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 9876 11540 9904 11580
rect 12897 11577 12909 11611
rect 12943 11608 12955 11611
rect 13446 11608 13452 11620
rect 12943 11580 13452 11608
rect 12943 11577 12955 11580
rect 12897 11571 12955 11577
rect 13446 11568 13452 11580
rect 13504 11568 13510 11620
rect 10502 11540 10508 11552
rect 9876 11512 10508 11540
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 11514 11500 11520 11552
rect 11572 11540 11578 11552
rect 13998 11540 14004 11552
rect 11572 11512 14004 11540
rect 11572 11500 11578 11512
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 16960 11540 16988 11716
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17589 11747 17647 11753
rect 17589 11744 17601 11747
rect 17092 11716 17601 11744
rect 17092 11704 17098 11716
rect 17589 11713 17601 11716
rect 17635 11713 17647 11747
rect 17696 11744 17724 11784
rect 19334 11772 19340 11824
rect 19392 11812 19398 11824
rect 19489 11815 19547 11821
rect 19489 11812 19501 11815
rect 19392 11784 19501 11812
rect 19392 11772 19398 11784
rect 19489 11781 19501 11784
rect 19535 11781 19547 11815
rect 19702 11812 19708 11824
rect 19663 11784 19708 11812
rect 19489 11775 19547 11781
rect 19702 11772 19708 11784
rect 19760 11772 19766 11824
rect 20732 11812 20760 11840
rect 19812 11784 20760 11812
rect 18693 11747 18751 11753
rect 18693 11744 18705 11747
rect 17696 11716 18705 11744
rect 17589 11707 17647 11713
rect 18693 11713 18705 11716
rect 18739 11713 18751 11747
rect 18693 11707 18751 11713
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11744 18935 11747
rect 18966 11744 18972 11756
rect 18923 11716 18972 11744
rect 18923 11713 18935 11716
rect 18877 11707 18935 11713
rect 18966 11704 18972 11716
rect 19024 11704 19030 11756
rect 19812 11744 19840 11784
rect 21542 11772 21548 11824
rect 21600 11812 21606 11824
rect 22002 11812 22008 11824
rect 21600 11784 22008 11812
rect 21600 11772 21606 11784
rect 22002 11772 22008 11784
rect 22060 11772 22066 11824
rect 22094 11772 22100 11824
rect 22152 11812 22158 11824
rect 22833 11815 22891 11821
rect 22833 11812 22845 11815
rect 22152 11784 22845 11812
rect 22152 11772 22158 11784
rect 22833 11781 22845 11784
rect 22879 11812 22891 11815
rect 24029 11815 24087 11821
rect 24029 11812 24041 11815
rect 22879 11784 24041 11812
rect 22879 11781 22891 11784
rect 22833 11775 22891 11781
rect 24029 11781 24041 11784
rect 24075 11781 24087 11815
rect 24136 11812 24164 11840
rect 25685 11815 25743 11821
rect 25685 11812 25697 11815
rect 24136 11784 25697 11812
rect 24029 11775 24087 11781
rect 25685 11781 25697 11784
rect 25731 11781 25743 11815
rect 25685 11775 25743 11781
rect 26329 11815 26387 11821
rect 26329 11781 26341 11815
rect 26375 11812 26387 11815
rect 27614 11812 27620 11824
rect 26375 11784 27620 11812
rect 26375 11781 26387 11784
rect 26329 11775 26387 11781
rect 27614 11772 27620 11784
rect 27672 11772 27678 11824
rect 19076 11716 19840 11744
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 17494 11676 17500 11688
rect 17175 11648 17500 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 19076 11676 19104 11716
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 20162 11744 20168 11756
rect 19944 11716 20168 11744
rect 19944 11704 19950 11716
rect 20162 11704 20168 11716
rect 20220 11704 20226 11756
rect 20349 11747 20407 11753
rect 20349 11713 20361 11747
rect 20395 11744 20407 11747
rect 20714 11744 20720 11756
rect 20395 11716 20720 11744
rect 20395 11713 20407 11716
rect 20349 11707 20407 11713
rect 20714 11704 20720 11716
rect 20772 11704 20778 11756
rect 20990 11744 20996 11756
rect 20951 11716 20996 11744
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 21177 11747 21235 11753
rect 21177 11713 21189 11747
rect 21223 11744 21235 11747
rect 21818 11744 21824 11756
rect 21223 11716 21824 11744
rect 21223 11713 21235 11716
rect 21177 11707 21235 11713
rect 21818 11704 21824 11716
rect 21876 11704 21882 11756
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11713 22247 11747
rect 22189 11707 22247 11713
rect 23017 11747 23075 11753
rect 23017 11713 23029 11747
rect 23063 11744 23075 11747
rect 24486 11744 24492 11756
rect 23063 11716 24492 11744
rect 23063 11713 23075 11716
rect 23017 11707 23075 11713
rect 17696 11648 19104 11676
rect 17037 11611 17095 11617
rect 17037 11577 17049 11611
rect 17083 11608 17095 11611
rect 17696 11608 17724 11648
rect 19150 11636 19156 11688
rect 19208 11676 19214 11688
rect 19702 11676 19708 11688
rect 19208 11648 19708 11676
rect 19208 11636 19214 11648
rect 19702 11636 19708 11648
rect 19760 11636 19766 11688
rect 20530 11676 20536 11688
rect 20088 11648 20536 11676
rect 17083 11580 17724 11608
rect 17083 11577 17095 11580
rect 17037 11571 17095 11577
rect 17770 11568 17776 11620
rect 17828 11608 17834 11620
rect 17865 11611 17923 11617
rect 17865 11608 17877 11611
rect 17828 11580 17877 11608
rect 17828 11568 17834 11580
rect 17865 11577 17877 11580
rect 17911 11577 17923 11611
rect 17865 11571 17923 11577
rect 19337 11611 19395 11617
rect 19337 11577 19349 11611
rect 19383 11608 19395 11611
rect 20088 11608 20116 11648
rect 20530 11636 20536 11648
rect 20588 11636 20594 11688
rect 20732 11676 20760 11704
rect 21910 11676 21916 11688
rect 20732 11648 21916 11676
rect 21910 11636 21916 11648
rect 21968 11636 21974 11688
rect 22204 11676 22232 11707
rect 24486 11704 24492 11716
rect 24544 11704 24550 11756
rect 27982 11704 27988 11756
rect 28040 11744 28046 11756
rect 29733 11747 29791 11753
rect 29733 11744 29745 11747
rect 28040 11716 29745 11744
rect 28040 11704 28046 11716
rect 29733 11713 29745 11716
rect 29779 11713 29791 11747
rect 29733 11707 29791 11713
rect 22204 11648 23612 11676
rect 20806 11608 20812 11620
rect 19383 11580 20116 11608
rect 20767 11580 20812 11608
rect 19383 11577 19395 11580
rect 19337 11571 19395 11577
rect 20806 11568 20812 11580
rect 20864 11568 20870 11620
rect 20990 11568 20996 11620
rect 21048 11608 21054 11620
rect 21726 11608 21732 11620
rect 21048 11580 21732 11608
rect 21048 11568 21054 11580
rect 21726 11568 21732 11580
rect 21784 11608 21790 11620
rect 22830 11608 22836 11620
rect 21784 11580 22836 11608
rect 21784 11568 21790 11580
rect 22830 11568 22836 11580
rect 22888 11568 22894 11620
rect 23584 11552 23612 11648
rect 28626 11636 28632 11688
rect 28684 11676 28690 11688
rect 29181 11679 29239 11685
rect 29181 11676 29193 11679
rect 28684 11648 29193 11676
rect 28684 11636 28690 11648
rect 29181 11645 29193 11648
rect 29227 11645 29239 11679
rect 29181 11639 29239 11645
rect 23658 11568 23664 11620
rect 23716 11608 23722 11620
rect 31294 11608 31300 11620
rect 23716 11580 31300 11608
rect 23716 11568 23722 11580
rect 31294 11568 31300 11580
rect 31352 11568 31358 11620
rect 17494 11540 17500 11552
rect 16960 11512 17500 11540
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 18049 11543 18107 11549
rect 18049 11509 18061 11543
rect 18095 11540 18107 11543
rect 18782 11540 18788 11552
rect 18095 11512 18788 11540
rect 18095 11509 18107 11512
rect 18049 11503 18107 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 19521 11543 19579 11549
rect 19521 11509 19533 11543
rect 19567 11540 19579 11543
rect 19610 11540 19616 11552
rect 19567 11512 19616 11540
rect 19567 11509 19579 11512
rect 19521 11503 19579 11509
rect 19610 11500 19616 11512
rect 19668 11500 19674 11552
rect 19702 11500 19708 11552
rect 19760 11540 19766 11552
rect 20070 11540 20076 11552
rect 19760 11512 20076 11540
rect 19760 11500 19766 11512
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 23566 11540 23572 11552
rect 23527 11512 23572 11540
rect 23566 11500 23572 11512
rect 23624 11500 23630 11552
rect 24486 11500 24492 11552
rect 24544 11540 24550 11552
rect 24581 11543 24639 11549
rect 24581 11540 24593 11543
rect 24544 11512 24593 11540
rect 24544 11500 24550 11512
rect 24581 11509 24593 11512
rect 24627 11509 24639 11543
rect 25222 11540 25228 11552
rect 25183 11512 25228 11540
rect 24581 11503 24639 11509
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 26970 11540 26976 11552
rect 26931 11512 26976 11540
rect 26970 11500 26976 11512
rect 27028 11500 27034 11552
rect 1104 11450 44896 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 44896 11450
rect 1104 11376 44896 11398
rect 1486 11296 1492 11348
rect 1544 11336 1550 11348
rect 1673 11339 1731 11345
rect 1673 11336 1685 11339
rect 1544 11308 1685 11336
rect 1544 11296 1550 11308
rect 1673 11305 1685 11308
rect 1719 11336 1731 11339
rect 2958 11336 2964 11348
rect 1719 11308 2964 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 3418 11336 3424 11348
rect 3068 11308 3424 11336
rect 2866 11228 2872 11280
rect 2924 11268 2930 11280
rect 3068 11268 3096 11308
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 5166 11336 5172 11348
rect 4663 11308 5172 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 6638 11296 6644 11348
rect 6696 11336 6702 11348
rect 12618 11336 12624 11348
rect 6696 11308 12434 11336
rect 12579 11308 12624 11336
rect 6696 11296 6702 11308
rect 2924 11240 3096 11268
rect 3145 11271 3203 11277
rect 2924 11228 2930 11240
rect 3145 11237 3157 11271
rect 3191 11268 3203 11271
rect 5077 11271 5135 11277
rect 5077 11268 5089 11271
rect 3191 11240 5089 11268
rect 3191 11237 3203 11240
rect 3145 11231 3203 11237
rect 5077 11237 5089 11240
rect 5123 11237 5135 11271
rect 5077 11231 5135 11237
rect 5810 11228 5816 11280
rect 5868 11268 5874 11280
rect 5868 11240 9168 11268
rect 5868 11228 5874 11240
rect 3237 11203 3295 11209
rect 3237 11169 3249 11203
rect 3283 11200 3295 11203
rect 4246 11200 4252 11212
rect 3283 11172 4252 11200
rect 3283 11169 3295 11172
rect 3237 11163 3295 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 5534 11200 5540 11212
rect 4356 11172 5304 11200
rect 5495 11172 5540 11200
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 2314 11132 2320 11144
rect 1903 11104 2320 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 3142 11092 3148 11144
rect 3200 11132 3206 11144
rect 3418 11132 3424 11144
rect 3200 11104 3424 11132
rect 3200 11092 3206 11104
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 4356 11141 4384 11172
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 2777 11067 2835 11073
rect 2777 11033 2789 11067
rect 2823 11064 2835 11067
rect 3878 11064 3884 11076
rect 2823 11036 3884 11064
rect 2823 11033 2835 11036
rect 2777 11027 2835 11033
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4448 11064 4476 11095
rect 4522 11064 4528 11076
rect 4448 11036 4528 11064
rect 4522 11024 4528 11036
rect 4580 11024 4586 11076
rect 4617 11067 4675 11073
rect 4617 11033 4629 11067
rect 4663 11064 4675 11067
rect 5276 11064 5304 11172
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5721 11203 5779 11209
rect 5721 11169 5733 11203
rect 5767 11200 5779 11203
rect 6546 11200 6552 11212
rect 5767 11172 5948 11200
rect 6507 11172 6552 11200
rect 5767 11169 5779 11172
rect 5721 11163 5779 11169
rect 5442 11132 5448 11144
rect 5403 11104 5448 11132
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 5534 11064 5540 11076
rect 4663 11036 5212 11064
rect 5276 11036 5540 11064
rect 4663 11033 4675 11036
rect 4617 11027 4675 11033
rect 4154 10996 4160 11008
rect 4115 10968 4160 10996
rect 4154 10956 4160 10968
rect 4212 10956 4218 11008
rect 5184 10996 5212 11036
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 5350 10996 5356 11008
rect 5184 10968 5356 10996
rect 5350 10956 5356 10968
rect 5408 10956 5414 11008
rect 5718 10956 5724 11008
rect 5776 10996 5782 11008
rect 5920 10996 5948 11172
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11200 7895 11203
rect 8018 11200 8024 11212
rect 7883 11172 8024 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 9140 11209 9168 11240
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 9306 11160 9312 11212
rect 9364 11200 9370 11212
rect 9401 11203 9459 11209
rect 9401 11200 9413 11203
rect 9364 11172 9413 11200
rect 9364 11160 9370 11172
rect 9401 11169 9413 11172
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 9732 11172 11376 11200
rect 9732 11160 9738 11172
rect 6270 11132 6276 11144
rect 6231 11104 6276 11132
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 7558 11132 7564 11144
rect 7519 11104 7564 11132
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11101 8999 11135
rect 11238 11132 11244 11144
rect 11199 11104 11244 11132
rect 8941 11095 8999 11101
rect 5994 11024 6000 11076
rect 6052 11064 6058 11076
rect 6362 11064 6368 11076
rect 6052 11036 6368 11064
rect 6052 11024 6058 11036
rect 6362 11024 6368 11036
rect 6420 11024 6426 11076
rect 6638 11024 6644 11076
rect 6696 11064 6702 11076
rect 8956 11064 8984 11095
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 11348 11132 11376 11172
rect 12406 11132 12434 11308
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 13044 11308 13093 11336
rect 13044 11296 13050 11308
rect 13081 11305 13093 11308
rect 13127 11305 13139 11339
rect 13081 11299 13139 11305
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11336 13599 11339
rect 14642 11336 14648 11348
rect 13587 11308 14648 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 15286 11296 15292 11348
rect 15344 11336 15350 11348
rect 15562 11336 15568 11348
rect 15344 11308 15568 11336
rect 15344 11296 15350 11308
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 16114 11296 16120 11348
rect 16172 11336 16178 11348
rect 16482 11336 16488 11348
rect 16172 11308 16488 11336
rect 16172 11296 16178 11308
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 17313 11339 17371 11345
rect 17313 11305 17325 11339
rect 17359 11336 17371 11339
rect 17862 11336 17868 11348
rect 17359 11308 17868 11336
rect 17359 11305 17371 11308
rect 17313 11299 17371 11305
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 19702 11336 19708 11348
rect 19392 11308 19708 11336
rect 19392 11296 19398 11308
rect 19702 11296 19708 11308
rect 19760 11296 19766 11348
rect 20070 11336 20076 11348
rect 20031 11308 20076 11336
rect 20070 11296 20076 11308
rect 20128 11296 20134 11348
rect 20993 11339 21051 11345
rect 20993 11305 21005 11339
rect 21039 11336 21051 11339
rect 21082 11336 21088 11348
rect 21039 11308 21088 11336
rect 21039 11305 21051 11308
rect 20993 11299 21051 11305
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 22554 11336 22560 11348
rect 22515 11308 22560 11336
rect 22554 11296 22560 11308
rect 22612 11296 22618 11348
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 23477 11339 23535 11345
rect 23256 11308 23428 11336
rect 23256 11296 23262 11308
rect 13630 11268 13636 11280
rect 13188 11240 13636 11268
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13188 11209 13216 11240
rect 13630 11228 13636 11240
rect 13688 11228 13694 11280
rect 13906 11228 13912 11280
rect 13964 11268 13970 11280
rect 14734 11268 14740 11280
rect 13964 11240 14740 11268
rect 13964 11228 13970 11240
rect 14734 11228 14740 11240
rect 14792 11228 14798 11280
rect 15473 11271 15531 11277
rect 15473 11237 15485 11271
rect 15519 11268 15531 11271
rect 23290 11268 23296 11280
rect 15519 11240 16252 11268
rect 15519 11237 15531 11240
rect 15473 11231 15531 11237
rect 13173 11203 13231 11209
rect 13173 11200 13185 11203
rect 12952 11172 13185 11200
rect 12952 11160 12958 11172
rect 13173 11169 13185 11172
rect 13219 11169 13231 11203
rect 15105 11203 15163 11209
rect 15105 11200 15117 11203
rect 13173 11163 13231 11169
rect 13280 11172 15117 11200
rect 13280 11132 13308 11172
rect 15105 11169 15117 11172
rect 15151 11169 15163 11203
rect 15105 11163 15163 11169
rect 15194 11160 15200 11212
rect 15252 11160 15258 11212
rect 15838 11200 15844 11212
rect 15304 11172 15844 11200
rect 11348 11104 11652 11132
rect 12406 11104 13308 11132
rect 6696 11036 8984 11064
rect 6696 11024 6702 11036
rect 9122 11024 9128 11076
rect 9180 11064 9186 11076
rect 11486 11067 11544 11073
rect 11486 11064 11498 11067
rect 9180 11036 11498 11064
rect 9180 11024 9186 11036
rect 11486 11033 11498 11036
rect 11532 11033 11544 11067
rect 11624 11064 11652 11104
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 13412 11104 13457 11132
rect 13412 11092 13418 11104
rect 13538 11092 13544 11144
rect 13596 11132 13602 11144
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 13596 11104 14381 11132
rect 13596 11092 13602 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 14734 11132 14740 11144
rect 14507 11104 14740 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 14734 11092 14740 11104
rect 14792 11092 14798 11144
rect 13081 11067 13139 11073
rect 13081 11064 13093 11067
rect 11624 11036 13093 11064
rect 11486 11027 11544 11033
rect 13081 11033 13093 11036
rect 13127 11064 13139 11067
rect 13170 11064 13176 11076
rect 13127 11036 13176 11064
rect 13127 11033 13139 11036
rect 13081 11027 13139 11033
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 13998 11024 14004 11076
rect 14056 11064 14062 11076
rect 14277 11067 14335 11073
rect 14277 11064 14289 11067
rect 14056 11036 14289 11064
rect 14056 11024 14062 11036
rect 14277 11033 14289 11036
rect 14323 11033 14335 11067
rect 14642 11064 14648 11076
rect 14555 11036 14648 11064
rect 14277 11027 14335 11033
rect 14642 11024 14648 11036
rect 14700 11064 14706 11076
rect 15212 11064 15240 11160
rect 15304 11141 15332 11172
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 16022 11200 16028 11212
rect 15983 11172 16028 11200
rect 16022 11160 16028 11172
rect 16080 11160 16086 11212
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11101 15623 11135
rect 15565 11095 15623 11101
rect 15580 11064 15608 11095
rect 15654 11092 15660 11144
rect 15712 11132 15718 11144
rect 16114 11132 16120 11144
rect 15712 11104 16120 11132
rect 15712 11092 15718 11104
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 14700 11036 15608 11064
rect 16224 11064 16252 11240
rect 16316 11240 20852 11268
rect 16316 11141 16344 11240
rect 17126 11160 17132 11212
rect 17184 11200 17190 11212
rect 18049 11203 18107 11209
rect 18049 11200 18061 11203
rect 17184 11172 18061 11200
rect 17184 11160 17190 11172
rect 18049 11169 18061 11172
rect 18095 11169 18107 11203
rect 20714 11200 20720 11212
rect 18049 11163 18107 11169
rect 18248 11172 20720 11200
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11101 16359 11135
rect 18248 11132 18276 11172
rect 20714 11160 20720 11172
rect 20772 11160 20778 11212
rect 20824 11200 20852 11240
rect 21468 11240 23296 11268
rect 21468 11200 21496 11240
rect 23290 11228 23296 11240
rect 23348 11228 23354 11280
rect 23400 11268 23428 11308
rect 23477 11305 23489 11339
rect 23523 11336 23535 11339
rect 23658 11336 23664 11348
rect 23523 11308 23664 11336
rect 23523 11305 23535 11308
rect 23477 11299 23535 11305
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 24394 11336 24400 11348
rect 24355 11308 24400 11336
rect 24394 11296 24400 11308
rect 24452 11296 24458 11348
rect 27246 11336 27252 11348
rect 27207 11308 27252 11336
rect 27246 11296 27252 11308
rect 27304 11296 27310 11348
rect 27801 11271 27859 11277
rect 27801 11268 27813 11271
rect 23400 11240 27813 11268
rect 27801 11237 27813 11240
rect 27847 11268 27859 11271
rect 28353 11271 28411 11277
rect 28353 11268 28365 11271
rect 27847 11240 28365 11268
rect 27847 11237 27859 11240
rect 27801 11231 27859 11237
rect 28353 11237 28365 11240
rect 28399 11268 28411 11271
rect 28997 11271 29055 11277
rect 28997 11268 29009 11271
rect 28399 11240 29009 11268
rect 28399 11237 28411 11240
rect 28353 11231 28411 11237
rect 28997 11237 29009 11240
rect 29043 11268 29055 11271
rect 32030 11268 32036 11280
rect 29043 11240 32036 11268
rect 29043 11237 29055 11240
rect 28997 11231 29055 11237
rect 32030 11228 32036 11240
rect 32088 11228 32094 11280
rect 20824 11172 21496 11200
rect 21637 11203 21695 11209
rect 21637 11169 21649 11203
rect 21683 11200 21695 11203
rect 23750 11200 23756 11212
rect 21683 11172 23756 11200
rect 21683 11169 21695 11172
rect 21637 11163 21695 11169
rect 23750 11160 23756 11172
rect 23808 11160 23814 11212
rect 24762 11160 24768 11212
rect 24820 11200 24826 11212
rect 25041 11203 25099 11209
rect 25041 11200 25053 11203
rect 24820 11172 25053 11200
rect 24820 11160 24826 11172
rect 25041 11169 25053 11172
rect 25087 11200 25099 11203
rect 26697 11203 26755 11209
rect 26697 11200 26709 11203
rect 25087 11172 26709 11200
rect 25087 11169 25099 11172
rect 25041 11163 25099 11169
rect 26697 11169 26709 11172
rect 26743 11169 26755 11203
rect 26697 11163 26755 11169
rect 18414 11132 18420 11144
rect 16301 11095 16359 11101
rect 16868 11104 18276 11132
rect 18375 11104 18420 11132
rect 16868 11064 16896 11104
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 18874 11092 18880 11144
rect 18932 11132 18938 11144
rect 19521 11135 19579 11141
rect 19521 11132 19533 11135
rect 18932 11104 19533 11132
rect 18932 11092 18938 11104
rect 19521 11101 19533 11104
rect 19567 11132 19579 11135
rect 20622 11132 20628 11144
rect 19567 11104 20628 11132
rect 19567 11101 19579 11104
rect 19521 11095 19579 11101
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 21358 11132 21364 11144
rect 20732 11104 21364 11132
rect 16224 11036 16896 11064
rect 16945 11067 17003 11073
rect 14700 11024 14706 11036
rect 16945 11033 16957 11067
rect 16991 11064 17003 11067
rect 17034 11064 17040 11076
rect 16991 11036 17040 11064
rect 16991 11033 17003 11036
rect 16945 11027 17003 11033
rect 17034 11024 17040 11036
rect 17092 11024 17098 11076
rect 17129 11067 17187 11073
rect 17129 11033 17141 11067
rect 17175 11064 17187 11067
rect 17175 11036 18000 11064
rect 17175 11033 17187 11036
rect 17129 11027 17187 11033
rect 8938 10996 8944 11008
rect 5776 10968 8944 10996
rect 5776 10956 5782 10968
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 12986 10996 12992 11008
rect 10836 10968 12992 10996
rect 10836 10956 10842 10968
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 14093 10999 14151 11005
rect 14093 10965 14105 10999
rect 14139 10996 14151 10999
rect 15010 10996 15016 11008
rect 14139 10968 15016 10996
rect 14139 10965 14151 10968
rect 14093 10959 14151 10965
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 15194 10956 15200 11008
rect 15252 10996 15258 11008
rect 16485 10999 16543 11005
rect 16485 10996 16497 10999
rect 15252 10968 16497 10996
rect 15252 10956 15258 10968
rect 16485 10965 16497 10968
rect 16531 10965 16543 10999
rect 16485 10959 16543 10965
rect 16666 10956 16672 11008
rect 16724 10996 16730 11008
rect 17144 10996 17172 11027
rect 16724 10968 17172 10996
rect 17972 10996 18000 11036
rect 18046 11024 18052 11076
rect 18104 11064 18110 11076
rect 18233 11067 18291 11073
rect 18233 11064 18245 11067
rect 18104 11036 18245 11064
rect 18104 11024 18110 11036
rect 18233 11033 18245 11036
rect 18279 11033 18291 11067
rect 18233 11027 18291 11033
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 19150 11064 19156 11076
rect 18748 11036 19156 11064
rect 18748 11024 18754 11036
rect 19150 11024 19156 11036
rect 19208 11024 19214 11076
rect 19337 11067 19395 11073
rect 19337 11033 19349 11067
rect 19383 11064 19395 11067
rect 20162 11064 20168 11076
rect 19383 11036 20168 11064
rect 19383 11033 19395 11036
rect 19337 11027 19395 11033
rect 20162 11024 20168 11036
rect 20220 11024 20226 11076
rect 20254 11024 20260 11076
rect 20312 11064 20318 11076
rect 20438 11064 20444 11076
rect 20312 11036 20357 11064
rect 20399 11036 20444 11064
rect 20312 11024 20318 11036
rect 20438 11024 20444 11036
rect 20496 11024 20502 11076
rect 20732 11064 20760 11104
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 22005 11135 22063 11141
rect 22005 11101 22017 11135
rect 22051 11132 22063 11135
rect 22830 11132 22836 11144
rect 22051 11104 22836 11132
rect 22051 11101 22063 11104
rect 22005 11095 22063 11101
rect 22830 11092 22836 11104
rect 22888 11092 22894 11144
rect 23658 11132 23664 11144
rect 23571 11104 23664 11132
rect 23658 11092 23664 11104
rect 23716 11132 23722 11144
rect 24210 11132 24216 11144
rect 23716 11104 24216 11132
rect 23716 11092 23722 11104
rect 24210 11092 24216 11104
rect 24268 11132 24274 11144
rect 24780 11132 24808 11160
rect 24268 11104 24808 11132
rect 24268 11092 24274 11104
rect 21082 11064 21088 11076
rect 20548 11036 20760 11064
rect 21043 11036 21088 11064
rect 18322 10996 18328 11008
rect 17972 10968 18328 10996
rect 16724 10956 16730 10968
rect 18322 10956 18328 10968
rect 18380 10956 18386 11008
rect 18782 10956 18788 11008
rect 18840 10996 18846 11008
rect 20548 10996 20576 11036
rect 21082 11024 21088 11036
rect 21140 11024 21146 11076
rect 21542 11024 21548 11076
rect 21600 11064 21606 11076
rect 21821 11067 21879 11073
rect 21821 11064 21833 11067
rect 21600 11036 21833 11064
rect 21600 11024 21606 11036
rect 21821 11033 21833 11036
rect 21867 11064 21879 11067
rect 21867 11036 22692 11064
rect 21867 11033 21879 11036
rect 21821 11027 21879 11033
rect 18840 10968 20576 10996
rect 18840 10956 18846 10968
rect 20622 10956 20628 11008
rect 20680 10996 20686 11008
rect 22462 10996 22468 11008
rect 20680 10968 22468 10996
rect 20680 10956 20686 10968
rect 22462 10956 22468 10968
rect 22520 10956 22526 11008
rect 22664 10996 22692 11036
rect 22738 11024 22744 11076
rect 22796 11064 22802 11076
rect 22922 11064 22928 11076
rect 22796 11036 22841 11064
rect 22883 11036 22928 11064
rect 22796 11024 22802 11036
rect 22922 11024 22928 11036
rect 22980 11024 22986 11076
rect 23845 11067 23903 11073
rect 23845 11033 23857 11067
rect 23891 11064 23903 11067
rect 24118 11064 24124 11076
rect 23891 11036 24124 11064
rect 23891 11033 23903 11036
rect 23845 11027 23903 11033
rect 24118 11024 24124 11036
rect 24176 11024 24182 11076
rect 24765 11067 24823 11073
rect 24765 11033 24777 11067
rect 24811 11064 24823 11067
rect 25682 11064 25688 11076
rect 24811 11036 25688 11064
rect 24811 11033 24823 11036
rect 24765 11027 24823 11033
rect 25682 11024 25688 11036
rect 25740 11024 25746 11076
rect 26234 11064 26240 11076
rect 26195 11036 26240 11064
rect 26234 11024 26240 11036
rect 26292 11024 26298 11076
rect 24302 10996 24308 11008
rect 22664 10968 24308 10996
rect 24302 10956 24308 10968
rect 24360 10956 24366 11008
rect 24670 10956 24676 11008
rect 24728 10996 24734 11008
rect 24857 10999 24915 11005
rect 24857 10996 24869 10999
rect 24728 10968 24869 10996
rect 24728 10956 24734 10968
rect 24857 10965 24869 10968
rect 24903 10965 24915 10999
rect 24857 10959 24915 10965
rect 1104 10906 44896 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 44896 10906
rect 1104 10832 44896 10854
rect 2130 10752 2136 10804
rect 2188 10752 2194 10804
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 2406 10792 2412 10804
rect 2363 10764 2412 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 2406 10752 2412 10764
rect 2464 10752 2470 10804
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3789 10795 3847 10801
rect 3789 10792 3801 10795
rect 3384 10764 3801 10792
rect 3384 10752 3390 10764
rect 3789 10761 3801 10764
rect 3835 10792 3847 10795
rect 5718 10792 5724 10804
rect 3835 10764 5724 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 7558 10792 7564 10804
rect 5859 10764 7564 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 7800 10764 8432 10792
rect 7800 10752 7806 10764
rect 2148 10724 2176 10752
rect 4433 10727 4491 10733
rect 4433 10724 4445 10727
rect 1412 10696 2452 10724
rect 1412 10665 1440 10696
rect 2424 10668 2452 10696
rect 2746 10696 4445 10724
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10625 1455 10659
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1397 10619 1455 10625
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 2130 10656 2136 10668
rect 2091 10628 2136 10656
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 2406 10616 2412 10668
rect 2464 10616 2470 10668
rect 566 10548 572 10600
rect 624 10588 630 10600
rect 624 10560 1716 10588
rect 624 10548 630 10560
rect 1578 10520 1584 10532
rect 1539 10492 1584 10520
rect 1578 10480 1584 10492
rect 1636 10480 1642 10532
rect 1688 10520 1716 10560
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 2746 10588 2774 10696
rect 4433 10693 4445 10696
rect 4479 10724 4491 10727
rect 5258 10724 5264 10736
rect 4479 10696 5264 10724
rect 4479 10693 4491 10696
rect 4433 10687 4491 10693
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 5534 10684 5540 10736
rect 5592 10724 5598 10736
rect 6454 10724 6460 10736
rect 5592 10696 5672 10724
rect 6415 10696 6460 10724
rect 5592 10684 5598 10696
rect 3234 10656 3240 10668
rect 3195 10628 3240 10656
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 3881 10659 3939 10665
rect 3881 10656 3893 10659
rect 3844 10628 3893 10656
rect 3844 10616 3850 10628
rect 3881 10625 3893 10628
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 4246 10616 4252 10668
rect 4304 10656 4310 10668
rect 4982 10656 4988 10668
rect 4304 10628 4988 10656
rect 4304 10616 4310 10628
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 5350 10656 5356 10668
rect 5311 10628 5356 10656
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5644 10665 5672 10696
rect 6454 10684 6460 10696
rect 6512 10684 6518 10736
rect 6638 10684 6644 10736
rect 6696 10724 6702 10736
rect 8294 10724 8300 10736
rect 6696 10696 8300 10724
rect 6696 10684 6702 10696
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 8404 10724 8432 10764
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 9585 10795 9643 10801
rect 9585 10792 9597 10795
rect 8536 10764 9597 10792
rect 8536 10752 8542 10764
rect 9585 10761 9597 10764
rect 9631 10792 9643 10795
rect 10502 10792 10508 10804
rect 9631 10764 10508 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 10594 10752 10600 10804
rect 10652 10792 10658 10804
rect 10870 10792 10876 10804
rect 10652 10764 10876 10792
rect 10652 10752 10658 10764
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12250 10792 12256 10804
rect 12032 10764 12256 10792
rect 12032 10752 12038 10764
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 13446 10792 13452 10804
rect 12492 10764 13452 10792
rect 12492 10752 12498 10764
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 14550 10792 14556 10804
rect 14511 10764 14556 10792
rect 14550 10752 14556 10764
rect 14608 10752 14614 10804
rect 14918 10792 14924 10804
rect 14879 10764 14924 10792
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 15286 10752 15292 10804
rect 15344 10792 15350 10804
rect 15654 10792 15660 10804
rect 15344 10764 15660 10792
rect 15344 10752 15350 10764
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 19426 10792 19432 10804
rect 15764 10764 19432 10792
rect 9490 10724 9496 10736
rect 8404 10696 9496 10724
rect 9490 10684 9496 10696
rect 9548 10684 9554 10736
rect 10134 10684 10140 10736
rect 10192 10724 10198 10736
rect 10192 10696 13492 10724
rect 10192 10684 10198 10696
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 5810 10656 5816 10668
rect 5675 10628 5816 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 6362 10656 6368 10668
rect 6323 10628 6368 10656
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 8573 10659 8631 10665
rect 7300 10628 8524 10656
rect 7300 10600 7328 10628
rect 2556 10560 2774 10588
rect 2556 10548 2562 10560
rect 4522 10548 4528 10600
rect 4580 10588 4586 10600
rect 5442 10588 5448 10600
rect 4580 10560 5448 10588
rect 4580 10548 4586 10560
rect 5442 10548 5448 10560
rect 5500 10588 5506 10600
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 5500 10560 5549 10588
rect 5500 10548 5506 10560
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 5537 10551 5595 10557
rect 6270 10548 6276 10600
rect 6328 10588 6334 10600
rect 7009 10591 7067 10597
rect 7009 10588 7021 10591
rect 6328 10560 7021 10588
rect 6328 10548 6334 10560
rect 7009 10557 7021 10560
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 7282 10548 7288 10600
rect 7340 10548 7346 10600
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 8297 10591 8355 10597
rect 8297 10588 8309 10591
rect 7432 10560 8309 10588
rect 7432 10548 7438 10560
rect 8297 10557 8309 10560
rect 8343 10557 8355 10591
rect 8297 10551 8355 10557
rect 3786 10520 3792 10532
rect 1688 10492 3792 10520
rect 3786 10480 3792 10492
rect 3844 10480 3850 10532
rect 4801 10523 4859 10529
rect 4801 10489 4813 10523
rect 4847 10520 4859 10523
rect 4847 10492 8340 10520
rect 4847 10489 4859 10492
rect 4801 10483 4859 10489
rect 8312 10464 8340 10492
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 2832 10424 3065 10452
rect 2832 10412 2838 10424
rect 3053 10421 3065 10424
rect 3099 10452 3111 10455
rect 3970 10452 3976 10464
rect 3099 10424 3976 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 4890 10452 4896 10464
rect 4851 10424 4896 10452
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 5534 10452 5540 10464
rect 5224 10424 5540 10452
rect 5224 10412 5230 10424
rect 5534 10412 5540 10424
rect 5592 10452 5598 10464
rect 5629 10455 5687 10461
rect 5629 10452 5641 10455
rect 5592 10424 5641 10452
rect 5592 10412 5598 10424
rect 5629 10421 5641 10424
rect 5675 10452 5687 10455
rect 6270 10452 6276 10464
rect 5675 10424 6276 10452
rect 5675 10421 5687 10424
rect 5629 10415 5687 10421
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7239 10455 7297 10461
rect 7239 10452 7251 10455
rect 7064 10424 7251 10452
rect 7064 10412 7070 10424
rect 7239 10421 7251 10424
rect 7285 10421 7297 10455
rect 7239 10415 7297 10421
rect 8294 10412 8300 10464
rect 8352 10412 8358 10464
rect 8496 10452 8524 10628
rect 8573 10625 8585 10659
rect 8619 10656 8631 10659
rect 10410 10656 10416 10668
rect 8619 10628 10416 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 10709 10659 10767 10665
rect 10709 10625 10721 10659
rect 10755 10656 10767 10659
rect 11606 10656 11612 10668
rect 10755 10628 11612 10656
rect 10755 10625 10767 10628
rect 10709 10619 10767 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 11784 10659 11842 10665
rect 11784 10625 11796 10659
rect 11830 10656 11842 10659
rect 13464 10656 13492 10696
rect 13538 10684 13544 10736
rect 13596 10724 13602 10736
rect 13596 10696 13641 10724
rect 15028 10696 15700 10724
rect 13596 10684 13602 10696
rect 13725 10659 13783 10665
rect 11830 10628 13400 10656
rect 13464 10628 13676 10656
rect 11830 10625 11842 10628
rect 11784 10619 11842 10625
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10588 11023 10591
rect 11238 10588 11244 10600
rect 11011 10560 11244 10588
rect 11011 10557 11023 10560
rect 10965 10551 11023 10557
rect 11238 10548 11244 10560
rect 11296 10588 11302 10600
rect 11514 10588 11520 10600
rect 11296 10560 11520 10588
rect 11296 10548 11302 10560
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 8662 10480 8668 10532
rect 8720 10520 8726 10532
rect 9766 10520 9772 10532
rect 8720 10492 9772 10520
rect 8720 10480 8726 10492
rect 9766 10480 9772 10492
rect 9824 10480 9830 10532
rect 12897 10523 12955 10529
rect 12897 10489 12909 10523
rect 12943 10520 12955 10523
rect 13262 10520 13268 10532
rect 12943 10492 13268 10520
rect 12943 10489 12955 10492
rect 12897 10483 12955 10489
rect 13262 10480 13268 10492
rect 13320 10480 13326 10532
rect 12710 10452 12716 10464
rect 8496 10424 12716 10452
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 13372 10452 13400 10628
rect 13446 10548 13452 10600
rect 13504 10588 13510 10600
rect 13648 10588 13676 10628
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 14274 10656 14280 10668
rect 13771 10628 14280 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10656 14795 10659
rect 14826 10656 14832 10668
rect 14783 10628 14832 10656
rect 14783 10625 14795 10628
rect 14737 10619 14795 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 15028 10665 15056 10696
rect 15013 10659 15071 10665
rect 15013 10625 15025 10659
rect 15059 10625 15071 10659
rect 15013 10619 15071 10625
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 13504 10560 13549 10588
rect 13648 10560 15485 10588
rect 13504 10548 13510 10560
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 15562 10548 15568 10600
rect 15620 10548 15626 10600
rect 15672 10588 15700 10696
rect 15764 10665 15792 10764
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 19705 10795 19763 10801
rect 19705 10761 19717 10795
rect 19751 10792 19763 10795
rect 19978 10792 19984 10804
rect 19751 10764 19984 10792
rect 19751 10761 19763 10764
rect 19705 10755 19763 10761
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 20717 10795 20775 10801
rect 20717 10761 20729 10795
rect 20763 10792 20775 10795
rect 21634 10792 21640 10804
rect 20763 10764 21640 10792
rect 20763 10761 20775 10764
rect 20717 10755 20775 10761
rect 21634 10752 21640 10764
rect 21692 10752 21698 10804
rect 22002 10752 22008 10804
rect 22060 10792 22066 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 22060 10764 22385 10792
rect 22060 10752 22066 10764
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 23385 10795 23443 10801
rect 23385 10761 23397 10795
rect 23431 10792 23443 10795
rect 23658 10792 23664 10804
rect 23431 10764 23664 10792
rect 23431 10761 23443 10764
rect 23385 10755 23443 10761
rect 23658 10752 23664 10764
rect 23716 10752 23722 10804
rect 24762 10752 24768 10804
rect 24820 10792 24826 10804
rect 25041 10795 25099 10801
rect 25041 10792 25053 10795
rect 24820 10764 25053 10792
rect 24820 10752 24826 10764
rect 25041 10761 25053 10764
rect 25087 10761 25099 10795
rect 25041 10755 25099 10761
rect 26694 10752 26700 10804
rect 26752 10792 26758 10804
rect 27525 10795 27583 10801
rect 27525 10792 27537 10795
rect 26752 10764 27537 10792
rect 26752 10752 26758 10764
rect 27525 10761 27537 10764
rect 27571 10761 27583 10795
rect 27525 10755 27583 10761
rect 28169 10795 28227 10801
rect 28169 10761 28181 10795
rect 28215 10792 28227 10795
rect 28258 10792 28264 10804
rect 28215 10764 28264 10792
rect 28215 10761 28227 10764
rect 28169 10755 28227 10761
rect 28258 10752 28264 10764
rect 28316 10752 28322 10804
rect 18233 10727 18291 10733
rect 18233 10724 18245 10727
rect 15856 10696 18245 10724
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 15856 10588 15884 10696
rect 18233 10693 18245 10696
rect 18279 10693 18291 10727
rect 19242 10724 19248 10736
rect 19155 10696 19248 10724
rect 18233 10687 18291 10693
rect 19242 10684 19248 10696
rect 19300 10724 19306 10736
rect 22186 10724 22192 10736
rect 19300 10696 22192 10724
rect 19300 10684 19306 10696
rect 22186 10684 22192 10696
rect 22244 10684 22250 10736
rect 22738 10684 22744 10736
rect 22796 10724 22802 10736
rect 23290 10724 23296 10736
rect 22796 10696 23296 10724
rect 22796 10684 22802 10696
rect 23290 10684 23296 10696
rect 23348 10724 23354 10736
rect 25498 10724 25504 10736
rect 23348 10696 25504 10724
rect 23348 10684 23354 10696
rect 25498 10684 25504 10696
rect 25556 10684 25562 10736
rect 25685 10727 25743 10733
rect 25685 10693 25697 10727
rect 25731 10724 25743 10727
rect 32122 10724 32128 10736
rect 25731 10696 32128 10724
rect 25731 10693 25743 10696
rect 25685 10687 25743 10693
rect 32122 10684 32128 10696
rect 32180 10684 32186 10736
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 18138 10656 18144 10668
rect 16632 10628 18144 10656
rect 16632 10616 16638 10628
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10656 18383 10659
rect 18371 10628 18644 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 17218 10588 17224 10600
rect 15672 10560 15884 10588
rect 17179 10560 17224 10588
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 17678 10588 17684 10600
rect 17639 10560 17684 10588
rect 17678 10548 17684 10560
rect 17736 10548 17742 10600
rect 18616 10588 18644 10628
rect 18690 10616 18696 10668
rect 18748 10656 18754 10668
rect 20346 10656 20352 10668
rect 18748 10628 20352 10656
rect 18748 10616 18754 10628
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 26970 10656 26976 10668
rect 20456 10628 26976 10656
rect 18966 10588 18972 10600
rect 18616 10560 18972 10588
rect 18966 10548 18972 10560
rect 19024 10588 19030 10600
rect 20165 10591 20223 10597
rect 19024 10560 20116 10588
rect 19024 10548 19030 10560
rect 13998 10520 14004 10532
rect 13959 10492 14004 10520
rect 13998 10480 14004 10492
rect 14056 10480 14062 10532
rect 14274 10480 14280 10532
rect 14332 10520 14338 10532
rect 14826 10520 14832 10532
rect 14332 10492 14832 10520
rect 14332 10480 14338 10492
rect 14826 10480 14832 10492
rect 14884 10480 14890 10532
rect 15580 10520 15608 10548
rect 16482 10520 16488 10532
rect 15580 10492 16488 10520
rect 16482 10480 16488 10492
rect 16540 10480 16546 10532
rect 17405 10523 17463 10529
rect 17405 10489 17417 10523
rect 17451 10520 17463 10523
rect 18506 10520 18512 10532
rect 17451 10492 18512 10520
rect 17451 10489 17463 10492
rect 17405 10483 17463 10489
rect 18506 10480 18512 10492
rect 18564 10480 18570 10532
rect 18874 10480 18880 10532
rect 18932 10520 18938 10532
rect 19886 10520 19892 10532
rect 18932 10492 18977 10520
rect 19847 10492 19892 10520
rect 18932 10480 18938 10492
rect 19886 10480 19892 10492
rect 19944 10480 19950 10532
rect 20088 10520 20116 10560
rect 20165 10557 20177 10591
rect 20211 10588 20223 10591
rect 20254 10588 20260 10600
rect 20211 10560 20260 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 20456 10520 20484 10628
rect 26970 10616 26976 10628
rect 27028 10616 27034 10668
rect 21358 10548 21364 10600
rect 21416 10588 21422 10600
rect 22002 10588 22008 10600
rect 21416 10560 22008 10588
rect 21416 10548 21422 10560
rect 22002 10548 22008 10560
rect 22060 10548 22066 10600
rect 24581 10591 24639 10597
rect 24581 10557 24593 10591
rect 24627 10588 24639 10591
rect 24670 10588 24676 10600
rect 24627 10560 24676 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 24670 10548 24676 10560
rect 24728 10548 24734 10600
rect 25590 10548 25596 10600
rect 25648 10588 25654 10600
rect 32214 10588 32220 10600
rect 25648 10560 32220 10588
rect 25648 10548 25654 10560
rect 32214 10548 32220 10560
rect 32272 10548 32278 10600
rect 20088 10492 20484 10520
rect 20530 10480 20536 10532
rect 20588 10520 20594 10532
rect 20588 10492 21956 10520
rect 20588 10480 20594 10492
rect 21928 10464 21956 10492
rect 23198 10480 23204 10532
rect 23256 10520 23262 10532
rect 30558 10520 30564 10532
rect 23256 10492 30564 10520
rect 23256 10480 23262 10492
rect 30558 10480 30564 10492
rect 30616 10480 30622 10532
rect 15194 10452 15200 10464
rect 13372 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 15930 10452 15936 10464
rect 15891 10424 15936 10452
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 16666 10452 16672 10464
rect 16627 10424 16672 10452
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 18782 10452 18788 10464
rect 18743 10424 18788 10452
rect 18782 10412 18788 10424
rect 18840 10412 18846 10464
rect 20990 10412 20996 10464
rect 21048 10452 21054 10464
rect 21177 10455 21235 10461
rect 21177 10452 21189 10455
rect 21048 10424 21189 10452
rect 21048 10412 21054 10424
rect 21177 10421 21189 10424
rect 21223 10421 21235 10455
rect 21910 10452 21916 10464
rect 21871 10424 21916 10452
rect 21177 10415 21235 10421
rect 21910 10412 21916 10424
rect 21968 10412 21974 10464
rect 24029 10455 24087 10461
rect 24029 10421 24041 10455
rect 24075 10452 24087 10455
rect 24118 10452 24124 10464
rect 24075 10424 24124 10452
rect 24075 10421 24087 10424
rect 24029 10415 24087 10421
rect 24118 10412 24124 10424
rect 24176 10412 24182 10464
rect 26237 10455 26295 10461
rect 26237 10421 26249 10455
rect 26283 10452 26295 10455
rect 26326 10452 26332 10464
rect 26283 10424 26332 10452
rect 26283 10421 26295 10424
rect 26237 10415 26295 10421
rect 26326 10412 26332 10424
rect 26384 10412 26390 10464
rect 1104 10362 44896 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 44896 10362
rect 1104 10288 44896 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 2682 10248 2688 10260
rect 1903 10220 2688 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 5534 10248 5540 10260
rect 2976 10220 5396 10248
rect 5495 10220 5540 10248
rect 2590 10180 2596 10192
rect 2551 10152 2596 10180
rect 2590 10140 2596 10152
rect 2648 10140 2654 10192
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 2314 10112 2320 10124
rect 1627 10084 2320 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 2314 10072 2320 10084
rect 2372 10072 2378 10124
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 2976 10044 3004 10220
rect 4157 10183 4215 10189
rect 4157 10149 4169 10183
rect 4203 10180 4215 10183
rect 4614 10180 4620 10192
rect 4203 10152 4620 10180
rect 4203 10149 4215 10152
rect 4157 10143 4215 10149
rect 4614 10140 4620 10152
rect 4672 10140 4678 10192
rect 4985 10183 5043 10189
rect 4985 10149 4997 10183
rect 5031 10180 5043 10183
rect 5074 10180 5080 10192
rect 5031 10152 5080 10180
rect 5031 10149 5043 10152
rect 4985 10143 5043 10149
rect 5074 10140 5080 10152
rect 5132 10140 5138 10192
rect 5368 10180 5396 10220
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 5997 10251 6055 10257
rect 5997 10217 6009 10251
rect 6043 10248 6055 10251
rect 6086 10248 6092 10260
rect 6043 10220 6092 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 6178 10208 6184 10260
rect 6236 10248 6242 10260
rect 7466 10248 7472 10260
rect 6236 10220 7472 10248
rect 6236 10208 6242 10220
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 8938 10248 8944 10260
rect 8899 10220 8944 10248
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 10594 10248 10600 10260
rect 9447 10220 10600 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 11606 10208 11612 10260
rect 11664 10248 11670 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 11664 10220 14105 10248
rect 11664 10208 11670 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 14461 10251 14519 10257
rect 14461 10217 14473 10251
rect 14507 10248 14519 10251
rect 14550 10248 14556 10260
rect 14507 10220 14556 10248
rect 14507 10217 14519 10220
rect 14461 10211 14519 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 15102 10208 15108 10260
rect 15160 10248 15166 10260
rect 17221 10251 17279 10257
rect 17221 10248 17233 10251
rect 15160 10220 17233 10248
rect 15160 10208 15166 10220
rect 17221 10217 17233 10220
rect 17267 10217 17279 10251
rect 17221 10211 17279 10217
rect 17586 10208 17592 10260
rect 17644 10248 17650 10260
rect 17954 10248 17960 10260
rect 17644 10220 17960 10248
rect 17644 10208 17650 10220
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 18138 10248 18144 10260
rect 18099 10220 18144 10248
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 18506 10208 18512 10260
rect 18564 10248 18570 10260
rect 18564 10220 21496 10248
rect 18564 10208 18570 10220
rect 7193 10183 7251 10189
rect 5368 10152 7144 10180
rect 3602 10112 3608 10124
rect 3068 10084 3608 10112
rect 3068 10053 3096 10084
rect 3602 10072 3608 10084
rect 3660 10072 3666 10124
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 4522 10112 4528 10124
rect 3936 10084 4528 10112
rect 3936 10072 3942 10084
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 5629 10115 5687 10121
rect 5629 10112 5641 10115
rect 5500 10084 5641 10112
rect 5500 10072 5506 10084
rect 5629 10081 5641 10084
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 5718 10072 5724 10124
rect 5776 10112 5782 10124
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 5776 10084 6561 10112
rect 5776 10072 5782 10084
rect 6549 10081 6561 10084
rect 6595 10081 6607 10115
rect 6549 10075 6607 10081
rect 6638 10072 6644 10124
rect 6696 10072 6702 10124
rect 2455 10016 3004 10044
rect 3053 10047 3111 10053
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 3053 10013 3065 10047
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 4062 10044 4068 10056
rect 3283 10016 4068 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 5810 10044 5816 10056
rect 4212 10016 5212 10044
rect 5771 10016 5816 10044
rect 4212 10004 4218 10016
rect 1397 9979 1455 9985
rect 1397 9945 1409 9979
rect 1443 9976 1455 9979
rect 2130 9976 2136 9988
rect 1443 9948 2136 9976
rect 1443 9945 1455 9948
rect 1397 9939 1455 9945
rect 2130 9936 2136 9948
rect 2188 9936 2194 9988
rect 2222 9936 2228 9988
rect 2280 9976 2286 9988
rect 3970 9976 3976 9988
rect 2280 9948 3976 9976
rect 2280 9936 2286 9948
rect 3970 9936 3976 9948
rect 4028 9936 4034 9988
rect 4522 9936 4528 9988
rect 4580 9976 4586 9988
rect 4617 9979 4675 9985
rect 4617 9976 4629 9979
rect 4580 9948 4629 9976
rect 4580 9936 4586 9948
rect 4617 9945 4629 9948
rect 4663 9945 4675 9979
rect 4617 9939 4675 9945
rect 3145 9911 3203 9917
rect 3145 9877 3157 9911
rect 3191 9908 3203 9911
rect 3878 9908 3884 9920
rect 3191 9880 3884 9908
rect 3191 9877 3203 9880
rect 3145 9871 3203 9877
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 5074 9908 5080 9920
rect 5035 9880 5080 9908
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5184 9908 5212 10016
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 6656 10044 6684 10072
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 6512 10016 6745 10044
rect 6512 10004 6518 10016
rect 6733 10013 6745 10016
rect 6779 10013 6791 10047
rect 7116 10044 7144 10152
rect 7193 10149 7205 10183
rect 7239 10180 7251 10183
rect 9214 10180 9220 10192
rect 7239 10152 9220 10180
rect 7239 10149 7251 10152
rect 7193 10143 7251 10149
rect 9214 10140 9220 10152
rect 9272 10140 9278 10192
rect 9861 10183 9919 10189
rect 9861 10149 9873 10183
rect 9907 10180 9919 10183
rect 10134 10180 10140 10192
rect 9907 10152 10140 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 12710 10140 12716 10192
rect 12768 10180 12774 10192
rect 12986 10180 12992 10192
rect 12768 10152 12992 10180
rect 12768 10140 12774 10152
rect 12986 10140 12992 10152
rect 13044 10180 13050 10192
rect 13081 10183 13139 10189
rect 13081 10180 13093 10183
rect 13044 10152 13093 10180
rect 13044 10140 13050 10152
rect 13081 10149 13093 10152
rect 13127 10149 13139 10183
rect 15286 10180 15292 10192
rect 15247 10152 15292 10180
rect 13081 10143 13139 10149
rect 15286 10140 15292 10152
rect 15344 10140 15350 10192
rect 15473 10183 15531 10189
rect 15473 10149 15485 10183
rect 15519 10180 15531 10183
rect 16758 10180 16764 10192
rect 15519 10152 16764 10180
rect 15519 10149 15531 10152
rect 15473 10143 15531 10149
rect 16758 10140 16764 10152
rect 16816 10140 16822 10192
rect 17405 10183 17463 10189
rect 17405 10149 17417 10183
rect 17451 10149 17463 10183
rect 17405 10143 17463 10149
rect 7742 10112 7748 10124
rect 7703 10084 7748 10112
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 7926 10112 7932 10124
rect 7887 10084 7932 10112
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 8018 10072 8024 10124
rect 8076 10112 8082 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8076 10084 9137 10112
rect 8076 10072 8082 10084
rect 9125 10081 9137 10084
rect 9171 10112 9183 10115
rect 9171 10084 9352 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 7116 10016 7411 10044
rect 6733 10007 6791 10013
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 5537 9979 5595 9985
rect 5537 9976 5549 9979
rect 5408 9948 5549 9976
rect 5408 9936 5414 9948
rect 5537 9945 5549 9948
rect 5583 9976 5595 9979
rect 6362 9976 6368 9988
rect 5583 9948 6368 9976
rect 5583 9945 5595 9948
rect 5537 9939 5595 9945
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 6638 9936 6644 9988
rect 6696 9976 6702 9988
rect 6825 9979 6883 9985
rect 6825 9976 6837 9979
rect 6696 9948 6837 9976
rect 6696 9936 6702 9948
rect 6825 9945 6837 9948
rect 6871 9976 6883 9979
rect 7282 9976 7288 9988
rect 6871 9948 7288 9976
rect 6871 9945 6883 9948
rect 6825 9939 6883 9945
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 7383 9976 7411 10016
rect 8938 10004 8944 10056
rect 8996 10044 9002 10056
rect 9217 10047 9275 10053
rect 8996 10016 9041 10044
rect 8996 10004 9002 10016
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9324 10044 9352 10084
rect 13538 10072 13544 10124
rect 13596 10112 13602 10124
rect 15562 10112 15568 10124
rect 13596 10084 15568 10112
rect 13596 10072 13602 10084
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 16393 10115 16451 10121
rect 16393 10112 16405 10115
rect 15712 10084 16405 10112
rect 15712 10072 15718 10084
rect 16393 10081 16405 10084
rect 16439 10081 16451 10115
rect 17420 10112 17448 10143
rect 17862 10140 17868 10192
rect 17920 10180 17926 10192
rect 18966 10180 18972 10192
rect 17920 10152 18972 10180
rect 17920 10140 17926 10152
rect 18966 10140 18972 10152
rect 19024 10140 19030 10192
rect 19334 10140 19340 10192
rect 19392 10180 19398 10192
rect 19521 10183 19579 10189
rect 19521 10180 19533 10183
rect 19392 10152 19533 10180
rect 19392 10140 19398 10152
rect 19521 10149 19533 10152
rect 19567 10149 19579 10183
rect 19521 10143 19579 10149
rect 19705 10183 19763 10189
rect 19705 10149 19717 10183
rect 19751 10180 19763 10183
rect 20530 10180 20536 10192
rect 19751 10152 20536 10180
rect 19751 10149 19763 10152
rect 19705 10143 19763 10149
rect 20530 10140 20536 10152
rect 20588 10140 20594 10192
rect 21468 10180 21496 10220
rect 21542 10208 21548 10260
rect 21600 10248 21606 10260
rect 22649 10251 22707 10257
rect 22649 10248 22661 10251
rect 21600 10220 22661 10248
rect 21600 10208 21606 10220
rect 22649 10217 22661 10220
rect 22695 10217 22707 10251
rect 23290 10248 23296 10260
rect 23251 10220 23296 10248
rect 22649 10211 22707 10217
rect 23290 10208 23296 10220
rect 23348 10208 23354 10260
rect 24854 10208 24860 10260
rect 24912 10248 24918 10260
rect 25041 10251 25099 10257
rect 25041 10248 25053 10251
rect 24912 10220 25053 10248
rect 24912 10208 24918 10220
rect 25041 10217 25053 10220
rect 25087 10217 25099 10251
rect 25041 10211 25099 10217
rect 26237 10251 26295 10257
rect 26237 10217 26249 10251
rect 26283 10248 26295 10251
rect 30650 10248 30656 10260
rect 26283 10220 30656 10248
rect 26283 10217 26295 10220
rect 26237 10211 26295 10217
rect 30650 10208 30656 10220
rect 30708 10208 30714 10260
rect 43346 10248 43352 10260
rect 43307 10220 43352 10248
rect 43346 10208 43352 10220
rect 43404 10208 43410 10260
rect 25498 10180 25504 10192
rect 21468 10152 25504 10180
rect 25498 10140 25504 10152
rect 25556 10180 25562 10192
rect 25593 10183 25651 10189
rect 25593 10180 25605 10183
rect 25556 10152 25605 10180
rect 25556 10140 25562 10152
rect 25593 10149 25605 10152
rect 25639 10149 25651 10183
rect 25593 10143 25651 10149
rect 25774 10140 25780 10192
rect 25832 10180 25838 10192
rect 26881 10183 26939 10189
rect 26881 10180 26893 10183
rect 25832 10152 26893 10180
rect 25832 10140 25838 10152
rect 26881 10149 26893 10152
rect 26927 10149 26939 10183
rect 26881 10143 26939 10149
rect 22646 10112 22652 10124
rect 17420 10084 22652 10112
rect 16393 10075 16451 10081
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 27246 10112 27252 10124
rect 27080 10084 27252 10112
rect 10410 10044 10416 10056
rect 9324 10016 10416 10044
rect 9217 10007 9275 10013
rect 7383 9948 8708 9976
rect 7650 9908 7656 9920
rect 5184 9880 7656 9908
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 8021 9911 8079 9917
rect 8021 9908 8033 9911
rect 7800 9880 8033 9908
rect 7800 9868 7806 9880
rect 8021 9877 8033 9880
rect 8067 9877 8079 9911
rect 8386 9908 8392 9920
rect 8347 9880 8392 9908
rect 8021 9871 8079 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8680 9908 8708 9948
rect 9030 9936 9036 9988
rect 9088 9976 9094 9988
rect 9232 9976 9260 10007
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10044 11299 10047
rect 11514 10044 11520 10056
rect 11287 10016 11520 10044
rect 11287 10013 11299 10016
rect 11241 10007 11299 10013
rect 11514 10004 11520 10016
rect 11572 10044 11578 10056
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11572 10016 11713 10044
rect 11572 10004 11578 10016
rect 11701 10013 11713 10016
rect 11747 10044 11759 10047
rect 12342 10044 12348 10056
rect 11747 10016 12348 10044
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 14274 10044 14280 10056
rect 14235 10016 14280 10044
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 14550 10004 14556 10056
rect 14608 10044 14614 10056
rect 15010 10044 15016 10056
rect 14608 10016 14653 10044
rect 14971 10016 15016 10044
rect 14608 10004 14614 10016
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 17678 10044 17684 10056
rect 16684 10016 17684 10044
rect 16684 9988 16712 10016
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 17862 10004 17868 10056
rect 17920 10044 17926 10056
rect 18690 10044 18696 10056
rect 17920 10016 18696 10044
rect 17920 10004 17926 10016
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 19242 10044 19248 10056
rect 19203 10016 19248 10044
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 20346 10004 20352 10056
rect 20404 10044 20410 10056
rect 21637 10047 21695 10053
rect 20404 10016 20760 10044
rect 20404 10004 20410 10016
rect 10594 9976 10600 9988
rect 9088 9948 9260 9976
rect 9646 9948 10600 9976
rect 9088 9936 9094 9948
rect 9646 9908 9674 9948
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 10996 9979 11054 9985
rect 10996 9945 11008 9979
rect 11042 9976 11054 9979
rect 11042 9948 11744 9976
rect 11042 9945 11054 9948
rect 10996 9939 11054 9945
rect 8680 9880 9674 9908
rect 11716 9908 11744 9948
rect 11790 9936 11796 9988
rect 11848 9976 11854 9988
rect 11946 9979 12004 9985
rect 11946 9976 11958 9979
rect 11848 9948 11958 9976
rect 11848 9936 11854 9948
rect 11946 9945 11958 9948
rect 11992 9945 12004 9979
rect 11946 9939 12004 9945
rect 16577 9979 16635 9985
rect 16577 9945 16589 9979
rect 16623 9976 16635 9979
rect 16666 9976 16672 9988
rect 16623 9948 16672 9976
rect 16623 9945 16635 9948
rect 16577 9939 16635 9945
rect 16666 9936 16672 9948
rect 16724 9936 16730 9988
rect 16758 9936 16764 9988
rect 16816 9976 16822 9988
rect 16816 9948 16861 9976
rect 16816 9936 16822 9948
rect 17218 9936 17224 9988
rect 17276 9976 17282 9988
rect 18325 9979 18383 9985
rect 18325 9976 18337 9979
rect 17276 9948 18337 9976
rect 17276 9936 17282 9948
rect 18325 9945 18337 9948
rect 18371 9945 18383 9979
rect 18506 9976 18512 9988
rect 18467 9948 18512 9976
rect 18325 9939 18383 9945
rect 18506 9936 18512 9948
rect 18564 9936 18570 9988
rect 20622 9985 20628 9988
rect 20441 9979 20499 9985
rect 20441 9945 20453 9979
rect 20487 9976 20499 9979
rect 20579 9979 20628 9985
rect 20487 9945 20516 9976
rect 20441 9939 20516 9945
rect 20579 9945 20591 9979
rect 20625 9945 20628 9979
rect 20579 9939 20628 9945
rect 12986 9908 12992 9920
rect 11716 9880 12992 9908
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 14274 9868 14280 9920
rect 14332 9908 14338 9920
rect 14918 9908 14924 9920
rect 14332 9880 14924 9908
rect 14332 9868 14338 9880
rect 14918 9868 14924 9880
rect 14976 9868 14982 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 19426 9908 19432 9920
rect 15252 9880 19432 9908
rect 15252 9868 15258 9880
rect 19426 9868 19432 9880
rect 19484 9868 19490 9920
rect 20488 9908 20516 9939
rect 20622 9936 20628 9939
rect 20680 9936 20686 9988
rect 20732 9985 20760 10016
rect 21637 10013 21649 10047
rect 21683 10044 21695 10047
rect 22462 10044 22468 10056
rect 21683 10016 22468 10044
rect 21683 10013 21695 10016
rect 21637 10007 21695 10013
rect 22462 10004 22468 10016
rect 22520 10004 22526 10056
rect 24581 10047 24639 10053
rect 24581 10013 24593 10047
rect 24627 10044 24639 10047
rect 25590 10044 25596 10056
rect 24627 10016 25596 10044
rect 24627 10013 24639 10016
rect 24581 10007 24639 10013
rect 25590 10004 25596 10016
rect 25648 10004 25654 10056
rect 27080 10053 27108 10084
rect 27246 10072 27252 10084
rect 27304 10112 27310 10124
rect 28350 10112 28356 10124
rect 27304 10084 28356 10112
rect 27304 10072 27310 10084
rect 28350 10072 28356 10084
rect 28408 10072 28414 10124
rect 27065 10047 27123 10053
rect 27065 10013 27077 10047
rect 27111 10013 27123 10047
rect 27065 10007 27123 10013
rect 27890 10004 27896 10056
rect 27948 10044 27954 10056
rect 28077 10047 28135 10053
rect 28077 10044 28089 10047
rect 27948 10016 28089 10044
rect 27948 10004 27954 10016
rect 28077 10013 28089 10016
rect 28123 10013 28135 10047
rect 28994 10044 29000 10056
rect 28955 10016 29000 10044
rect 28077 10007 28135 10013
rect 28994 10004 29000 10016
rect 29052 10044 29058 10056
rect 29549 10047 29607 10053
rect 29549 10044 29561 10047
rect 29052 10016 29561 10044
rect 29052 10004 29058 10016
rect 29549 10013 29561 10016
rect 29595 10013 29607 10047
rect 29549 10007 29607 10013
rect 43346 10004 43352 10056
rect 43404 10044 43410 10056
rect 43901 10047 43959 10053
rect 43901 10044 43913 10047
rect 43404 10016 43913 10044
rect 43404 10004 43410 10016
rect 43901 10013 43913 10016
rect 43947 10013 43959 10047
rect 43901 10007 43959 10013
rect 20717 9979 20775 9985
rect 20717 9945 20729 9979
rect 20763 9945 20775 9979
rect 20717 9939 20775 9945
rect 21011 9979 21069 9985
rect 21011 9945 21023 9979
rect 21057 9976 21069 9979
rect 21174 9976 21180 9988
rect 21057 9948 21180 9976
rect 21057 9945 21069 9948
rect 21011 9939 21069 9945
rect 21174 9936 21180 9948
rect 21232 9936 21238 9988
rect 24854 9976 24860 9988
rect 21284 9948 24860 9976
rect 21284 9908 21312 9948
rect 24854 9936 24860 9948
rect 24912 9936 24918 9988
rect 25498 9936 25504 9988
rect 25556 9976 25562 9988
rect 26786 9976 26792 9988
rect 25556 9948 26792 9976
rect 25556 9936 25562 9948
rect 26786 9936 26792 9948
rect 26844 9936 26850 9988
rect 20488 9880 21312 9908
rect 21726 9868 21732 9920
rect 21784 9908 21790 9920
rect 22002 9908 22008 9920
rect 21784 9880 22008 9908
rect 21784 9868 21790 9880
rect 22002 9868 22008 9880
rect 22060 9908 22066 9920
rect 22097 9911 22155 9917
rect 22097 9908 22109 9911
rect 22060 9880 22109 9908
rect 22060 9868 22066 9880
rect 22097 9877 22109 9880
rect 22143 9877 22155 9911
rect 22097 9871 22155 9877
rect 22186 9868 22192 9920
rect 22244 9908 22250 9920
rect 23753 9911 23811 9917
rect 23753 9908 23765 9911
rect 22244 9880 23765 9908
rect 22244 9868 22250 9880
rect 23753 9877 23765 9880
rect 23799 9908 23811 9911
rect 24026 9908 24032 9920
rect 23799 9880 24032 9908
rect 23799 9877 23811 9880
rect 23753 9871 23811 9877
rect 24026 9868 24032 9880
rect 24084 9868 24090 9920
rect 24302 9868 24308 9920
rect 24360 9908 24366 9920
rect 24397 9911 24455 9917
rect 24397 9908 24409 9911
rect 24360 9880 24409 9908
rect 24360 9868 24366 9880
rect 24397 9877 24409 9880
rect 24443 9877 24455 9911
rect 24397 9871 24455 9877
rect 27614 9868 27620 9920
rect 27672 9908 27678 9920
rect 27893 9911 27951 9917
rect 27893 9908 27905 9911
rect 27672 9880 27905 9908
rect 27672 9868 27678 9880
rect 27893 9877 27905 9880
rect 27939 9877 27951 9911
rect 27893 9871 27951 9877
rect 27982 9868 27988 9920
rect 28040 9908 28046 9920
rect 28813 9911 28871 9917
rect 28813 9908 28825 9911
rect 28040 9880 28825 9908
rect 28040 9868 28046 9880
rect 28813 9877 28825 9880
rect 28859 9877 28871 9911
rect 44082 9908 44088 9920
rect 44043 9880 44088 9908
rect 28813 9871 28871 9877
rect 44082 9868 44088 9880
rect 44140 9868 44146 9920
rect 1104 9818 44896 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 44896 9818
rect 1104 9744 44896 9766
rect 2222 9664 2228 9716
rect 2280 9704 2286 9716
rect 2406 9704 2412 9716
rect 2280 9676 2412 9704
rect 2280 9664 2286 9676
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 3602 9664 3608 9716
rect 3660 9704 3666 9716
rect 4338 9704 4344 9716
rect 3660 9676 4344 9704
rect 3660 9664 3666 9676
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 7009 9707 7067 9713
rect 6604 9676 6960 9704
rect 6604 9664 6610 9676
rect 1946 9596 1952 9648
rect 2004 9636 2010 9648
rect 2004 9608 2774 9636
rect 2004 9596 2010 9608
rect 1762 9568 1768 9580
rect 1723 9540 1768 9568
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 2406 9568 2412 9580
rect 2367 9540 2412 9568
rect 2406 9528 2412 9540
rect 2464 9528 2470 9580
rect 2746 9568 2774 9608
rect 3786 9596 3792 9648
rect 3844 9636 3850 9648
rect 3844 9608 5672 9636
rect 3844 9596 3850 9608
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 2746 9540 3341 9568
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4338 9568 4344 9580
rect 4203 9540 4344 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 4338 9528 4344 9540
rect 4396 9568 4402 9580
rect 4614 9568 4620 9580
rect 4396 9540 4620 9568
rect 4396 9528 4402 9540
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5166 9568 5172 9580
rect 4939 9540 5172 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 4908 9500 4936 9531
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 5644 9577 5672 9608
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 6932 9636 6960 9676
rect 7009 9673 7021 9707
rect 7055 9704 7067 9707
rect 7374 9704 7380 9716
rect 7055 9676 7380 9704
rect 7055 9673 7067 9676
rect 7009 9667 7067 9673
rect 7374 9664 7380 9676
rect 7432 9664 7438 9716
rect 8757 9707 8815 9713
rect 8757 9673 8769 9707
rect 8803 9704 8815 9707
rect 9122 9704 9128 9716
rect 8803 9676 9128 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 9306 9664 9312 9716
rect 9364 9664 9370 9716
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 9950 9704 9956 9716
rect 9824 9676 9956 9704
rect 9824 9664 9830 9676
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 10686 9704 10692 9716
rect 10560 9676 10692 9704
rect 10560 9664 10566 9676
rect 10686 9664 10692 9676
rect 10744 9704 10750 9716
rect 14550 9704 14556 9716
rect 10744 9676 14556 9704
rect 10744 9664 10750 9676
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 16942 9704 16948 9716
rect 15120 9676 16948 9704
rect 7282 9636 7288 9648
rect 5868 9608 6868 9636
rect 6932 9608 7288 9636
rect 5868 9596 5874 9608
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 5994 9568 6000 9580
rect 5675 9540 6000 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6362 9528 6368 9580
rect 6420 9568 6426 9580
rect 6840 9577 6868 9608
rect 7282 9596 7288 9608
rect 7340 9636 7346 9648
rect 7469 9639 7527 9645
rect 7469 9636 7481 9639
rect 7340 9608 7481 9636
rect 7340 9596 7346 9608
rect 7469 9605 7481 9608
rect 7515 9605 7527 9639
rect 9324 9636 9352 9664
rect 12989 9639 13047 9645
rect 12989 9636 13001 9639
rect 7469 9599 7527 9605
rect 7579 9608 8064 9636
rect 9324 9608 9720 9636
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6420 9540 6561 9568
rect 6420 9528 6426 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 7374 9568 7380 9580
rect 6871 9540 7380 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 3476 9472 4936 9500
rect 3476 9460 3482 9472
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 6733 9503 6791 9509
rect 6733 9500 6745 9503
rect 5500 9472 6745 9500
rect 5500 9460 5506 9472
rect 6733 9469 6745 9472
rect 6779 9500 6791 9503
rect 7579 9500 7607 9608
rect 7785 9571 7843 9577
rect 7785 9537 7797 9571
rect 7831 9568 7843 9571
rect 7926 9568 7932 9580
rect 7831 9540 7932 9568
rect 7831 9537 7843 9540
rect 7785 9531 7843 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 8036 9568 8064 9608
rect 8202 9568 8208 9580
rect 8036 9540 8208 9568
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 9364 9540 9597 9568
rect 9364 9528 9370 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 6779 9472 7607 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 7708 9472 7753 9500
rect 7708 9460 7714 9472
rect 8478 9460 8484 9512
rect 8536 9500 8542 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8536 9472 8861 9500
rect 8536 9460 8542 9472
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9490 9500 9496 9512
rect 9079 9472 9496 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 9692 9500 9720 9608
rect 12544 9608 13001 9636
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 9824 9540 11928 9568
rect 9824 9528 9830 9540
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9692 9472 9873 9500
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 10226 9460 10232 9512
rect 10284 9500 10290 9512
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 10284 9472 11529 9500
rect 10284 9460 10290 9472
rect 11517 9469 11529 9472
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 11793 9503 11851 9509
rect 11793 9500 11805 9503
rect 11664 9472 11805 9500
rect 11664 9460 11670 9472
rect 11793 9469 11805 9472
rect 11839 9469 11851 9503
rect 11900 9500 11928 9540
rect 12544 9500 12572 9608
rect 12989 9605 13001 9608
rect 13035 9605 13047 9639
rect 12989 9599 13047 9605
rect 14461 9639 14519 9645
rect 14461 9605 14473 9639
rect 14507 9636 14519 9639
rect 15120 9636 15148 9676
rect 16942 9664 16948 9676
rect 17000 9664 17006 9716
rect 17770 9664 17776 9716
rect 17828 9704 17834 9716
rect 17828 9676 18828 9704
rect 17828 9664 17834 9676
rect 14507 9608 15148 9636
rect 14507 9605 14519 9608
rect 14461 9599 14519 9605
rect 15838 9596 15844 9648
rect 15896 9636 15902 9648
rect 15933 9639 15991 9645
rect 15933 9636 15945 9639
rect 15896 9608 15945 9636
rect 15896 9596 15902 9608
rect 15933 9605 15945 9608
rect 15979 9605 15991 9639
rect 15933 9599 15991 9605
rect 16669 9639 16727 9645
rect 16669 9605 16681 9639
rect 16715 9636 16727 9639
rect 17678 9636 17684 9648
rect 16715 9608 17684 9636
rect 16715 9605 16727 9608
rect 16669 9599 16727 9605
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 17957 9639 18015 9645
rect 17957 9605 17969 9639
rect 18003 9636 18015 9639
rect 18003 9608 18276 9636
rect 18003 9605 18015 9608
rect 17957 9599 18015 9605
rect 13173 9571 13231 9577
rect 13173 9537 13185 9571
rect 13219 9568 13231 9571
rect 13906 9568 13912 9580
rect 13219 9540 13912 9568
rect 13219 9537 13231 9540
rect 13173 9531 13231 9537
rect 13906 9528 13912 9540
rect 13964 9528 13970 9580
rect 14093 9571 14151 9577
rect 14093 9537 14105 9571
rect 14139 9568 14151 9571
rect 14139 9540 14964 9568
rect 14139 9537 14151 9540
rect 14093 9531 14151 9537
rect 11900 9472 12572 9500
rect 12897 9503 12955 9509
rect 11793 9463 11851 9469
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 12986 9500 12992 9512
rect 12943 9472 12992 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 14185 9503 14243 9509
rect 14185 9469 14197 9503
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9500 14335 9503
rect 14936 9500 14964 9540
rect 15010 9528 15016 9580
rect 15068 9568 15074 9580
rect 15105 9571 15163 9577
rect 15105 9568 15117 9571
rect 15068 9540 15117 9568
rect 15068 9528 15074 9540
rect 15105 9537 15117 9540
rect 15151 9537 15163 9571
rect 15286 9568 15292 9580
rect 15247 9540 15292 9568
rect 15105 9531 15163 9537
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 15746 9568 15752 9580
rect 15707 9540 15752 9568
rect 15746 9528 15752 9540
rect 15804 9528 15810 9580
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 16390 9568 16396 9580
rect 16163 9540 16396 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16500 9540 16865 9568
rect 15194 9500 15200 9512
rect 14323 9472 14780 9500
rect 14936 9472 15200 9500
rect 14323 9469 14335 9472
rect 14277 9463 14335 9469
rect 1026 9392 1032 9444
rect 1084 9432 1090 9444
rect 2593 9435 2651 9441
rect 2593 9432 2605 9435
rect 1084 9404 2605 9432
rect 1084 9392 1090 9404
rect 2593 9401 2605 9404
rect 2639 9401 2651 9435
rect 3510 9432 3516 9444
rect 3471 9404 3516 9432
rect 2593 9395 2651 9401
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 3602 9392 3608 9444
rect 3660 9432 3666 9444
rect 3973 9435 4031 9441
rect 3973 9432 3985 9435
rect 3660 9404 3985 9432
rect 3660 9392 3666 9404
rect 3973 9401 3985 9404
rect 4019 9432 4031 9435
rect 5813 9435 5871 9441
rect 4019 9404 5764 9432
rect 4019 9401 4031 9404
rect 3973 9395 4031 9401
rect 1946 9364 1952 9376
rect 1907 9336 1952 9364
rect 1946 9324 1952 9336
rect 2004 9324 2010 9376
rect 5077 9367 5135 9373
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 5350 9364 5356 9376
rect 5123 9336 5356 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 5736 9364 5764 9404
rect 5813 9401 5825 9435
rect 5859 9432 5871 9435
rect 7834 9432 7840 9444
rect 5859 9404 7840 9432
rect 5859 9401 5871 9404
rect 5813 9395 5871 9401
rect 7834 9392 7840 9404
rect 7892 9392 7898 9444
rect 7929 9435 7987 9441
rect 7929 9401 7941 9435
rect 7975 9432 7987 9435
rect 13354 9432 13360 9444
rect 7975 9404 13360 9432
rect 7975 9401 7987 9404
rect 7929 9395 7987 9401
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 14200 9432 14228 9463
rect 14458 9432 14464 9444
rect 14200 9404 14464 9432
rect 14458 9392 14464 9404
rect 14516 9432 14522 9444
rect 14642 9432 14648 9444
rect 14516 9404 14648 9432
rect 14516 9392 14522 9404
rect 14642 9392 14648 9404
rect 14700 9392 14706 9444
rect 6178 9364 6184 9376
rect 5736 9336 6184 9364
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6328 9336 6561 9364
rect 6328 9324 6334 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 7466 9364 7472 9376
rect 7427 9336 7472 9364
rect 6549 9327 6607 9333
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 8018 9364 8024 9376
rect 7708 9336 8024 9364
rect 7708 9324 7714 9336
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 8352 9336 8401 9364
rect 8352 9324 8358 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 10870 9364 10876 9376
rect 10831 9336 10876 9364
rect 8389 9327 8447 9333
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 11940 9336 13461 9364
rect 11940 9324 11946 9336
rect 13449 9333 13461 9336
rect 13495 9333 13507 9367
rect 14752 9364 14780 9472
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 16500 9500 16528 9540
rect 16853 9537 16865 9540
rect 16899 9568 16911 9571
rect 17862 9568 17868 9580
rect 16899 9540 17868 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 17862 9528 17868 9540
rect 17920 9528 17926 9580
rect 18248 9568 18276 9608
rect 18322 9596 18328 9648
rect 18380 9636 18386 9648
rect 18506 9636 18512 9648
rect 18380 9608 18512 9636
rect 18380 9596 18386 9608
rect 18506 9596 18512 9608
rect 18564 9596 18570 9648
rect 18800 9636 18828 9676
rect 19058 9664 19064 9716
rect 19116 9704 19122 9716
rect 19153 9707 19211 9713
rect 19153 9704 19165 9707
rect 19116 9676 19165 9704
rect 19116 9664 19122 9676
rect 19153 9673 19165 9676
rect 19199 9673 19211 9707
rect 21910 9704 21916 9716
rect 19153 9667 19211 9673
rect 19260 9676 21916 9704
rect 19260 9636 19288 9676
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 22094 9704 22100 9716
rect 22020 9676 22100 9704
rect 18800 9608 19288 9636
rect 18248 9540 18644 9568
rect 15764 9472 16528 9500
rect 15764 9444 15792 9472
rect 16574 9460 16580 9512
rect 16632 9460 16638 9512
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 17218 9500 17224 9512
rect 16724 9472 17224 9500
rect 16724 9460 16730 9472
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 18046 9460 18052 9472
rect 18104 9460 18110 9512
rect 18233 9503 18291 9509
rect 18233 9469 18245 9503
rect 18279 9500 18291 9503
rect 18322 9500 18328 9512
rect 18279 9472 18328 9500
rect 18279 9469 18291 9472
rect 18233 9463 18291 9469
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 14918 9432 14924 9444
rect 14879 9404 14924 9432
rect 14918 9392 14924 9404
rect 14976 9392 14982 9444
rect 15746 9392 15752 9444
rect 15804 9392 15810 9444
rect 16482 9392 16488 9444
rect 16540 9432 16546 9444
rect 16592 9432 16620 9460
rect 16540 9404 16620 9432
rect 16540 9392 16546 9404
rect 17034 9392 17040 9444
rect 17092 9432 17098 9444
rect 17586 9432 17592 9444
rect 17092 9404 17137 9432
rect 17547 9404 17592 9432
rect 17092 9392 17098 9404
rect 17586 9392 17592 9404
rect 17644 9392 17650 9444
rect 18616 9432 18644 9540
rect 18800 9512 18828 9608
rect 20346 9596 20352 9648
rect 20404 9636 20410 9648
rect 20714 9636 20720 9648
rect 20404 9608 20720 9636
rect 20404 9596 20410 9608
rect 20714 9596 20720 9608
rect 20772 9636 20778 9648
rect 22020 9645 22048 9676
rect 22094 9664 22100 9676
rect 22152 9664 22158 9716
rect 25222 9704 25228 9716
rect 22204 9676 25228 9704
rect 21085 9639 21143 9645
rect 21085 9636 21097 9639
rect 20772 9608 21097 9636
rect 20772 9596 20778 9608
rect 21085 9605 21097 9608
rect 21131 9605 21143 9639
rect 21085 9599 21143 9605
rect 21997 9639 22055 9645
rect 21997 9605 22009 9639
rect 22043 9605 22055 9639
rect 22204 9636 22232 9676
rect 25222 9664 25228 9676
rect 25280 9664 25286 9716
rect 27246 9704 27252 9716
rect 27207 9676 27252 9704
rect 27246 9664 27252 9676
rect 27304 9664 27310 9716
rect 27890 9664 27896 9716
rect 27948 9704 27954 9716
rect 28169 9707 28227 9713
rect 28169 9704 28181 9707
rect 27948 9676 28181 9704
rect 27948 9664 27954 9676
rect 28169 9673 28181 9676
rect 28215 9673 28227 9707
rect 28169 9667 28227 9673
rect 24210 9636 24216 9648
rect 21997 9599 22055 9605
rect 22112 9608 22232 9636
rect 24171 9608 24216 9636
rect 20898 9568 20904 9580
rect 20859 9540 20904 9568
rect 20898 9528 20904 9540
rect 20956 9528 20962 9580
rect 21726 9568 21732 9580
rect 21008 9540 21732 9568
rect 18782 9500 18788 9512
rect 18695 9472 18788 9500
rect 18782 9460 18788 9472
rect 18840 9500 18846 9512
rect 18877 9503 18935 9509
rect 18877 9500 18889 9503
rect 18840 9472 18889 9500
rect 18840 9460 18846 9472
rect 18877 9469 18889 9472
rect 18923 9469 18935 9503
rect 19058 9500 19064 9512
rect 19019 9472 19064 9500
rect 18877 9463 18935 9469
rect 19058 9460 19064 9472
rect 19116 9460 19122 9512
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 19981 9503 20039 9509
rect 19981 9500 19993 9503
rect 19300 9472 19993 9500
rect 19300 9460 19306 9472
rect 19981 9469 19993 9472
rect 20027 9469 20039 9503
rect 21008 9500 21036 9540
rect 21726 9528 21732 9540
rect 21784 9528 21790 9580
rect 22112 9568 22140 9608
rect 24210 9596 24216 9608
rect 24268 9636 24274 9648
rect 24765 9639 24823 9645
rect 24765 9636 24777 9639
rect 24268 9608 24777 9636
rect 24268 9596 24274 9608
rect 24765 9605 24777 9608
rect 24811 9605 24823 9639
rect 25958 9636 25964 9648
rect 25919 9608 25964 9636
rect 24765 9599 24823 9605
rect 25958 9596 25964 9608
rect 26016 9596 26022 9648
rect 22020 9540 22140 9568
rect 22170 9571 22228 9577
rect 19981 9463 20039 9469
rect 20272 9472 21036 9500
rect 19886 9432 19892 9444
rect 18616 9404 19892 9432
rect 19886 9392 19892 9404
rect 19944 9392 19950 9444
rect 20272 9441 20300 9472
rect 20257 9435 20315 9441
rect 20257 9401 20269 9435
rect 20303 9401 20315 9435
rect 22020 9432 22048 9540
rect 22170 9537 22182 9571
rect 22216 9568 22228 9571
rect 22216 9540 22324 9568
rect 22216 9537 22228 9540
rect 22170 9531 22228 9537
rect 22296 9500 22324 9540
rect 22738 9528 22744 9580
rect 22796 9568 22802 9580
rect 23293 9571 23351 9577
rect 23293 9568 23305 9571
rect 22796 9540 23305 9568
rect 22796 9528 22802 9540
rect 23293 9537 23305 9540
rect 23339 9568 23351 9571
rect 26694 9568 26700 9580
rect 23339 9540 26700 9568
rect 23339 9537 23351 9540
rect 23293 9531 23351 9537
rect 26694 9528 26700 9540
rect 26752 9528 26758 9580
rect 23382 9500 23388 9512
rect 22296 9472 23388 9500
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 27338 9500 27344 9512
rect 23492 9472 27344 9500
rect 20257 9395 20315 9401
rect 20364 9404 22048 9432
rect 15102 9364 15108 9376
rect 14752 9336 15108 9364
rect 13449 9327 13507 9333
rect 15102 9324 15108 9336
rect 15160 9364 15166 9376
rect 16666 9364 16672 9376
rect 15160 9336 16672 9364
rect 15160 9324 15166 9336
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 16942 9324 16948 9376
rect 17000 9364 17006 9376
rect 17954 9364 17960 9376
rect 17000 9336 17960 9364
rect 17000 9324 17006 9336
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 19521 9367 19579 9373
rect 19521 9333 19533 9367
rect 19567 9364 19579 9367
rect 20364 9364 20392 9404
rect 22094 9392 22100 9444
rect 22152 9432 22158 9444
rect 22370 9432 22376 9444
rect 22152 9404 22376 9432
rect 22152 9392 22158 9404
rect 22370 9392 22376 9404
rect 22428 9392 22434 9444
rect 22462 9392 22468 9444
rect 22520 9432 22526 9444
rect 23492 9432 23520 9472
rect 27338 9460 27344 9472
rect 27396 9460 27402 9512
rect 22520 9404 23520 9432
rect 26145 9435 26203 9441
rect 22520 9392 22526 9404
rect 26145 9401 26157 9435
rect 26191 9432 26203 9435
rect 26191 9404 35894 9432
rect 26191 9401 26203 9404
rect 26145 9395 26203 9401
rect 19567 9336 20392 9364
rect 20441 9367 20499 9373
rect 19567 9333 19579 9336
rect 19521 9327 19579 9333
rect 20441 9333 20453 9367
rect 20487 9364 20499 9367
rect 20622 9364 20628 9376
rect 20487 9336 20628 9364
rect 20487 9333 20499 9336
rect 20441 9327 20499 9333
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 21269 9367 21327 9373
rect 21269 9333 21281 9367
rect 21315 9364 21327 9367
rect 21450 9364 21456 9376
rect 21315 9336 21456 9364
rect 21315 9333 21327 9336
rect 21269 9327 21327 9333
rect 21450 9324 21456 9336
rect 21508 9324 21514 9376
rect 21821 9367 21879 9373
rect 21821 9333 21833 9367
rect 21867 9364 21879 9367
rect 22554 9364 22560 9376
rect 21867 9336 22560 9364
rect 21867 9333 21879 9336
rect 21821 9327 21879 9333
rect 22554 9324 22560 9336
rect 22612 9324 22618 9376
rect 22646 9324 22652 9376
rect 22704 9364 22710 9376
rect 24857 9367 24915 9373
rect 22704 9336 22749 9364
rect 22704 9324 22710 9336
rect 24857 9333 24869 9367
rect 24903 9364 24915 9367
rect 27062 9364 27068 9376
rect 24903 9336 27068 9364
rect 24903 9333 24915 9336
rect 24857 9327 24915 9333
rect 27062 9324 27068 9336
rect 27120 9324 27126 9376
rect 35866 9364 35894 9404
rect 42150 9364 42156 9376
rect 35866 9336 42156 9364
rect 42150 9324 42156 9336
rect 42208 9324 42214 9376
rect 1104 9274 44896 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 44896 9274
rect 1104 9200 44896 9222
rect 1394 9160 1400 9172
rect 1355 9132 1400 9160
rect 1394 9120 1400 9132
rect 1452 9120 1458 9172
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 2041 9163 2099 9169
rect 2041 9160 2053 9163
rect 1728 9132 2053 9160
rect 1728 9120 1734 9132
rect 2041 9129 2053 9132
rect 2087 9129 2099 9163
rect 2041 9123 2099 9129
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 2685 9163 2743 9169
rect 2685 9160 2697 9163
rect 2188 9132 2697 9160
rect 2188 9120 2194 9132
rect 2685 9129 2697 9132
rect 2731 9129 2743 9163
rect 2685 9123 2743 9129
rect 4433 9163 4491 9169
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 5442 9160 5448 9172
rect 4479 9132 5448 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 5813 9163 5871 9169
rect 5813 9129 5825 9163
rect 5859 9160 5871 9163
rect 6730 9160 6736 9172
rect 5859 9132 6736 9160
rect 5859 9129 5871 9132
rect 5813 9123 5871 9129
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 6886 9132 7227 9160
rect 4985 9095 5043 9101
rect 4985 9061 4997 9095
rect 5031 9092 5043 9095
rect 5718 9092 5724 9104
rect 5031 9064 5724 9092
rect 5031 9061 5043 9064
rect 4985 9055 5043 9061
rect 5718 9052 5724 9064
rect 5776 9052 5782 9104
rect 6178 9052 6184 9104
rect 6236 9092 6242 9104
rect 6886 9092 6914 9132
rect 7098 9092 7104 9104
rect 6236 9064 6914 9092
rect 7059 9064 7104 9092
rect 6236 9052 6242 9064
rect 7098 9052 7104 9064
rect 7156 9052 7162 9104
rect 7199 9092 7227 9132
rect 7466 9120 7472 9172
rect 7524 9160 7530 9172
rect 7929 9163 7987 9169
rect 7929 9160 7941 9163
rect 7524 9132 7941 9160
rect 7524 9120 7530 9132
rect 7929 9129 7941 9132
rect 7975 9129 7987 9163
rect 7929 9123 7987 9129
rect 8389 9163 8447 9169
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 9030 9160 9036 9172
rect 8435 9132 9036 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9129 9183 9163
rect 11054 9160 11060 9172
rect 9125 9123 9183 9129
rect 9232 9132 11060 9160
rect 7650 9092 7656 9104
rect 7199 9064 7656 9092
rect 7650 9052 7656 9064
rect 7708 9092 7714 9104
rect 7834 9092 7840 9104
rect 7708 9064 7840 9092
rect 7708 9052 7714 9064
rect 7834 9052 7840 9064
rect 7892 9092 7898 9104
rect 7892 9064 8241 9092
rect 7892 9052 7898 9064
rect 1762 8984 1768 9036
rect 1820 9024 1826 9036
rect 1820 8996 7972 9024
rect 1820 8984 1826 8996
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 1544 8928 1593 8956
rect 1544 8916 1550 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 1762 8848 1768 8900
rect 1820 8888 1826 8900
rect 2240 8888 2268 8919
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 2924 8928 2969 8956
rect 2924 8916 2930 8928
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3786 8956 3792 8968
rect 3292 8928 3792 8956
rect 3292 8916 3298 8928
rect 3786 8916 3792 8928
rect 3844 8956 3850 8968
rect 4249 8959 4307 8965
rect 4249 8956 4261 8959
rect 3844 8928 4261 8956
rect 3844 8916 3850 8928
rect 4249 8925 4261 8928
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 4672 8928 5181 8956
rect 4672 8916 4678 8928
rect 5169 8925 5181 8928
rect 5215 8956 5227 8959
rect 5442 8956 5448 8968
rect 5215 8928 5448 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 5626 8956 5632 8968
rect 5587 8928 5632 8956
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 6273 8959 6331 8965
rect 6273 8956 6285 8959
rect 6144 8928 6285 8956
rect 6144 8916 6150 8928
rect 6273 8925 6285 8928
rect 6319 8925 6331 8959
rect 6454 8956 6460 8968
rect 6415 8928 6460 8956
rect 6273 8919 6331 8925
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 3326 8888 3332 8900
rect 1820 8860 3332 8888
rect 1820 8848 1826 8860
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 6178 8848 6184 8900
rect 6236 8888 6242 8900
rect 6564 8888 6592 8919
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 7282 8956 7288 8968
rect 6788 8928 7288 8956
rect 6788 8916 6794 8928
rect 7282 8916 7288 8928
rect 7340 8956 7346 8968
rect 7944 8956 7972 8996
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 8076 8996 8121 9024
rect 8076 8984 8082 8996
rect 8213 8965 8241 9064
rect 8662 9052 8668 9104
rect 8720 9092 8726 9104
rect 9140 9092 9168 9123
rect 8720 9064 9168 9092
rect 8720 9052 8726 9064
rect 8570 8984 8576 9036
rect 8628 9024 8634 9036
rect 9232 9033 9260 9132
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11974 9160 11980 9172
rect 11935 9132 11980 9160
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 13078 9120 13084 9172
rect 13136 9160 13142 9172
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 13136 9132 13185 9160
rect 13136 9120 13142 9132
rect 13173 9129 13185 9132
rect 13219 9129 13231 9163
rect 13173 9123 13231 9129
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 14182 9160 14188 9172
rect 14139 9132 14188 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 14366 9120 14372 9172
rect 14424 9160 14430 9172
rect 14737 9163 14795 9169
rect 14737 9160 14749 9163
rect 14424 9132 14749 9160
rect 14424 9120 14430 9132
rect 14737 9129 14749 9132
rect 14783 9129 14795 9163
rect 16482 9160 16488 9172
rect 16443 9132 16488 9160
rect 14737 9123 14795 9129
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16574 9120 16580 9172
rect 16632 9160 16638 9172
rect 16850 9160 16856 9172
rect 16632 9132 16856 9160
rect 16632 9120 16638 9132
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 17586 9160 17592 9172
rect 17276 9132 17592 9160
rect 17276 9120 17282 9132
rect 17586 9120 17592 9132
rect 17644 9120 17650 9172
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 19337 9163 19395 9169
rect 19337 9160 19349 9163
rect 18564 9132 19349 9160
rect 18564 9120 18570 9132
rect 19337 9129 19349 9132
rect 19383 9129 19395 9163
rect 19337 9123 19395 9129
rect 19797 9163 19855 9169
rect 19797 9129 19809 9163
rect 19843 9160 19855 9163
rect 20070 9160 20076 9172
rect 19843 9132 20076 9160
rect 19843 9129 19855 9132
rect 19797 9123 19855 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 20530 9160 20536 9172
rect 20272 9132 20536 9160
rect 9585 9095 9643 9101
rect 9585 9061 9597 9095
rect 9631 9092 9643 9095
rect 9950 9092 9956 9104
rect 9631 9064 9956 9092
rect 9631 9061 9643 9064
rect 9585 9055 9643 9061
rect 9950 9052 9956 9064
rect 10008 9052 10014 9104
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 10778 9092 10784 9104
rect 10284 9064 10784 9092
rect 10284 9052 10290 9064
rect 10778 9052 10784 9064
rect 10836 9092 10842 9104
rect 13538 9092 13544 9104
rect 10836 9064 13544 9092
rect 10836 9052 10842 9064
rect 13538 9052 13544 9064
rect 13596 9052 13602 9104
rect 13998 9052 14004 9104
rect 14056 9092 14062 9104
rect 14918 9092 14924 9104
rect 14056 9064 14924 9092
rect 14056 9052 14062 9064
rect 14918 9052 14924 9064
rect 14976 9052 14982 9104
rect 15930 9092 15936 9104
rect 15891 9064 15936 9092
rect 15930 9052 15936 9064
rect 15988 9052 15994 9104
rect 16025 9095 16083 9101
rect 16025 9061 16037 9095
rect 16071 9092 16083 9095
rect 16758 9092 16764 9104
rect 16071 9064 16764 9092
rect 16071 9061 16083 9064
rect 16025 9055 16083 9061
rect 16758 9052 16764 9064
rect 16816 9052 16822 9104
rect 18690 9092 18696 9104
rect 16960 9064 18696 9092
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 8628 8996 9229 9024
rect 8628 8984 8634 8996
rect 9217 8993 9229 8996
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 9364 8996 10333 9024
rect 9364 8984 9370 8996
rect 10321 8993 10333 8996
rect 10367 9024 10379 9027
rect 10962 9024 10968 9036
rect 10367 8996 10968 9024
rect 10367 8993 10379 8996
rect 10321 8987 10379 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 11974 9024 11980 9036
rect 11664 8996 11980 9024
rect 11664 8984 11670 8996
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 12618 9024 12624 9036
rect 12579 8996 12624 9024
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 13446 8984 13452 9036
rect 13504 9024 13510 9036
rect 16960 9024 16988 9064
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 19978 9092 19984 9104
rect 19939 9064 19984 9092
rect 19978 9052 19984 9064
rect 20036 9052 20042 9104
rect 13504 8996 16988 9024
rect 17037 9027 17095 9033
rect 13504 8984 13510 8996
rect 17037 8993 17049 9027
rect 17083 9024 17095 9027
rect 18417 9027 18475 9033
rect 17083 8996 18368 9024
rect 17083 8993 17095 8996
rect 17037 8987 17095 8993
rect 8198 8959 8256 8965
rect 7340 8928 7696 8956
rect 7944 8928 8156 8956
rect 7340 8916 7346 8928
rect 6236 8860 6592 8888
rect 6886 8860 7411 8888
rect 6236 8848 6242 8860
rect 6549 8823 6607 8829
rect 6549 8789 6561 8823
rect 6595 8820 6607 8823
rect 6886 8820 6914 8860
rect 6595 8792 6914 8820
rect 7009 8823 7067 8829
rect 6595 8789 6607 8792
rect 6549 8783 6607 8789
rect 7009 8789 7021 8823
rect 7055 8820 7067 8823
rect 7282 8820 7288 8832
rect 7055 8792 7288 8820
rect 7055 8789 7067 8792
rect 7009 8783 7067 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 7383 8820 7411 8860
rect 7466 8848 7472 8900
rect 7524 8888 7530 8900
rect 7668 8888 7696 8928
rect 7929 8891 7987 8897
rect 7929 8888 7941 8891
rect 7524 8860 7569 8888
rect 7668 8860 7941 8888
rect 7524 8848 7530 8860
rect 7929 8857 7941 8860
rect 7975 8857 7987 8891
rect 8128 8888 8156 8928
rect 8198 8925 8210 8959
rect 8244 8925 8256 8959
rect 8198 8919 8256 8925
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8478 8956 8484 8968
rect 8352 8928 8484 8956
rect 8352 8916 8358 8928
rect 8478 8916 8484 8928
rect 8536 8956 8542 8968
rect 8536 8928 9168 8956
rect 8536 8916 8542 8928
rect 9030 8888 9036 8900
rect 8128 8860 9036 8888
rect 7929 8851 7987 8857
rect 9030 8848 9036 8860
rect 9088 8848 9094 8900
rect 9140 8897 9168 8928
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 10045 8959 10103 8965
rect 9456 8928 9501 8956
rect 9456 8916 9462 8928
rect 10045 8925 10057 8959
rect 10091 8956 10103 8959
rect 10134 8956 10140 8968
rect 10091 8928 10140 8956
rect 10091 8925 10103 8928
rect 10045 8919 10103 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 10560 8928 12756 8956
rect 10560 8916 10566 8928
rect 9125 8891 9183 8897
rect 9125 8857 9137 8891
rect 9171 8888 9183 8891
rect 9674 8888 9680 8900
rect 9171 8860 9352 8888
rect 9171 8857 9183 8860
rect 9125 8851 9183 8857
rect 8110 8820 8116 8832
rect 7383 8792 8116 8820
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 9324 8820 9352 8860
rect 9508 8860 9680 8888
rect 9508 8820 9536 8860
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 11238 8848 11244 8900
rect 11296 8888 11302 8900
rect 11425 8891 11483 8897
rect 11425 8888 11437 8891
rect 11296 8860 11437 8888
rect 11296 8848 11302 8860
rect 11425 8857 11437 8860
rect 11471 8888 11483 8891
rect 11606 8888 11612 8900
rect 11471 8860 11612 8888
rect 11471 8857 11483 8860
rect 11425 8851 11483 8857
rect 11606 8848 11612 8860
rect 11664 8848 11670 8900
rect 11701 8891 11759 8897
rect 11701 8857 11713 8891
rect 11747 8888 11759 8891
rect 11790 8888 11796 8900
rect 11747 8860 11796 8888
rect 11747 8857 11759 8860
rect 11701 8851 11759 8857
rect 11790 8848 11796 8860
rect 11848 8848 11854 8900
rect 12728 8897 12756 8928
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 13412 8928 14289 8956
rect 13412 8916 13418 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14918 8956 14924 8968
rect 14277 8919 14335 8925
rect 14375 8928 14596 8956
rect 14879 8928 14924 8956
rect 12713 8891 12771 8897
rect 12713 8857 12725 8891
rect 12759 8857 12771 8891
rect 12713 8851 12771 8857
rect 12897 8891 12955 8897
rect 12897 8857 12909 8891
rect 12943 8888 12955 8891
rect 14375 8888 14403 8928
rect 12943 8860 14403 8888
rect 12943 8857 12955 8860
rect 12897 8851 12955 8857
rect 14568 8832 14596 8928
rect 14918 8916 14924 8928
rect 14976 8916 14982 8968
rect 16758 8916 16764 8968
rect 16816 8956 16822 8968
rect 17052 8956 17080 8987
rect 16816 8928 17080 8956
rect 16816 8916 16822 8928
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 17494 8956 17500 8968
rect 17276 8928 17500 8956
rect 17276 8916 17282 8928
rect 17494 8916 17500 8928
rect 17552 8916 17558 8968
rect 18340 8956 18368 8996
rect 18417 8993 18429 9027
rect 18463 9024 18475 9027
rect 20272 9024 20300 9132
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 24397 9163 24455 9169
rect 24397 9160 24409 9163
rect 22152 9132 24409 9160
rect 22152 9120 22158 9132
rect 24397 9129 24409 9132
rect 24443 9160 24455 9163
rect 24486 9160 24492 9172
rect 24443 9132 24492 9160
rect 24443 9129 24455 9132
rect 24397 9123 24455 9129
rect 24486 9120 24492 9132
rect 24544 9120 24550 9172
rect 25777 9163 25835 9169
rect 25777 9129 25789 9163
rect 25823 9160 25835 9163
rect 25958 9160 25964 9172
rect 25823 9132 25964 9160
rect 25823 9129 25835 9132
rect 25777 9123 25835 9129
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 26418 9120 26424 9172
rect 26476 9160 26482 9172
rect 26970 9160 26976 9172
rect 26476 9132 26976 9160
rect 26476 9120 26482 9132
rect 26970 9120 26976 9132
rect 27028 9120 27034 9172
rect 27062 9120 27068 9172
rect 27120 9160 27126 9172
rect 41414 9160 41420 9172
rect 27120 9132 41420 9160
rect 27120 9120 27126 9132
rect 41414 9120 41420 9132
rect 41472 9120 41478 9172
rect 20806 9052 20812 9104
rect 20864 9092 20870 9104
rect 21085 9095 21143 9101
rect 21085 9092 21097 9095
rect 20864 9064 21097 9092
rect 20864 9052 20870 9064
rect 21085 9061 21097 9064
rect 21131 9061 21143 9095
rect 21085 9055 21143 9061
rect 21177 9095 21235 9101
rect 21177 9061 21189 9095
rect 21223 9092 21235 9095
rect 22462 9092 22468 9104
rect 21223 9064 22468 9092
rect 21223 9061 21235 9064
rect 21177 9055 21235 9061
rect 22462 9052 22468 9064
rect 22520 9052 22526 9104
rect 23109 9095 23167 9101
rect 23109 9061 23121 9095
rect 23155 9092 23167 9095
rect 23658 9092 23664 9104
rect 23155 9064 23664 9092
rect 23155 9061 23167 9064
rect 23109 9055 23167 9061
rect 23658 9052 23664 9064
rect 23716 9092 23722 9104
rect 31202 9092 31208 9104
rect 23716 9064 31208 9092
rect 23716 9052 23722 9064
rect 31202 9052 31208 9064
rect 31260 9052 31266 9104
rect 33318 9092 33324 9104
rect 31726 9064 33324 9092
rect 20990 9024 20996 9036
rect 18463 8996 20300 9024
rect 20824 8996 20996 9024
rect 18463 8993 18475 8996
rect 18417 8987 18475 8993
rect 20824 8956 20852 8996
rect 20990 8984 20996 8996
rect 21048 8984 21054 9036
rect 22554 9024 22560 9036
rect 22515 8996 22560 9024
rect 22554 8984 22560 8996
rect 22612 8984 22618 9036
rect 24118 8984 24124 9036
rect 24176 9024 24182 9036
rect 27430 9024 27436 9036
rect 24176 8996 27436 9024
rect 24176 8984 24182 8996
rect 27430 8984 27436 8996
rect 27488 8984 27494 9036
rect 21634 8956 21640 8968
rect 18340 8928 20852 8956
rect 21595 8928 21640 8956
rect 21634 8916 21640 8928
rect 21692 8916 21698 8968
rect 22005 8959 22063 8965
rect 22005 8925 22017 8959
rect 22051 8956 22063 8959
rect 31726 8956 31754 9064
rect 33318 9052 33324 9064
rect 33376 9052 33382 9104
rect 22051 8928 31754 8956
rect 22051 8925 22063 8928
rect 22005 8919 22063 8925
rect 15105 8891 15163 8897
rect 15105 8857 15117 8891
rect 15151 8888 15163 8891
rect 15194 8888 15200 8900
rect 15151 8860 15200 8888
rect 15151 8857 15163 8860
rect 15105 8851 15163 8857
rect 15194 8848 15200 8860
rect 15252 8848 15258 8900
rect 15565 8891 15623 8897
rect 15565 8857 15577 8891
rect 15611 8888 15623 8891
rect 15746 8888 15752 8900
rect 15611 8860 15752 8888
rect 15611 8857 15623 8860
rect 15565 8851 15623 8857
rect 15746 8848 15752 8860
rect 15804 8848 15810 8900
rect 16853 8891 16911 8897
rect 16853 8857 16865 8891
rect 16899 8888 16911 8891
rect 17034 8888 17040 8900
rect 16899 8860 17040 8888
rect 16899 8857 16911 8860
rect 16853 8851 16911 8857
rect 17034 8848 17040 8860
rect 17092 8848 17098 8900
rect 18046 8888 18052 8900
rect 18007 8860 18052 8888
rect 18046 8848 18052 8860
rect 18104 8848 18110 8900
rect 18233 8891 18291 8897
rect 18233 8857 18245 8891
rect 18279 8888 18291 8891
rect 18506 8888 18512 8900
rect 18279 8860 18512 8888
rect 18279 8857 18291 8860
rect 18233 8851 18291 8857
rect 18506 8848 18512 8860
rect 18564 8888 18570 8900
rect 18564 8860 19334 8888
rect 18564 8848 18570 8860
rect 9324 8792 9536 8820
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 11517 8823 11575 8829
rect 11517 8820 11529 8823
rect 11388 8792 11529 8820
rect 11388 8780 11394 8792
rect 11517 8789 11529 8792
rect 11563 8789 11575 8823
rect 11517 8783 11575 8789
rect 12986 8780 12992 8832
rect 13044 8820 13050 8832
rect 13354 8820 13360 8832
rect 13044 8792 13360 8820
rect 13044 8780 13050 8792
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 14550 8780 14556 8832
rect 14608 8780 14614 8832
rect 14918 8780 14924 8832
rect 14976 8820 14982 8832
rect 16206 8820 16212 8832
rect 14976 8792 16212 8820
rect 14976 8780 14982 8792
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 16945 8823 17003 8829
rect 16945 8789 16957 8823
rect 16991 8820 17003 8823
rect 17494 8820 17500 8832
rect 16991 8792 17500 8820
rect 16991 8789 17003 8792
rect 16945 8783 17003 8789
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 19306 8820 19334 8860
rect 20070 8848 20076 8900
rect 20128 8848 20134 8900
rect 20254 8888 20260 8900
rect 20215 8860 20260 8888
rect 20254 8848 20260 8860
rect 20312 8848 20318 8900
rect 20346 8848 20352 8900
rect 20404 8888 20410 8900
rect 20717 8891 20775 8897
rect 20717 8888 20729 8891
rect 20404 8860 20729 8888
rect 20404 8848 20410 8860
rect 20717 8857 20729 8860
rect 20763 8857 20775 8891
rect 21821 8891 21879 8897
rect 21821 8888 21833 8891
rect 20717 8851 20775 8857
rect 20824 8860 21833 8888
rect 20088 8820 20116 8848
rect 20824 8820 20852 8860
rect 21821 8857 21833 8860
rect 21867 8857 21879 8891
rect 21821 8851 21879 8857
rect 23658 8848 23664 8900
rect 23716 8888 23722 8900
rect 23716 8860 23761 8888
rect 23716 8848 23722 8860
rect 26970 8848 26976 8900
rect 27028 8888 27034 8900
rect 27617 8891 27675 8897
rect 27617 8888 27629 8891
rect 27028 8860 27629 8888
rect 27028 8848 27034 8860
rect 27617 8857 27629 8860
rect 27663 8857 27675 8891
rect 27617 8851 27675 8857
rect 23750 8820 23756 8832
rect 19306 8792 20852 8820
rect 23711 8792 23756 8820
rect 23750 8780 23756 8792
rect 23808 8780 23814 8832
rect 23842 8780 23848 8832
rect 23900 8820 23906 8832
rect 24210 8820 24216 8832
rect 23900 8792 24216 8820
rect 23900 8780 23906 8792
rect 24210 8780 24216 8792
rect 24268 8780 24274 8832
rect 25038 8820 25044 8832
rect 24999 8792 25044 8820
rect 25038 8780 25044 8792
rect 25096 8780 25102 8832
rect 27706 8820 27712 8832
rect 27667 8792 27712 8820
rect 27706 8780 27712 8792
rect 27764 8780 27770 8832
rect 1104 8730 44896 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 44896 8730
rect 1104 8656 44896 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1854 8616 1860 8628
rect 1627 8588 1860 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 2372 8588 2697 8616
rect 2372 8576 2378 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 3418 8616 3424 8628
rect 3379 8588 3424 8616
rect 2685 8579 2743 8585
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4798 8616 4804 8628
rect 4571 8588 4804 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 5169 8619 5227 8625
rect 5169 8585 5181 8619
rect 5215 8616 5227 8619
rect 7190 8616 7196 8628
rect 5215 8588 7196 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 7300 8588 7389 8616
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 6641 8551 6699 8557
rect 6641 8548 6653 8551
rect 4028 8520 6653 8548
rect 4028 8508 4034 8520
rect 6641 8517 6653 8520
rect 6687 8517 6699 8551
rect 6822 8548 6828 8560
rect 6783 8520 6828 8548
rect 6641 8511 6699 8517
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 6914 8508 6920 8560
rect 6972 8548 6978 8560
rect 7300 8548 7328 8588
rect 7377 8585 7389 8588
rect 7423 8585 7435 8619
rect 7377 8579 7435 8585
rect 8496 8588 8708 8616
rect 6972 8520 7328 8548
rect 7561 8551 7619 8557
rect 6972 8508 6978 8520
rect 7208 8492 7236 8520
rect 7561 8517 7573 8551
rect 7607 8548 7619 8551
rect 7834 8548 7840 8560
rect 7607 8520 7840 8548
rect 7607 8517 7619 8520
rect 7561 8511 7619 8517
rect 7834 8508 7840 8520
rect 7892 8548 7898 8560
rect 7892 8520 8156 8548
rect 7892 8508 7898 8520
rect 1394 8480 1400 8492
rect 1355 8452 1400 8480
rect 1394 8440 1400 8452
rect 1452 8440 1458 8492
rect 2222 8480 2228 8492
rect 2183 8452 2228 8480
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 3142 8480 3148 8492
rect 2915 8452 3148 8480
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4706 8480 4712 8492
rect 4387 8452 4712 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 4982 8480 4988 8492
rect 4943 8452 4988 8480
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5684 8452 5825 8480
rect 5684 8440 5690 8452
rect 5813 8449 5825 8452
rect 5859 8480 5871 8483
rect 7006 8480 7012 8492
rect 5859 8452 7012 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7190 8440 7196 8492
rect 7248 8440 7254 8492
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 8128 8480 8156 8520
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 8496 8548 8524 8588
rect 8260 8520 8524 8548
rect 8680 8548 8708 8588
rect 8754 8576 8760 8628
rect 8812 8616 8818 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 8812 8588 8953 8616
rect 8812 8576 8818 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 8941 8579 8999 8585
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9950 8616 9956 8628
rect 9355 8588 9956 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10594 8616 10600 8628
rect 10555 8588 10600 8616
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 11422 8576 11428 8628
rect 11480 8616 11486 8628
rect 11609 8619 11667 8625
rect 11609 8616 11621 8619
rect 11480 8588 11621 8616
rect 11480 8576 11486 8588
rect 11609 8585 11621 8588
rect 11655 8585 11667 8619
rect 11609 8579 11667 8585
rect 12158 8576 12164 8628
rect 12216 8616 12222 8628
rect 12216 8588 12434 8616
rect 12216 8576 12222 8588
rect 8680 8520 10364 8548
rect 8260 8508 8266 8520
rect 9306 8480 9312 8492
rect 8128 8452 9312 8480
rect 7285 8443 7343 8449
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 7300 8412 7328 8443
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 10134 8480 10140 8492
rect 9548 8452 9628 8480
rect 10095 8452 10140 8480
rect 9548 8440 9554 8452
rect 7374 8412 7380 8424
rect 5316 8384 6040 8412
rect 7300 8384 7380 8412
rect 5316 8372 5322 8384
rect 3234 8304 3240 8356
rect 3292 8344 3298 8356
rect 5902 8344 5908 8356
rect 3292 8316 5908 8344
rect 3292 8304 3298 8316
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 6012 8344 6040 8384
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8381 8079 8415
rect 8294 8412 8300 8424
rect 8021 8375 8079 8381
rect 8128 8384 8300 8412
rect 6914 8344 6920 8356
rect 6012 8316 6920 8344
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 4062 8276 4068 8288
rect 3936 8248 4068 8276
rect 3936 8236 3942 8248
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 5442 8276 5448 8288
rect 5316 8248 5448 8276
rect 5316 8236 5322 8248
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 5629 8279 5687 8285
rect 5629 8245 5641 8279
rect 5675 8276 5687 8279
rect 6012 8276 6040 8316
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7561 8347 7619 8353
rect 7561 8313 7573 8347
rect 7607 8344 7619 8347
rect 7742 8344 7748 8356
rect 7607 8316 7748 8344
rect 7607 8313 7619 8316
rect 7561 8307 7619 8313
rect 7742 8304 7748 8316
rect 7800 8304 7806 8356
rect 8036 8288 8064 8375
rect 8128 8356 8156 8384
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 9122 8412 9128 8424
rect 8680 8384 9128 8412
rect 8680 8356 8708 8384
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9600 8421 9628 8452
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 10336 8489 10364 8520
rect 10778 8508 10784 8560
rect 10836 8548 10842 8560
rect 12176 8548 12204 8576
rect 10836 8520 12204 8548
rect 10836 8508 10842 8520
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 12158 8480 12164 8492
rect 12023 8452 12164 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 9401 8415 9459 8421
rect 9401 8381 9413 8415
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 8110 8304 8116 8356
rect 8168 8304 8174 8356
rect 8386 8344 8392 8356
rect 8347 8316 8392 8344
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 8662 8304 8668 8356
rect 8720 8304 8726 8356
rect 9416 8344 9444 8375
rect 9950 8372 9956 8424
rect 10008 8412 10014 8424
rect 10428 8412 10456 8443
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 12406 8480 12434 8588
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 15749 8619 15807 8625
rect 12768 8588 14596 8616
rect 12768 8576 12774 8588
rect 12802 8548 12808 8560
rect 12763 8520 12808 8548
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 13021 8551 13079 8557
rect 13021 8517 13033 8551
rect 13067 8548 13079 8551
rect 13446 8548 13452 8560
rect 13067 8520 13452 8548
rect 13067 8517 13079 8520
rect 13021 8511 13079 8517
rect 13446 8508 13452 8520
rect 13504 8508 13510 8560
rect 13633 8551 13691 8557
rect 13633 8517 13645 8551
rect 13679 8517 13691 8551
rect 13633 8511 13691 8517
rect 13849 8551 13907 8557
rect 13849 8517 13861 8551
rect 13895 8548 13907 8551
rect 14090 8548 14096 8560
rect 13895 8520 14096 8548
rect 13895 8517 13907 8520
rect 13849 8511 13907 8517
rect 13648 8480 13676 8511
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 14568 8557 14596 8588
rect 15749 8585 15761 8619
rect 15795 8616 15807 8619
rect 17862 8616 17868 8628
rect 15795 8588 17868 8616
rect 15795 8585 15807 8588
rect 15749 8579 15807 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 19150 8576 19156 8628
rect 19208 8616 19214 8628
rect 19337 8619 19395 8625
rect 19337 8616 19349 8619
rect 19208 8588 19349 8616
rect 19208 8576 19214 8588
rect 19337 8585 19349 8588
rect 19383 8585 19395 8619
rect 19337 8579 19395 8585
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 21634 8616 21640 8628
rect 20220 8588 21640 8616
rect 20220 8576 20226 8588
rect 21634 8576 21640 8588
rect 21692 8576 21698 8628
rect 21726 8576 21732 8628
rect 21784 8616 21790 8628
rect 22738 8616 22744 8628
rect 21784 8588 22744 8616
rect 21784 8576 21790 8588
rect 22738 8576 22744 8588
rect 22796 8576 22802 8628
rect 25498 8616 25504 8628
rect 25459 8588 25504 8616
rect 25498 8576 25504 8588
rect 25556 8576 25562 8628
rect 27706 8576 27712 8628
rect 27764 8616 27770 8628
rect 42978 8616 42984 8628
rect 27764 8588 42984 8616
rect 27764 8576 27770 8588
rect 42978 8576 42984 8588
rect 43036 8576 43042 8628
rect 14553 8551 14611 8557
rect 14553 8517 14565 8551
rect 14599 8517 14611 8551
rect 14553 8511 14611 8517
rect 14737 8551 14795 8557
rect 14737 8517 14749 8551
rect 14783 8548 14795 8551
rect 14918 8548 14924 8560
rect 14783 8520 14924 8548
rect 14783 8517 14795 8520
rect 14737 8511 14795 8517
rect 14918 8508 14924 8520
rect 14976 8508 14982 8560
rect 16206 8508 16212 8560
rect 16264 8548 16270 8560
rect 19242 8548 19248 8560
rect 16264 8520 19248 8548
rect 16264 8508 16270 8520
rect 19242 8508 19248 8520
rect 19300 8548 19306 8560
rect 19797 8551 19855 8557
rect 19797 8548 19809 8551
rect 19300 8520 19809 8548
rect 19300 8508 19306 8520
rect 19797 8517 19809 8520
rect 19843 8517 19855 8551
rect 19797 8511 19855 8517
rect 20070 8508 20076 8560
rect 20128 8548 20134 8560
rect 22554 8548 22560 8560
rect 20128 8520 22416 8548
rect 22515 8520 22560 8548
rect 20128 8508 20134 8520
rect 22388 8492 22416 8520
rect 22554 8508 22560 8520
rect 22612 8508 22618 8560
rect 23750 8508 23756 8560
rect 23808 8548 23814 8560
rect 40770 8548 40776 8560
rect 23808 8520 40776 8548
rect 23808 8508 23814 8520
rect 40770 8508 40776 8520
rect 40828 8508 40834 8560
rect 15562 8480 15568 8492
rect 12406 8452 13676 8480
rect 15304 8452 15568 8480
rect 10008 8384 10456 8412
rect 10008 8372 10014 8384
rect 11054 8372 11060 8424
rect 11112 8412 11118 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 11112 8384 12081 8412
rect 11112 8372 11118 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12342 8412 12348 8424
rect 12299 8384 12348 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 15102 8412 15108 8424
rect 13188 8384 15108 8412
rect 12710 8344 12716 8356
rect 9416 8316 12716 8344
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 13188 8353 13216 8384
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 13173 8347 13231 8353
rect 13173 8313 13185 8347
rect 13219 8313 13231 8347
rect 13173 8307 13231 8313
rect 14001 8347 14059 8353
rect 14001 8313 14013 8347
rect 14047 8344 14059 8347
rect 15304 8344 15332 8452
rect 15562 8440 15568 8452
rect 15620 8440 15626 8492
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 15804 8452 16681 8480
rect 15804 8440 15810 8452
rect 16669 8449 16681 8452
rect 16715 8480 16727 8483
rect 17589 8483 17647 8489
rect 17589 8480 17601 8483
rect 16715 8452 17601 8480
rect 16715 8449 16727 8452
rect 16669 8443 16727 8449
rect 17589 8449 17601 8452
rect 17635 8449 17647 8483
rect 17589 8443 17647 8449
rect 17770 8440 17776 8492
rect 17828 8480 17834 8492
rect 18325 8483 18383 8489
rect 18325 8480 18337 8483
rect 17828 8452 18337 8480
rect 17828 8440 17834 8452
rect 18325 8449 18337 8452
rect 18371 8449 18383 8483
rect 18506 8480 18512 8492
rect 18467 8452 18512 8480
rect 18325 8443 18383 8449
rect 18506 8440 18512 8452
rect 18564 8440 18570 8492
rect 18690 8480 18696 8492
rect 18651 8452 18696 8480
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 21266 8480 21272 8492
rect 19168 8452 21272 8480
rect 15841 8415 15899 8421
rect 15841 8412 15853 8415
rect 15672 8384 15853 8412
rect 14047 8316 15332 8344
rect 14047 8313 14059 8316
rect 14001 8307 14059 8313
rect 15378 8304 15384 8356
rect 15436 8344 15442 8356
rect 15436 8316 15481 8344
rect 15436 8304 15442 8316
rect 5675 8248 6040 8276
rect 5675 8245 5687 8248
rect 5629 8239 5687 8245
rect 8018 8236 8024 8288
rect 8076 8236 8082 8288
rect 8202 8236 8208 8288
rect 8260 8276 8266 8288
rect 8481 8279 8539 8285
rect 8481 8276 8493 8279
rect 8260 8248 8493 8276
rect 8260 8236 8266 8248
rect 8481 8245 8493 8248
rect 8527 8245 8539 8279
rect 8481 8239 8539 8245
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 10137 8279 10195 8285
rect 10137 8276 10149 8279
rect 9180 8248 10149 8276
rect 9180 8236 9186 8248
rect 10137 8245 10149 8248
rect 10183 8245 10195 8279
rect 12986 8276 12992 8288
rect 12947 8248 12992 8276
rect 10137 8239 10195 8245
rect 12986 8236 12992 8248
rect 13044 8236 13050 8288
rect 13538 8236 13544 8288
rect 13596 8276 13602 8288
rect 13817 8279 13875 8285
rect 13817 8276 13829 8279
rect 13596 8248 13829 8276
rect 13596 8236 13602 8248
rect 13817 8245 13829 8248
rect 13863 8245 13875 8279
rect 13817 8239 13875 8245
rect 15562 8236 15568 8288
rect 15620 8276 15626 8288
rect 15672 8276 15700 8384
rect 15841 8381 15853 8384
rect 15887 8381 15899 8415
rect 16022 8412 16028 8424
rect 15983 8384 16028 8412
rect 15841 8375 15899 8381
rect 16022 8372 16028 8384
rect 16080 8412 16086 8424
rect 16574 8412 16580 8424
rect 16080 8384 16580 8412
rect 16080 8372 16086 8384
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8412 17187 8415
rect 19168 8412 19196 8452
rect 21266 8440 21272 8452
rect 21324 8440 21330 8492
rect 22370 8440 22376 8492
rect 22428 8480 22434 8492
rect 23293 8483 23351 8489
rect 23293 8480 23305 8483
rect 22428 8452 23305 8480
rect 22428 8440 22434 8452
rect 23293 8449 23305 8452
rect 23339 8480 23351 8483
rect 24397 8483 24455 8489
rect 24397 8480 24409 8483
rect 23339 8452 24409 8480
rect 23339 8449 23351 8452
rect 23293 8443 23351 8449
rect 24397 8449 24409 8452
rect 24443 8480 24455 8483
rect 26326 8480 26332 8492
rect 24443 8452 26332 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 26326 8440 26332 8452
rect 26384 8440 26390 8492
rect 20254 8412 20260 8424
rect 17175 8384 19196 8412
rect 20215 8384 20260 8412
rect 17175 8381 17187 8384
rect 17129 8375 17187 8381
rect 20254 8372 20260 8384
rect 20312 8372 20318 8424
rect 20717 8415 20775 8421
rect 20717 8381 20729 8415
rect 20763 8412 20775 8415
rect 25958 8412 25964 8424
rect 20763 8384 25084 8412
rect 25919 8384 25964 8412
rect 20763 8381 20775 8384
rect 20717 8375 20775 8381
rect 16942 8344 16948 8356
rect 16903 8316 16948 8344
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 17586 8304 17592 8356
rect 17644 8344 17650 8356
rect 19518 8344 19524 8356
rect 17644 8316 19380 8344
rect 19479 8316 19524 8344
rect 17644 8304 17650 8316
rect 15620 8248 15700 8276
rect 15620 8236 15626 8248
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 16850 8276 16856 8288
rect 16724 8248 16856 8276
rect 16724 8236 16730 8248
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 17954 8236 17960 8288
rect 18012 8276 18018 8288
rect 18598 8276 18604 8288
rect 18012 8248 18604 8276
rect 18012 8236 18018 8248
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 19352 8276 19380 8316
rect 19518 8304 19524 8316
rect 19576 8304 19582 8356
rect 19886 8304 19892 8356
rect 19944 8344 19950 8356
rect 20346 8344 20352 8356
rect 19944 8316 20352 8344
rect 19944 8304 19950 8316
rect 20346 8304 20352 8316
rect 20404 8304 20410 8356
rect 20530 8344 20536 8356
rect 20491 8316 20536 8344
rect 20530 8304 20536 8316
rect 20588 8304 20594 8356
rect 20806 8304 20812 8356
rect 20864 8344 20870 8356
rect 20990 8344 20996 8356
rect 20864 8316 20996 8344
rect 20864 8304 20870 8316
rect 20990 8304 20996 8316
rect 21048 8304 21054 8356
rect 21266 8344 21272 8356
rect 21227 8316 21272 8344
rect 21266 8304 21272 8316
rect 21324 8304 21330 8356
rect 22738 8344 22744 8356
rect 21744 8316 22600 8344
rect 22699 8316 22744 8344
rect 21744 8276 21772 8316
rect 21910 8276 21916 8288
rect 19352 8248 21772 8276
rect 21871 8248 21916 8276
rect 21910 8236 21916 8248
rect 21968 8236 21974 8288
rect 22572 8276 22600 8316
rect 22738 8304 22744 8316
rect 22796 8304 22802 8356
rect 23474 8344 23480 8356
rect 23308 8316 23480 8344
rect 23308 8276 23336 8316
rect 23474 8304 23480 8316
rect 23532 8304 23538 8356
rect 23842 8344 23848 8356
rect 23803 8316 23848 8344
rect 23842 8304 23848 8316
rect 23900 8304 23906 8356
rect 25056 8344 25084 8384
rect 25958 8372 25964 8384
rect 26016 8372 26022 8424
rect 26878 8344 26884 8356
rect 25056 8316 26884 8344
rect 26878 8304 26884 8316
rect 26936 8304 26942 8356
rect 22572 8248 23336 8276
rect 23382 8236 23388 8288
rect 23440 8276 23446 8288
rect 24949 8279 25007 8285
rect 24949 8276 24961 8279
rect 23440 8248 24961 8276
rect 23440 8236 23446 8248
rect 24949 8245 24961 8248
rect 24995 8276 25007 8279
rect 28626 8276 28632 8288
rect 24995 8248 28632 8276
rect 24995 8245 25007 8248
rect 24949 8239 25007 8245
rect 28626 8236 28632 8248
rect 28684 8236 28690 8288
rect 1104 8186 44896 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 44896 8186
rect 1104 8112 44896 8134
rect 2038 8072 2044 8084
rect 1999 8044 2044 8072
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 2590 8072 2596 8084
rect 2551 8044 2596 8072
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 3234 8072 3240 8084
rect 3195 8044 3240 8072
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 3786 8072 3792 8084
rect 3747 8044 3792 8072
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 6178 8072 6184 8084
rect 6139 8044 6184 8072
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 6641 8075 6699 8081
rect 6641 8041 6653 8075
rect 6687 8072 6699 8075
rect 6730 8072 6736 8084
rect 6687 8044 6736 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7466 8072 7472 8084
rect 6972 8044 7472 8072
rect 6972 8032 6978 8044
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 7616 8044 9137 8072
rect 7616 8032 7622 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 10008 8044 10149 8072
rect 10008 8032 10014 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12124 8044 12633 8072
rect 12124 8032 12130 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 13044 8044 16574 8072
rect 13044 8032 13050 8044
rect 1210 7964 1216 8016
rect 1268 8004 1274 8016
rect 8205 8007 8263 8013
rect 8205 8004 8217 8007
rect 1268 7976 8217 8004
rect 1268 7964 1274 7976
rect 8205 7973 8217 7976
rect 8251 7973 8263 8007
rect 8205 7967 8263 7973
rect 8294 7964 8300 8016
rect 8352 8004 8358 8016
rect 9398 8004 9404 8016
rect 8352 7976 9404 8004
rect 8352 7964 8358 7976
rect 9398 7964 9404 7976
rect 9456 8004 9462 8016
rect 13262 8004 13268 8016
rect 9456 7976 13268 8004
rect 9456 7964 9462 7976
rect 13262 7964 13268 7976
rect 13320 7964 13326 8016
rect 15378 7964 15384 8016
rect 15436 8004 15442 8016
rect 15746 8004 15752 8016
rect 15436 7976 15752 8004
rect 15436 7964 15442 7976
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 16546 8004 16574 8044
rect 17402 8032 17408 8084
rect 17460 8072 17466 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17460 8044 17785 8072
rect 17460 8032 17466 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 18598 8072 18604 8084
rect 18559 8044 18604 8072
rect 17773 8035 17831 8041
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 19150 8032 19156 8084
rect 19208 8072 19214 8084
rect 22002 8072 22008 8084
rect 19208 8044 22008 8072
rect 19208 8032 19214 8044
rect 22002 8032 22008 8044
rect 22060 8032 22066 8084
rect 25038 8072 25044 8084
rect 24999 8044 25044 8072
rect 25038 8032 25044 8044
rect 25096 8032 25102 8084
rect 25590 8072 25596 8084
rect 25551 8044 25596 8072
rect 25590 8032 25596 8044
rect 25648 8032 25654 8084
rect 18414 8004 18420 8016
rect 16546 7976 18420 8004
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 25406 8004 25412 8016
rect 21008 7976 25412 8004
rect 5166 7896 5172 7948
rect 5224 7936 5230 7948
rect 5224 7908 6868 7936
rect 5224 7896 5230 7908
rect 6840 7880 6868 7908
rect 7926 7896 7932 7948
rect 7984 7936 7990 7948
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 7984 7908 9229 7936
rect 7984 7896 7990 7908
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10505 7939 10563 7945
rect 10008 7908 10456 7936
rect 10008 7896 10014 7908
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 5132 7840 6009 7868
rect 5132 7828 5138 7840
rect 5997 7837 6009 7840
rect 6043 7837 6055 7871
rect 6822 7868 6828 7880
rect 6783 7840 6828 7868
rect 5997 7831 6055 7837
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 7285 7871 7343 7877
rect 7285 7868 7297 7871
rect 7248 7840 7297 7868
rect 7248 7828 7254 7840
rect 7285 7837 7297 7840
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 7708 7840 9413 7868
rect 7708 7828 7714 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 10318 7868 10324 7880
rect 10279 7840 10324 7868
rect 9401 7831 9459 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10428 7868 10456 7908
rect 10505 7905 10517 7939
rect 10551 7936 10563 7939
rect 10686 7936 10692 7948
rect 10551 7908 10692 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 11977 7939 12035 7945
rect 11977 7936 11989 7939
rect 11572 7908 11989 7936
rect 11572 7896 11578 7908
rect 11977 7905 11989 7908
rect 12023 7905 12035 7939
rect 13170 7936 13176 7948
rect 13131 7908 13176 7936
rect 11977 7899 12035 7905
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 13354 7896 13360 7948
rect 13412 7936 13418 7948
rect 18138 7936 18144 7948
rect 13412 7908 17172 7936
rect 13412 7896 13418 7908
rect 10597 7871 10655 7877
rect 10597 7868 10609 7871
rect 10428 7840 10609 7868
rect 10597 7837 10609 7840
rect 10643 7868 10655 7871
rect 10778 7868 10784 7880
rect 10643 7840 10784 7868
rect 10643 7837 10655 7840
rect 10597 7831 10655 7837
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 13081 7871 13139 7877
rect 13081 7868 13093 7871
rect 11204 7840 13093 7868
rect 11204 7828 11210 7840
rect 13081 7837 13093 7840
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13872 7840 14289 7868
rect 13872 7828 13878 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 15010 7868 15016 7880
rect 14971 7840 15016 7868
rect 14277 7831 14335 7837
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15102 7828 15108 7880
rect 15160 7868 15166 7880
rect 15470 7868 15476 7880
rect 15160 7840 15476 7868
rect 15160 7828 15166 7840
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 15654 7868 15660 7880
rect 15615 7840 15660 7868
rect 15654 7828 15660 7840
rect 15712 7828 15718 7880
rect 16298 7868 16304 7880
rect 16259 7840 16304 7868
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 16942 7868 16948 7880
rect 16903 7840 16948 7868
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17144 7877 17172 7908
rect 17972 7908 18144 7936
rect 17972 7877 18000 7908
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7868 17187 7871
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17175 7840 17969 7868
rect 17175 7837 17187 7840
rect 17129 7831 17187 7837
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 19794 7868 19800 7880
rect 19755 7840 19800 7868
rect 17957 7831 18015 7837
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 21008 7877 21036 7976
rect 25406 7964 25412 7976
rect 25464 7964 25470 8016
rect 22370 7936 22376 7948
rect 22331 7908 22376 7936
rect 22370 7896 22376 7908
rect 22428 7896 22434 7948
rect 25130 7936 25136 7948
rect 22572 7908 25136 7936
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20993 7871 21051 7877
rect 20993 7837 21005 7871
rect 21039 7837 21051 7871
rect 20993 7831 21051 7837
rect 21453 7871 21511 7877
rect 21453 7837 21465 7871
rect 21499 7868 21511 7871
rect 21910 7868 21916 7880
rect 21499 7840 21916 7868
rect 21499 7837 21511 7840
rect 21453 7831 21511 7837
rect 1581 7803 1639 7809
rect 1581 7769 1593 7803
rect 1627 7800 1639 7803
rect 4893 7803 4951 7809
rect 4893 7800 4905 7803
rect 1627 7772 4905 7800
rect 1627 7769 1639 7772
rect 1581 7763 1639 7769
rect 4893 7769 4905 7772
rect 4939 7800 4951 7803
rect 4982 7800 4988 7812
rect 4939 7772 4988 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 4982 7760 4988 7772
rect 5040 7760 5046 7812
rect 6730 7760 6736 7812
rect 6788 7800 6794 7812
rect 7926 7800 7932 7812
rect 6788 7772 7788 7800
rect 7887 7772 7932 7800
rect 6788 7760 6794 7772
rect 3602 7692 3608 7744
rect 3660 7732 3666 7744
rect 4338 7732 4344 7744
rect 3660 7704 4344 7732
rect 3660 7692 3666 7704
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 5534 7732 5540 7744
rect 5495 7704 5540 7732
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 7469 7735 7527 7741
rect 7469 7701 7481 7735
rect 7515 7732 7527 7735
rect 7558 7732 7564 7744
rect 7515 7704 7564 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 7760 7732 7788 7772
rect 7926 7760 7932 7772
rect 7984 7760 7990 7812
rect 9125 7803 9183 7809
rect 9125 7800 9137 7803
rect 8036 7772 9137 7800
rect 8036 7732 8064 7772
rect 9125 7769 9137 7772
rect 9171 7769 9183 7803
rect 11885 7803 11943 7809
rect 11885 7800 11897 7803
rect 9125 7763 9183 7769
rect 10796 7772 11897 7800
rect 10796 7744 10824 7772
rect 11885 7769 11897 7772
rect 11931 7769 11943 7803
rect 14090 7800 14096 7812
rect 14051 7772 14096 7800
rect 11885 7763 11943 7769
rect 14090 7760 14096 7772
rect 14148 7760 14154 7812
rect 16022 7760 16028 7812
rect 16080 7800 16086 7812
rect 17313 7803 17371 7809
rect 16080 7772 17264 7800
rect 16080 7760 16086 7772
rect 7760 7704 8064 7732
rect 8386 7692 8392 7744
rect 8444 7732 8450 7744
rect 9582 7732 9588 7744
rect 8444 7704 8489 7732
rect 9543 7704 9588 7732
rect 8444 7692 8450 7704
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 10778 7692 10784 7744
rect 10836 7692 10842 7744
rect 11422 7732 11428 7744
rect 11383 7704 11428 7732
rect 11422 7692 11428 7704
rect 11480 7692 11486 7744
rect 11790 7732 11796 7744
rect 11751 7704 11796 7732
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 12989 7735 13047 7741
rect 12989 7701 13001 7735
rect 13035 7732 13047 7735
rect 13078 7732 13084 7744
rect 13035 7704 13084 7732
rect 13035 7701 13047 7704
rect 12989 7695 13047 7701
rect 13078 7692 13084 7704
rect 13136 7692 13142 7744
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 14829 7735 14887 7741
rect 14829 7732 14841 7735
rect 14056 7704 14841 7732
rect 14056 7692 14062 7704
rect 14829 7701 14841 7704
rect 14875 7701 14887 7735
rect 15470 7732 15476 7744
rect 15431 7704 15476 7732
rect 14829 7695 14887 7701
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 15562 7692 15568 7744
rect 15620 7732 15626 7744
rect 16117 7735 16175 7741
rect 16117 7732 16129 7735
rect 15620 7704 16129 7732
rect 15620 7692 15626 7704
rect 16117 7701 16129 7704
rect 16163 7701 16175 7735
rect 17236 7732 17264 7772
rect 17313 7769 17325 7803
rect 17359 7800 17371 7803
rect 17402 7800 17408 7812
rect 17359 7772 17408 7800
rect 17359 7769 17371 7772
rect 17313 7763 17371 7769
rect 17402 7760 17408 7772
rect 17460 7760 17466 7812
rect 18138 7800 18144 7812
rect 18099 7772 18144 7800
rect 18138 7760 18144 7772
rect 18196 7760 18202 7812
rect 20088 7800 20116 7831
rect 21910 7828 21916 7840
rect 21968 7828 21974 7880
rect 22002 7828 22008 7880
rect 22060 7868 22066 7880
rect 22572 7868 22600 7908
rect 25130 7896 25136 7908
rect 25188 7896 25194 7948
rect 22060 7840 22600 7868
rect 22649 7871 22707 7877
rect 22060 7828 22066 7840
rect 22649 7837 22661 7871
rect 22695 7868 22707 7871
rect 23382 7868 23388 7880
rect 22695 7840 23388 7868
rect 22695 7837 22707 7840
rect 22649 7831 22707 7837
rect 23382 7828 23388 7840
rect 23440 7828 23446 7880
rect 21266 7800 21272 7812
rect 20088 7772 21272 7800
rect 21266 7760 21272 7772
rect 21324 7760 21330 7812
rect 21358 7760 21364 7812
rect 21416 7800 21422 7812
rect 29178 7800 29184 7812
rect 21416 7772 29184 7800
rect 21416 7760 21422 7772
rect 29178 7760 29184 7772
rect 29236 7760 29242 7812
rect 20070 7732 20076 7744
rect 17236 7704 20076 7732
rect 16117 7695 16175 7701
rect 20070 7692 20076 7704
rect 20128 7692 20134 7744
rect 20806 7732 20812 7744
rect 20767 7704 20812 7732
rect 20806 7692 20812 7704
rect 20864 7692 20870 7744
rect 21634 7732 21640 7744
rect 21595 7704 21640 7732
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 22094 7692 22100 7744
rect 22152 7732 22158 7744
rect 23198 7732 23204 7744
rect 22152 7704 23204 7732
rect 22152 7692 22158 7704
rect 23198 7692 23204 7704
rect 23256 7692 23262 7744
rect 23750 7732 23756 7744
rect 23711 7704 23756 7732
rect 23750 7692 23756 7704
rect 23808 7692 23814 7744
rect 24394 7732 24400 7744
rect 24355 7704 24400 7732
rect 24394 7692 24400 7704
rect 24452 7692 24458 7744
rect 1104 7642 44896 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 44896 7642
rect 1104 7568 44896 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 3602 7528 3608 7540
rect 2179 7500 3608 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 3602 7488 3608 7500
rect 3660 7488 3666 7540
rect 3786 7488 3792 7540
rect 3844 7528 3850 7540
rect 4065 7531 4123 7537
rect 4065 7528 4077 7531
rect 3844 7500 4077 7528
rect 3844 7488 3850 7500
rect 4065 7497 4077 7500
rect 4111 7497 4123 7531
rect 4065 7491 4123 7497
rect 4985 7531 5043 7537
rect 4985 7497 4997 7531
rect 5031 7528 5043 7531
rect 5074 7528 5080 7540
rect 5031 7500 5080 7528
rect 5031 7497 5043 7500
rect 4985 7491 5043 7497
rect 2685 7463 2743 7469
rect 2685 7429 2697 7463
rect 2731 7460 2743 7463
rect 3237 7463 3295 7469
rect 2731 7432 3188 7460
rect 2731 7429 2743 7432
rect 2685 7423 2743 7429
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7392 1458 7404
rect 2866 7392 2872 7404
rect 1452 7364 2872 7392
rect 1452 7352 1458 7364
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 3160 7392 3188 7432
rect 3237 7429 3249 7463
rect 3283 7460 3295 7463
rect 5000 7460 5028 7491
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 6457 7531 6515 7537
rect 6457 7497 6469 7531
rect 6503 7528 6515 7531
rect 8113 7531 8171 7537
rect 8113 7528 8125 7531
rect 6503 7500 8125 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 8113 7497 8125 7500
rect 8159 7528 8171 7531
rect 8294 7528 8300 7540
rect 8159 7500 8300 7528
rect 8159 7497 8171 7500
rect 8113 7491 8171 7497
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 8846 7528 8852 7540
rect 8807 7500 8852 7528
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9309 7531 9367 7537
rect 9309 7497 9321 7531
rect 9355 7528 9367 7531
rect 9490 7528 9496 7540
rect 9355 7500 9496 7528
rect 9355 7497 9367 7500
rect 9309 7491 9367 7497
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 14458 7528 14464 7540
rect 10244 7500 13492 7528
rect 14419 7500 14464 7528
rect 3283 7432 5028 7460
rect 5813 7463 5871 7469
rect 3283 7429 3295 7432
rect 3237 7423 3295 7429
rect 5813 7429 5825 7463
rect 5859 7460 5871 7463
rect 8573 7463 8631 7469
rect 8573 7460 8585 7463
rect 5859 7432 8585 7460
rect 5859 7429 5871 7432
rect 5813 7423 5871 7429
rect 8573 7429 8585 7432
rect 8619 7460 8631 7463
rect 10244 7460 10272 7500
rect 10410 7460 10416 7472
rect 8619 7432 9168 7460
rect 8619 7429 8631 7432
rect 8573 7423 8631 7429
rect 9140 7416 9168 7432
rect 9416 7432 10272 7460
rect 10371 7432 10416 7460
rect 9416 7416 9444 7432
rect 10410 7420 10416 7432
rect 10468 7420 10474 7472
rect 12710 7420 12716 7472
rect 12768 7460 12774 7472
rect 12805 7463 12863 7469
rect 12805 7460 12817 7463
rect 12768 7432 12817 7460
rect 12768 7420 12774 7432
rect 12805 7429 12817 7432
rect 12851 7429 12863 7463
rect 12805 7423 12863 7429
rect 12989 7463 13047 7469
rect 12989 7429 13001 7463
rect 13035 7460 13047 7463
rect 13170 7460 13176 7472
rect 13035 7432 13176 7460
rect 13035 7429 13047 7432
rect 12989 7423 13047 7429
rect 13170 7420 13176 7432
rect 13228 7460 13234 7472
rect 13354 7460 13360 7472
rect 13228 7432 13360 7460
rect 13228 7420 13234 7432
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 13464 7460 13492 7500
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 21174 7528 21180 7540
rect 17236 7500 21180 7528
rect 14642 7460 14648 7472
rect 13464 7432 14648 7460
rect 14642 7420 14648 7432
rect 14700 7420 14706 7472
rect 14829 7463 14887 7469
rect 14829 7429 14841 7463
rect 14875 7460 14887 7463
rect 15930 7460 15936 7472
rect 14875 7432 15936 7460
rect 14875 7429 14887 7432
rect 14829 7423 14887 7429
rect 15930 7420 15936 7432
rect 15988 7420 15994 7472
rect 16942 7420 16948 7472
rect 17000 7460 17006 7472
rect 17236 7469 17264 7500
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 21634 7488 21640 7540
rect 21692 7528 21698 7540
rect 29546 7528 29552 7540
rect 21692 7500 29552 7528
rect 21692 7488 21698 7500
rect 29546 7488 29552 7500
rect 29604 7488 29610 7540
rect 17037 7463 17095 7469
rect 17037 7460 17049 7463
rect 17000 7432 17049 7460
rect 17000 7420 17006 7432
rect 17037 7429 17049 7432
rect 17083 7429 17095 7463
rect 17037 7423 17095 7429
rect 17221 7463 17279 7469
rect 17221 7429 17233 7463
rect 17267 7429 17279 7463
rect 17221 7423 17279 7429
rect 17586 7420 17592 7472
rect 17644 7460 17650 7472
rect 18414 7460 18420 7472
rect 17644 7432 18420 7460
rect 17644 7420 17650 7432
rect 18414 7420 18420 7432
rect 18472 7420 18478 7472
rect 18598 7420 18604 7472
rect 18656 7460 18662 7472
rect 18656 7432 18920 7460
rect 18656 7420 18662 7432
rect 5534 7392 5540 7404
rect 3160 7364 5540 7392
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6880 7364 6929 7392
rect 6880 7352 6886 7364
rect 6917 7361 6929 7364
rect 6963 7361 6975 7395
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 6917 7355 6975 7361
rect 7024 7364 7941 7392
rect 5258 7284 5264 7336
rect 5316 7324 5322 7336
rect 7024 7324 7052 7364
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8202 7352 8208 7404
rect 8260 7392 8266 7404
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8260 7364 8769 7392
rect 8260 7352 8266 7364
rect 8757 7361 8769 7364
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7392 8907 7395
rect 8938 7392 8944 7404
rect 8895 7364 8944 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 5316 7296 7052 7324
rect 5316 7284 5322 7296
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8864 7324 8892 7355
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9140 7388 9444 7416
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 11514 7392 11520 7404
rect 10643 7364 11520 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 9784 7324 9812 7355
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 11882 7392 11888 7404
rect 11843 7364 11888 7392
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 13630 7392 13636 7404
rect 13591 7364 13636 7392
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7392 15899 7395
rect 16482 7392 16488 7404
rect 15887 7364 16488 7392
rect 15887 7361 15899 7364
rect 15841 7355 15899 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 18892 7401 18920 7432
rect 19242 7420 19248 7472
rect 19300 7460 19306 7472
rect 21542 7460 21548 7472
rect 19300 7432 21548 7460
rect 19300 7420 19306 7432
rect 21542 7420 21548 7432
rect 21600 7420 21606 7472
rect 18877 7395 18935 7401
rect 16960 7364 18828 7392
rect 8352 7296 8892 7324
rect 9416 7296 9812 7324
rect 10321 7327 10379 7333
rect 8352 7284 8358 7296
rect 7466 7216 7472 7268
rect 7524 7256 7530 7268
rect 9416 7256 9444 7296
rect 10321 7293 10333 7327
rect 10367 7324 10379 7327
rect 10778 7324 10784 7336
rect 10367 7296 10784 7324
rect 10367 7293 10379 7296
rect 10321 7287 10379 7293
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 11974 7324 11980 7336
rect 11935 7296 11980 7324
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7324 12219 7327
rect 12250 7324 12256 7336
rect 12207 7296 12256 7324
rect 12207 7293 12219 7296
rect 12161 7287 12219 7293
rect 12250 7284 12256 7296
rect 12308 7324 12314 7336
rect 12710 7324 12716 7336
rect 12308 7296 12716 7324
rect 12308 7284 12314 7296
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14921 7327 14979 7333
rect 14921 7324 14933 7327
rect 13872 7296 14933 7324
rect 13872 7284 13878 7296
rect 14921 7293 14933 7296
rect 14967 7293 14979 7327
rect 14921 7287 14979 7293
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7324 15163 7327
rect 16022 7324 16028 7336
rect 15151 7296 16028 7324
rect 15151 7293 15163 7296
rect 15105 7287 15163 7293
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 16960 7333 16988 7364
rect 16945 7327 17003 7333
rect 16945 7293 16957 7327
rect 16991 7293 17003 7327
rect 16945 7287 17003 7293
rect 18601 7327 18659 7333
rect 18601 7293 18613 7327
rect 18647 7293 18659 7327
rect 18800 7324 18828 7364
rect 18877 7361 18889 7395
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7392 19395 7395
rect 19426 7392 19432 7404
rect 19383 7364 19432 7392
rect 19383 7361 19395 7364
rect 19337 7355 19395 7361
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 20254 7392 20260 7404
rect 19536 7364 20260 7392
rect 19536 7324 19564 7364
rect 20254 7352 20260 7364
rect 20312 7352 20318 7404
rect 20809 7396 20867 7401
rect 20809 7395 20944 7396
rect 20809 7361 20821 7395
rect 20855 7392 20944 7395
rect 22002 7392 22008 7404
rect 20855 7368 22008 7392
rect 20855 7361 20867 7368
rect 20916 7364 22008 7368
rect 20809 7355 20867 7361
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 22094 7352 22100 7404
rect 22152 7392 22158 7404
rect 23385 7395 23443 7401
rect 22152 7364 22197 7392
rect 22152 7352 22158 7364
rect 23385 7361 23397 7395
rect 23431 7392 23443 7395
rect 23750 7392 23756 7404
rect 23431 7364 23756 7392
rect 23431 7361 23443 7364
rect 23385 7355 23443 7361
rect 23750 7352 23756 7364
rect 23808 7392 23814 7404
rect 32582 7392 32588 7404
rect 23808 7364 32588 7392
rect 23808 7352 23814 7364
rect 32582 7352 32588 7364
rect 32640 7352 32646 7404
rect 18800 7296 19564 7324
rect 19613 7327 19671 7333
rect 18601 7287 18659 7293
rect 19613 7293 19625 7327
rect 19659 7324 19671 7327
rect 20714 7324 20720 7336
rect 19659 7296 20720 7324
rect 19659 7293 19671 7296
rect 19613 7287 19671 7293
rect 7524 7228 9444 7256
rect 7524 7216 7530 7228
rect 9490 7216 9496 7268
rect 9548 7256 9554 7268
rect 10873 7259 10931 7265
rect 9548 7228 9593 7256
rect 9548 7216 9554 7228
rect 10873 7225 10885 7259
rect 10919 7256 10931 7259
rect 11606 7256 11612 7268
rect 10919 7228 11612 7256
rect 10919 7225 10931 7228
rect 10873 7219 10931 7225
rect 11606 7216 11612 7228
rect 11664 7216 11670 7268
rect 17954 7256 17960 7268
rect 12268 7228 17960 7256
rect 12268 7200 12296 7228
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 18616 7256 18644 7287
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 22370 7324 22376 7336
rect 22331 7296 22376 7324
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 23661 7327 23719 7333
rect 23661 7293 23673 7327
rect 23707 7324 23719 7327
rect 24118 7324 24124 7336
rect 23707 7296 24124 7324
rect 23707 7293 23719 7296
rect 23661 7287 23719 7293
rect 24118 7284 24124 7296
rect 24176 7284 24182 7336
rect 28350 7256 28356 7268
rect 18616 7228 28356 7256
rect 28350 7216 28356 7228
rect 28408 7216 28414 7268
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 7101 7191 7159 7197
rect 7101 7188 7113 7191
rect 6420 7160 7113 7188
rect 6420 7148 6426 7160
rect 7101 7157 7113 7160
rect 7147 7188 7159 7191
rect 10134 7188 10140 7200
rect 7147 7160 10140 7188
rect 7147 7157 7159 7160
rect 7101 7151 7159 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 11480 7160 11529 7188
rect 11480 7148 11486 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 12250 7148 12256 7200
rect 12308 7148 12314 7200
rect 12986 7148 12992 7200
rect 13044 7188 13050 7200
rect 13449 7191 13507 7197
rect 13449 7188 13461 7191
rect 13044 7160 13461 7188
rect 13044 7148 13050 7160
rect 13449 7157 13461 7160
rect 13495 7157 13507 7191
rect 13449 7151 13507 7157
rect 14458 7148 14464 7200
rect 14516 7188 14522 7200
rect 15286 7188 15292 7200
rect 14516 7160 15292 7188
rect 14516 7148 14522 7160
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15657 7191 15715 7197
rect 15657 7157 15669 7191
rect 15703 7188 15715 7191
rect 15746 7188 15752 7200
rect 15703 7160 15752 7188
rect 15703 7157 15715 7160
rect 15657 7151 15715 7157
rect 15746 7148 15752 7160
rect 15804 7148 15810 7200
rect 17497 7191 17555 7197
rect 17497 7157 17509 7191
rect 17543 7188 17555 7191
rect 19978 7188 19984 7200
rect 17543 7160 19984 7188
rect 17543 7157 17555 7160
rect 17497 7151 17555 7157
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 20622 7188 20628 7200
rect 20583 7160 20628 7188
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 24762 7188 24768 7200
rect 24723 7160 24768 7188
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 1104 7098 44896 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 44896 7098
rect 1104 7024 44896 7046
rect 3326 6944 3332 6996
rect 3384 6984 3390 6996
rect 4798 6984 4804 6996
rect 3384 6956 4804 6984
rect 3384 6944 3390 6956
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 6270 6944 6276 6996
rect 6328 6984 6334 6996
rect 8389 6987 8447 6993
rect 8389 6984 8401 6987
rect 6328 6956 8401 6984
rect 6328 6944 6334 6956
rect 8389 6953 8401 6956
rect 8435 6984 8447 6987
rect 9122 6984 9128 6996
rect 8435 6956 9128 6984
rect 8435 6953 8447 6956
rect 8389 6947 8447 6953
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 9766 6984 9772 6996
rect 9272 6956 9772 6984
rect 9272 6944 9278 6956
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 10594 6944 10600 6996
rect 10652 6984 10658 6996
rect 10689 6987 10747 6993
rect 10689 6984 10701 6987
rect 10652 6956 10701 6984
rect 10652 6944 10658 6956
rect 10689 6953 10701 6956
rect 10735 6953 10747 6987
rect 10689 6947 10747 6953
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 12621 6987 12679 6993
rect 12621 6984 12633 6987
rect 12492 6956 12633 6984
rect 12492 6944 12498 6956
rect 12621 6953 12633 6956
rect 12667 6953 12679 6987
rect 12621 6947 12679 6953
rect 13262 6944 13268 6996
rect 13320 6984 13326 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 13320 6956 14105 6984
rect 13320 6944 13326 6956
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 17310 6984 17316 6996
rect 15252 6956 17316 6984
rect 15252 6944 15258 6956
rect 17310 6944 17316 6956
rect 17368 6944 17374 6996
rect 20438 6944 20444 6996
rect 20496 6984 20502 6996
rect 22646 6984 22652 6996
rect 20496 6956 22652 6984
rect 20496 6944 20502 6956
rect 22646 6944 22652 6956
rect 22704 6944 22710 6996
rect 2866 6876 2872 6928
rect 2924 6916 2930 6928
rect 7558 6916 7564 6928
rect 2924 6888 7564 6916
rect 2924 6876 2930 6888
rect 7558 6876 7564 6888
rect 7616 6876 7622 6928
rect 8570 6876 8576 6928
rect 8628 6916 8634 6928
rect 8754 6916 8760 6928
rect 8628 6888 8760 6916
rect 8628 6876 8634 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 9309 6919 9367 6925
rect 9309 6885 9321 6919
rect 9355 6885 9367 6919
rect 10962 6916 10968 6928
rect 9309 6879 9367 6885
rect 9600 6888 10968 6916
rect 4430 6848 4436 6860
rect 4391 6820 4436 6848
rect 4430 6808 4436 6820
rect 4488 6808 4494 6860
rect 5166 6848 5172 6860
rect 5127 6820 5172 6848
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 5721 6851 5779 6857
rect 5721 6817 5733 6851
rect 5767 6848 5779 6851
rect 6086 6848 6092 6860
rect 5767 6820 6092 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 7190 6848 7196 6860
rect 6871 6820 7196 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 7190 6808 7196 6820
rect 7248 6848 7254 6860
rect 9324 6848 9352 6879
rect 9600 6860 9628 6888
rect 10962 6876 10968 6888
rect 11020 6876 11026 6928
rect 11072 6888 13124 6916
rect 9398 6848 9404 6860
rect 7248 6820 8248 6848
rect 9324 6820 9404 6848
rect 7248 6808 7254 6820
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6780 1455 6783
rect 1486 6780 1492 6792
rect 1443 6752 1492 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 1486 6740 1492 6752
rect 1544 6740 1550 6792
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6780 6331 6783
rect 7098 6780 7104 6792
rect 6319 6752 7104 6780
rect 6319 6749 6331 6752
rect 6273 6743 6331 6749
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 7282 6780 7288 6792
rect 7243 6752 7288 6780
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 8220 6789 8248 6820
rect 9398 6808 9404 6820
rect 9456 6808 9462 6860
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 9640 6820 9733 6848
rect 9640 6808 9646 6820
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 11072 6848 11100 6888
rect 10744 6820 11100 6848
rect 11977 6851 12035 6857
rect 10744 6808 10750 6820
rect 11977 6817 11989 6851
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 11992 6780 12020 6811
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 12894 6848 12900 6860
rect 12124 6820 12900 6848
rect 12124 6808 12130 6820
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13096 6848 13124 6888
rect 14642 6876 14648 6928
rect 14700 6916 14706 6928
rect 17954 6916 17960 6928
rect 14700 6888 17960 6916
rect 14700 6876 14706 6888
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 19889 6919 19947 6925
rect 19889 6885 19901 6919
rect 19935 6885 19947 6919
rect 19889 6879 19947 6885
rect 13096 6820 13400 6848
rect 13096 6792 13124 6820
rect 8205 6743 8263 6749
rect 9140 6752 11008 6780
rect 11992 6752 12112 6780
rect 2593 6715 2651 6721
rect 2593 6681 2605 6715
rect 2639 6712 2651 6715
rect 2774 6712 2780 6724
rect 2639 6684 2780 6712
rect 2639 6681 2651 6684
rect 2593 6675 2651 6681
rect 2774 6672 2780 6684
rect 2832 6672 2838 6724
rect 2866 6672 2872 6724
rect 2924 6712 2930 6724
rect 3694 6712 3700 6724
rect 2924 6684 3700 6712
rect 2924 6672 2930 6684
rect 3694 6672 3700 6684
rect 3752 6712 3758 6724
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 3752 6684 3801 6712
rect 3752 6672 3758 6684
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3789 6675 3847 6681
rect 6914 6672 6920 6724
rect 6972 6712 6978 6724
rect 9140 6712 9168 6752
rect 6972 6684 9168 6712
rect 6972 6672 6978 6684
rect 9950 6672 9956 6724
rect 10008 6712 10014 6724
rect 10686 6721 10692 6724
rect 10673 6715 10692 6721
rect 10008 6684 10640 6712
rect 10008 6672 10014 6684
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 3050 6644 3056 6656
rect 3011 6616 3056 6644
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 7466 6644 7472 6656
rect 7427 6616 7472 6644
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 8294 6644 8300 6656
rect 7984 6616 8300 6644
rect 7984 6604 7990 6616
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 8628 6616 9137 6644
rect 8628 6604 8634 6616
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 9125 6607 9183 6613
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 10505 6647 10563 6653
rect 10505 6644 10517 6647
rect 10284 6616 10517 6644
rect 10284 6604 10290 6616
rect 10505 6613 10517 6616
rect 10551 6613 10563 6647
rect 10612 6644 10640 6684
rect 10673 6681 10685 6715
rect 10673 6675 10692 6681
rect 10686 6672 10692 6675
rect 10744 6672 10750 6724
rect 10873 6715 10931 6721
rect 10873 6681 10885 6715
rect 10919 6681 10931 6715
rect 10980 6712 11008 6752
rect 12084 6724 12112 6752
rect 13078 6740 13084 6792
rect 13136 6740 13142 6792
rect 13262 6780 13268 6792
rect 13188 6752 13268 6780
rect 11793 6715 11851 6721
rect 11793 6712 11805 6715
rect 10980 6684 11805 6712
rect 10873 6675 10931 6681
rect 11793 6681 11805 6684
rect 11839 6681 11851 6715
rect 11793 6675 11851 6681
rect 10888 6644 10916 6675
rect 12066 6672 12072 6724
rect 12124 6672 12130 6724
rect 12434 6672 12440 6724
rect 12492 6712 12498 6724
rect 12713 6715 12771 6721
rect 12713 6712 12725 6715
rect 12492 6684 12725 6712
rect 12492 6672 12498 6684
rect 12713 6681 12725 6684
rect 12759 6681 12771 6715
rect 12713 6675 12771 6681
rect 10612 6616 10916 6644
rect 10505 6607 10563 6613
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11333 6647 11391 6653
rect 11333 6644 11345 6647
rect 11204 6616 11345 6644
rect 11204 6604 11210 6616
rect 11333 6613 11345 6616
rect 11379 6613 11391 6647
rect 11333 6607 11391 6613
rect 11701 6647 11759 6653
rect 11701 6613 11713 6647
rect 11747 6644 11759 6647
rect 13188 6644 13216 6752
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 11747 6616 13216 6644
rect 13265 6647 13323 6653
rect 11747 6613 11759 6616
rect 11701 6607 11759 6613
rect 13265 6613 13277 6647
rect 13311 6644 13323 6647
rect 13372 6644 13400 6820
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 13780 6820 14749 6848
rect 13780 6808 13786 6820
rect 14737 6817 14749 6820
rect 14783 6817 14795 6851
rect 14737 6811 14795 6817
rect 15289 6851 15347 6857
rect 15289 6817 15301 6851
rect 15335 6848 15347 6851
rect 16298 6848 16304 6860
rect 15335 6820 16304 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 19702 6848 19708 6860
rect 17420 6820 19708 6848
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 15102 6780 15108 6792
rect 13495 6752 15108 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 17420 6789 17448 6820
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 19904 6848 19932 6879
rect 20714 6876 20720 6928
rect 20772 6916 20778 6928
rect 31018 6916 31024 6928
rect 20772 6888 31024 6916
rect 20772 6876 20778 6888
rect 31018 6876 31024 6888
rect 31076 6876 31082 6928
rect 21358 6848 21364 6860
rect 19904 6820 21364 6848
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 22189 6851 22247 6857
rect 22189 6817 22201 6851
rect 22235 6848 22247 6851
rect 23014 6848 23020 6860
rect 22235 6820 23020 6848
rect 22235 6817 22247 6820
rect 22189 6811 22247 6817
rect 23014 6808 23020 6820
rect 23072 6808 23078 6860
rect 24486 6808 24492 6860
rect 24544 6848 24550 6860
rect 31110 6848 31116 6860
rect 24544 6820 31116 6848
rect 24544 6808 24550 6820
rect 31110 6808 31116 6820
rect 31168 6808 31174 6860
rect 42058 6808 42064 6860
rect 42116 6848 42122 6860
rect 42702 6848 42708 6860
rect 42116 6820 42708 6848
rect 42116 6808 42122 6820
rect 42702 6808 42708 6820
rect 42760 6848 42766 6860
rect 43717 6851 43775 6857
rect 43717 6848 43729 6851
rect 42760 6820 43729 6848
rect 42760 6808 42766 6820
rect 43717 6817 43729 6820
rect 43763 6817 43775 6851
rect 43717 6811 43775 6817
rect 17405 6783 17463 6789
rect 17405 6749 17417 6783
rect 17451 6749 17463 6783
rect 17405 6743 17463 6749
rect 18417 6783 18475 6789
rect 18417 6749 18429 6783
rect 18463 6780 18475 6783
rect 18598 6780 18604 6792
rect 18463 6752 18604 6780
rect 18463 6749 18475 6752
rect 18417 6743 18475 6749
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 18230 6672 18236 6724
rect 18288 6712 18294 6724
rect 18708 6712 18736 6743
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 20622 6780 20628 6792
rect 19116 6752 20484 6780
rect 20583 6752 20628 6780
rect 19116 6740 19122 6752
rect 18288 6684 18736 6712
rect 18288 6672 18294 6684
rect 19242 6672 19248 6724
rect 19300 6712 19306 6724
rect 19337 6715 19395 6721
rect 19337 6712 19349 6715
rect 19300 6684 19349 6712
rect 19300 6672 19306 6684
rect 19337 6681 19349 6684
rect 19383 6681 19395 6715
rect 19337 6675 19395 6681
rect 19518 6672 19524 6724
rect 19576 6712 19582 6724
rect 19613 6715 19671 6721
rect 19613 6712 19625 6715
rect 19576 6684 19625 6712
rect 19576 6672 19582 6684
rect 19613 6681 19625 6684
rect 19659 6681 19671 6715
rect 19613 6675 19671 6681
rect 13630 6644 13636 6656
rect 13311 6616 13636 6644
rect 13311 6613 13323 6616
rect 13265 6607 13323 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 14090 6604 14096 6656
rect 14148 6644 14154 6656
rect 14366 6644 14372 6656
rect 14148 6616 14372 6644
rect 14148 6604 14154 6616
rect 14366 6604 14372 6616
rect 14424 6644 14430 6656
rect 15749 6647 15807 6653
rect 15749 6644 15761 6647
rect 14424 6616 15761 6644
rect 14424 6604 14430 6616
rect 15749 6613 15761 6616
rect 15795 6613 15807 6647
rect 16666 6644 16672 6656
rect 16627 6616 16672 6644
rect 15749 6607 15807 6613
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 17218 6644 17224 6656
rect 17179 6616 17224 6644
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 19429 6647 19487 6653
rect 19429 6613 19441 6647
rect 19475 6644 19487 6647
rect 20254 6644 20260 6656
rect 19475 6616 20260 6644
rect 19475 6613 19487 6616
rect 19429 6607 19487 6613
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 20456 6653 20484 6752
rect 20622 6740 20628 6752
rect 20680 6740 20686 6792
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 22465 6783 22523 6789
rect 21591 6752 22094 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 20441 6647 20499 6653
rect 20441 6613 20453 6647
rect 20487 6613 20499 6647
rect 21726 6644 21732 6656
rect 21687 6616 21732 6644
rect 20441 6607 20499 6613
rect 21726 6604 21732 6616
rect 21784 6604 21790 6656
rect 22066 6644 22094 6752
rect 22465 6749 22477 6783
rect 22511 6749 22523 6783
rect 22465 6743 22523 6749
rect 23661 6783 23719 6789
rect 23661 6749 23673 6783
rect 23707 6780 23719 6783
rect 23934 6780 23940 6792
rect 23707 6752 23940 6780
rect 23707 6749 23719 6752
rect 23661 6743 23719 6749
rect 22480 6712 22508 6743
rect 23934 6740 23940 6752
rect 23992 6740 23998 6792
rect 24578 6780 24584 6792
rect 24539 6752 24584 6780
rect 24578 6740 24584 6752
rect 24636 6740 24642 6792
rect 27890 6712 27896 6724
rect 22480 6684 27896 6712
rect 27890 6672 27896 6684
rect 27948 6672 27954 6724
rect 23198 6644 23204 6656
rect 22066 6616 23204 6644
rect 23198 6604 23204 6616
rect 23256 6604 23262 6656
rect 23474 6644 23480 6656
rect 23435 6616 23480 6644
rect 23474 6604 23480 6616
rect 23532 6604 23538 6656
rect 23750 6604 23756 6656
rect 23808 6644 23814 6656
rect 24397 6647 24455 6653
rect 24397 6644 24409 6647
rect 23808 6616 24409 6644
rect 23808 6604 23814 6616
rect 24397 6613 24409 6616
rect 24443 6613 24455 6647
rect 25130 6644 25136 6656
rect 25091 6616 25136 6644
rect 24397 6607 24455 6613
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 25222 6604 25228 6656
rect 25280 6644 25286 6656
rect 25593 6647 25651 6653
rect 25593 6644 25605 6647
rect 25280 6616 25605 6644
rect 25280 6604 25286 6616
rect 25593 6613 25605 6616
rect 25639 6613 25651 6647
rect 25593 6607 25651 6613
rect 1104 6554 44896 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 44896 6554
rect 1104 6480 44896 6502
rect 1857 6443 1915 6449
rect 1857 6409 1869 6443
rect 1903 6440 1915 6443
rect 2498 6440 2504 6452
rect 1903 6412 2504 6440
rect 1903 6409 1915 6412
rect 1857 6403 1915 6409
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 2958 6440 2964 6452
rect 2823 6412 2964 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3878 6440 3884 6452
rect 3839 6412 3884 6440
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 4341 6443 4399 6449
rect 4341 6440 4353 6443
rect 4120 6412 4353 6440
rect 4120 6400 4126 6412
rect 4341 6409 4353 6412
rect 4387 6409 4399 6443
rect 5810 6440 5816 6452
rect 5771 6412 5816 6440
rect 4341 6403 4399 6409
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 7190 6440 7196 6452
rect 7151 6412 7196 6440
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 7984 6412 8309 6440
rect 7984 6400 7990 6412
rect 8297 6409 8309 6412
rect 8343 6409 8355 6443
rect 8297 6403 8355 6409
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 8941 6443 8999 6449
rect 8941 6440 8953 6443
rect 8720 6412 8953 6440
rect 8720 6400 8726 6412
rect 8941 6409 8953 6412
rect 8987 6409 8999 6443
rect 8941 6403 8999 6409
rect 9585 6443 9643 6449
rect 9585 6409 9597 6443
rect 9631 6440 9643 6443
rect 10042 6440 10048 6452
rect 9631 6412 10048 6440
rect 9631 6409 9643 6412
rect 9585 6403 9643 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 11054 6440 11060 6452
rect 10434 6412 11060 6440
rect 2406 6332 2412 6384
rect 2464 6372 2470 6384
rect 8570 6372 8576 6384
rect 2464 6344 8576 6372
rect 2464 6332 2470 6344
rect 8570 6332 8576 6344
rect 8628 6332 8634 6384
rect 10434 6372 10462 6412
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 11882 6440 11888 6452
rect 11164 6412 11888 6440
rect 10060 6344 10462 6372
rect 10060 6316 10088 6344
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 11164 6372 11192 6412
rect 11882 6400 11888 6412
rect 11940 6440 11946 6452
rect 12253 6443 12311 6449
rect 12253 6440 12265 6443
rect 11940 6412 12265 6440
rect 11940 6400 11946 6412
rect 12253 6409 12265 6412
rect 12299 6409 12311 6443
rect 12253 6403 12311 6409
rect 12989 6443 13047 6449
rect 12989 6409 13001 6443
rect 13035 6440 13047 6443
rect 14458 6440 14464 6452
rect 13035 6412 14464 6440
rect 13035 6409 13047 6412
rect 12989 6403 13047 6409
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 14829 6443 14887 6449
rect 14829 6409 14841 6443
rect 14875 6440 14887 6443
rect 15286 6440 15292 6452
rect 14875 6412 15292 6440
rect 14875 6409 14887 6412
rect 14829 6403 14887 6409
rect 15286 6400 15292 6412
rect 15344 6440 15350 6452
rect 15654 6440 15660 6452
rect 15344 6412 15660 6440
rect 15344 6400 15350 6412
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 15933 6443 15991 6449
rect 15933 6409 15945 6443
rect 15979 6440 15991 6443
rect 16114 6440 16120 6452
rect 15979 6412 16120 6440
rect 15979 6409 15991 6412
rect 15933 6403 15991 6409
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 17313 6443 17371 6449
rect 17313 6409 17325 6443
rect 17359 6440 17371 6443
rect 17862 6440 17868 6452
rect 17359 6412 17868 6440
rect 17359 6409 17371 6412
rect 17313 6403 17371 6409
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 20346 6440 20352 6452
rect 18248 6412 20352 6440
rect 10560 6344 10605 6372
rect 10980 6344 11192 6372
rect 11793 6375 11851 6381
rect 10560 6332 10566 6344
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6264 1458 6316
rect 1578 6304 1584 6316
rect 1539 6276 1584 6304
rect 1578 6264 1584 6276
rect 1636 6264 1642 6316
rect 1670 6264 1676 6316
rect 1728 6304 1734 6316
rect 1728 6276 1773 6304
rect 1728 6264 1734 6276
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3237 6307 3295 6313
rect 3237 6304 3249 6307
rect 2832 6276 3249 6304
rect 2832 6264 2838 6276
rect 3237 6273 3249 6276
rect 3283 6273 3295 6307
rect 3237 6267 3295 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6304 6791 6307
rect 7742 6304 7748 6316
rect 6779 6276 7748 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6304 7895 6307
rect 8110 6304 8116 6316
rect 7883 6276 8116 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8481 6307 8539 6313
rect 8481 6273 8493 6307
rect 8527 6304 8539 6307
rect 9030 6304 9036 6316
rect 8527 6276 9036 6304
rect 8527 6273 8539 6276
rect 8481 6267 8539 6273
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9766 6304 9772 6316
rect 9727 6276 9772 6304
rect 9125 6267 9183 6273
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 9140 6236 9168 6267
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 10042 6264 10048 6316
rect 10100 6264 10106 6316
rect 10318 6264 10324 6316
rect 10376 6304 10382 6316
rect 10597 6307 10655 6313
rect 10376 6276 10421 6304
rect 10376 6264 10382 6276
rect 10597 6273 10609 6307
rect 10643 6304 10655 6307
rect 10686 6304 10692 6316
rect 10643 6276 10692 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 10686 6264 10692 6276
rect 10744 6304 10750 6316
rect 10980 6304 11008 6344
rect 11793 6341 11805 6375
rect 11839 6372 11851 6375
rect 12342 6372 12348 6384
rect 11839 6344 12348 6372
rect 11839 6341 11851 6344
rect 11793 6335 11851 6341
rect 12342 6332 12348 6344
rect 12400 6332 12406 6384
rect 14182 6372 14188 6384
rect 12452 6344 14188 6372
rect 10744 6276 11008 6304
rect 10744 6264 10750 6276
rect 11054 6264 11060 6316
rect 11112 6304 11118 6316
rect 11606 6304 11612 6316
rect 11112 6276 11612 6304
rect 11112 6264 11118 6276
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 12452 6313 12480 6344
rect 14182 6332 14188 6344
rect 14240 6332 14246 6384
rect 15102 6332 15108 6384
rect 15160 6372 15166 6384
rect 18141 6375 18199 6381
rect 18141 6372 18153 6375
rect 15160 6344 18153 6372
rect 15160 6332 15166 6344
rect 18141 6341 18153 6344
rect 18187 6341 18199 6375
rect 18141 6335 18199 6341
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6273 12495 6307
rect 12894 6304 12900 6316
rect 12855 6276 12900 6304
rect 12437 6267 12495 6273
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 13078 6304 13084 6316
rect 13039 6276 13084 6304
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13529 6308 13587 6313
rect 13464 6307 13587 6308
rect 13464 6280 13541 6307
rect 13464 6236 13492 6280
rect 13529 6273 13541 6280
rect 13575 6273 13587 6307
rect 13529 6267 13587 6273
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 14642 6304 14648 6316
rect 13771 6276 14648 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 18248 6304 18276 6412
rect 19812 6384 19840 6412
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 31754 6440 31760 6452
rect 20680 6412 31760 6440
rect 20680 6400 20686 6412
rect 31754 6400 31760 6412
rect 31812 6400 31818 6452
rect 19702 6372 19708 6384
rect 19663 6344 19708 6372
rect 19702 6332 19708 6344
rect 19760 6332 19766 6384
rect 19794 6332 19800 6384
rect 19852 6332 19858 6384
rect 21910 6372 21916 6384
rect 21871 6344 21916 6372
rect 21910 6332 21916 6344
rect 21968 6332 21974 6384
rect 23566 6372 23572 6384
rect 23527 6344 23572 6372
rect 23566 6332 23572 6344
rect 23624 6332 23630 6384
rect 24026 6332 24032 6384
rect 24084 6372 24090 6384
rect 24084 6344 35894 6372
rect 24084 6332 24090 6344
rect 17696 6276 18276 6304
rect 18325 6307 18383 6313
rect 4948 6208 9168 6236
rect 12084 6208 13492 6236
rect 4948 6196 4954 6208
rect 2130 6128 2136 6180
rect 2188 6168 2194 6180
rect 5261 6171 5319 6177
rect 5261 6168 5273 6171
rect 2188 6140 5273 6168
rect 2188 6128 2194 6140
rect 5261 6137 5273 6140
rect 5307 6168 5319 6171
rect 8018 6168 8024 6180
rect 5307 6140 8024 6168
rect 5307 6137 5319 6140
rect 5261 6131 5319 6137
rect 8018 6128 8024 6140
rect 8076 6168 8082 6180
rect 12084 6168 12112 6208
rect 8076 6140 12112 6168
rect 8076 6128 8082 6140
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 8110 6060 8116 6112
rect 8168 6100 8174 6112
rect 10226 6100 10232 6112
rect 8168 6072 10232 6100
rect 8168 6060 8174 6072
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10321 6103 10379 6109
rect 10321 6069 10333 6103
rect 10367 6100 10379 6103
rect 11054 6100 11060 6112
rect 10367 6072 11060 6100
rect 10367 6069 10379 6072
rect 10321 6063 10379 6069
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 13464 6100 13492 6208
rect 13633 6239 13691 6245
rect 13633 6205 13645 6239
rect 13679 6236 13691 6239
rect 15378 6236 15384 6248
rect 13679 6208 14596 6236
rect 15339 6208 15384 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 14182 6168 14188 6180
rect 14143 6140 14188 6168
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 13814 6100 13820 6112
rect 13464 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 14568 6100 14596 6208
rect 15378 6196 15384 6208
rect 15436 6196 15442 6248
rect 17696 6236 17724 6276
rect 18325 6273 18337 6307
rect 18371 6304 18383 6307
rect 18598 6304 18604 6316
rect 18371 6276 18604 6304
rect 18371 6273 18383 6276
rect 18325 6267 18383 6273
rect 18598 6264 18604 6276
rect 18656 6264 18662 6316
rect 19613 6307 19671 6313
rect 19613 6273 19625 6307
rect 19659 6304 19671 6307
rect 19886 6304 19892 6316
rect 19659 6276 19892 6304
rect 19659 6273 19671 6276
rect 19613 6267 19671 6273
rect 19886 6264 19892 6276
rect 19944 6304 19950 6316
rect 23290 6304 23296 6316
rect 19944 6276 23296 6304
rect 19944 6264 19950 6276
rect 23290 6264 23296 6276
rect 23348 6264 23354 6316
rect 15856 6208 17724 6236
rect 14642 6128 14648 6180
rect 14700 6168 14706 6180
rect 15856 6168 15884 6208
rect 17862 6196 17868 6248
rect 17920 6236 17926 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17920 6208 18061 6236
rect 17920 6196 17926 6208
rect 18049 6205 18061 6208
rect 18095 6236 18107 6239
rect 19150 6236 19156 6248
rect 18095 6208 19156 6236
rect 18095 6205 18107 6208
rect 18049 6199 18107 6205
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 19797 6239 19855 6245
rect 19797 6205 19809 6239
rect 19843 6236 19855 6239
rect 20070 6236 20076 6248
rect 19843 6208 20076 6236
rect 19843 6205 19855 6208
rect 19797 6199 19855 6205
rect 20070 6196 20076 6208
rect 20128 6196 20134 6248
rect 20809 6239 20867 6245
rect 20809 6205 20821 6239
rect 20855 6236 20867 6239
rect 21450 6236 21456 6248
rect 20855 6208 21456 6236
rect 20855 6205 20867 6208
rect 20809 6199 20867 6205
rect 21450 6196 21456 6208
rect 21508 6236 21514 6248
rect 21634 6236 21640 6248
rect 21508 6208 21640 6236
rect 21508 6196 21514 6208
rect 21634 6196 21640 6208
rect 21692 6196 21698 6248
rect 29822 6236 29828 6248
rect 22066 6208 29828 6236
rect 14700 6140 15884 6168
rect 14700 6128 14706 6140
rect 15930 6128 15936 6180
rect 15988 6168 15994 6180
rect 16761 6171 16819 6177
rect 16761 6168 16773 6171
rect 15988 6140 16773 6168
rect 15988 6128 15994 6140
rect 16761 6137 16773 6140
rect 16807 6168 16819 6171
rect 18601 6171 18659 6177
rect 16807 6140 17908 6168
rect 16807 6137 16819 6140
rect 16761 6131 16819 6137
rect 17586 6100 17592 6112
rect 14568 6072 17592 6100
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 17880 6100 17908 6140
rect 18601 6137 18613 6171
rect 18647 6168 18659 6171
rect 19978 6168 19984 6180
rect 18647 6140 19984 6168
rect 18647 6137 18659 6140
rect 18601 6131 18659 6137
rect 19978 6128 19984 6140
rect 20036 6128 20042 6180
rect 20165 6171 20223 6177
rect 20165 6137 20177 6171
rect 20211 6168 20223 6171
rect 22066 6168 22094 6208
rect 29822 6196 29828 6208
rect 29880 6196 29886 6248
rect 20211 6140 22094 6168
rect 24121 6171 24179 6177
rect 20211 6137 20223 6140
rect 20165 6131 20223 6137
rect 24121 6137 24133 6171
rect 24167 6168 24179 6171
rect 24486 6168 24492 6180
rect 24167 6140 24492 6168
rect 24167 6137 24179 6140
rect 24121 6131 24179 6137
rect 24486 6128 24492 6140
rect 24544 6128 24550 6180
rect 35866 6168 35894 6344
rect 42794 6168 42800 6180
rect 35866 6140 42800 6168
rect 42794 6128 42800 6140
rect 42852 6128 42858 6180
rect 20714 6100 20720 6112
rect 17880 6072 20720 6100
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 21082 6060 21088 6112
rect 21140 6100 21146 6112
rect 22373 6103 22431 6109
rect 22373 6100 22385 6103
rect 21140 6072 22385 6100
rect 21140 6060 21146 6072
rect 22373 6069 22385 6072
rect 22419 6069 22431 6103
rect 22922 6100 22928 6112
rect 22883 6072 22928 6100
rect 22373 6063 22431 6069
rect 22922 6060 22928 6072
rect 22980 6060 22986 6112
rect 24578 6100 24584 6112
rect 24539 6072 24584 6100
rect 24578 6060 24584 6072
rect 24636 6060 24642 6112
rect 25225 6103 25283 6109
rect 25225 6069 25237 6103
rect 25271 6100 25283 6103
rect 25406 6100 25412 6112
rect 25271 6072 25412 6100
rect 25271 6069 25283 6072
rect 25225 6063 25283 6069
rect 25406 6060 25412 6072
rect 25464 6060 25470 6112
rect 25682 6100 25688 6112
rect 25643 6072 25688 6100
rect 25682 6060 25688 6072
rect 25740 6060 25746 6112
rect 26234 6100 26240 6112
rect 26195 6072 26240 6100
rect 26234 6060 26240 6072
rect 26292 6060 26298 6112
rect 42978 6060 42984 6112
rect 43036 6100 43042 6112
rect 43073 6103 43131 6109
rect 43073 6100 43085 6103
rect 43036 6072 43085 6100
rect 43036 6060 43042 6072
rect 43073 6069 43085 6072
rect 43119 6100 43131 6103
rect 43162 6100 43168 6112
rect 43119 6072 43168 6100
rect 43119 6069 43131 6072
rect 43073 6063 43131 6069
rect 43162 6060 43168 6072
rect 43220 6060 43226 6112
rect 43625 6103 43683 6109
rect 43625 6069 43637 6103
rect 43671 6100 43683 6103
rect 43806 6100 43812 6112
rect 43671 6072 43812 6100
rect 43671 6069 43683 6072
rect 43625 6063 43683 6069
rect 43806 6060 43812 6072
rect 43864 6060 43870 6112
rect 44174 6100 44180 6112
rect 44135 6072 44180 6100
rect 44174 6060 44180 6072
rect 44232 6060 44238 6112
rect 1104 6010 44896 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 44896 6010
rect 1104 5936 44896 5958
rect 1394 5896 1400 5908
rect 1355 5868 1400 5896
rect 1394 5856 1400 5868
rect 1452 5856 1458 5908
rect 2685 5899 2743 5905
rect 2685 5865 2697 5899
rect 2731 5896 2743 5899
rect 3050 5896 3056 5908
rect 2731 5868 3056 5896
rect 2731 5865 2743 5868
rect 2685 5859 2743 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 3752 5868 3801 5896
rect 3752 5856 3758 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 3789 5859 3847 5865
rect 6454 5856 6460 5908
rect 6512 5896 6518 5908
rect 6641 5899 6699 5905
rect 6641 5896 6653 5899
rect 6512 5868 6653 5896
rect 6512 5856 6518 5868
rect 6641 5865 6653 5868
rect 6687 5865 6699 5899
rect 6641 5859 6699 5865
rect 7837 5899 7895 5905
rect 7837 5865 7849 5899
rect 7883 5896 7895 5899
rect 8202 5896 8208 5908
rect 7883 5868 8208 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 8754 5896 8760 5908
rect 8435 5868 8760 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 9217 5899 9275 5905
rect 9217 5865 9229 5899
rect 9263 5896 9275 5899
rect 9398 5896 9404 5908
rect 9263 5868 9404 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 10594 5896 10600 5908
rect 10555 5868 10600 5896
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 11241 5899 11299 5905
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11330 5896 11336 5908
rect 11287 5868 11336 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 11790 5856 11796 5908
rect 11848 5896 11854 5908
rect 12250 5896 12256 5908
rect 11848 5868 12256 5896
rect 11848 5856 11854 5868
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 13538 5896 13544 5908
rect 12406 5868 12940 5896
rect 13499 5868 13544 5896
rect 2133 5831 2191 5837
rect 2133 5797 2145 5831
rect 2179 5828 2191 5831
rect 2866 5828 2872 5840
rect 2179 5800 2872 5828
rect 2179 5797 2191 5800
rect 2133 5791 2191 5797
rect 2866 5788 2872 5800
rect 2924 5788 2930 5840
rect 2958 5788 2964 5840
rect 3016 5828 3022 5840
rect 3145 5831 3203 5837
rect 3145 5828 3157 5831
rect 3016 5800 3157 5828
rect 3016 5788 3022 5800
rect 3145 5797 3157 5800
rect 3191 5797 3203 5831
rect 3145 5791 3203 5797
rect 8266 5800 10824 5828
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1544 5664 1593 5692
rect 1544 5652 1550 5664
rect 1581 5661 1593 5664
rect 1627 5692 1639 5695
rect 4062 5692 4068 5704
rect 1627 5664 4068 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4893 5627 4951 5633
rect 4893 5593 4905 5627
rect 4939 5624 4951 5627
rect 5074 5624 5080 5636
rect 4939 5596 5080 5624
rect 4939 5593 4951 5596
rect 4893 5587 4951 5593
rect 5074 5584 5080 5596
rect 5132 5624 5138 5636
rect 5718 5624 5724 5636
rect 5132 5596 5724 5624
rect 5132 5584 5138 5596
rect 5718 5584 5724 5596
rect 5776 5584 5782 5636
rect 7285 5627 7343 5633
rect 7285 5593 7297 5627
rect 7331 5624 7343 5627
rect 7374 5624 7380 5636
rect 7331 5596 7380 5624
rect 7331 5593 7343 5596
rect 7285 5587 7343 5593
rect 7374 5584 7380 5596
rect 7432 5624 7438 5636
rect 8018 5624 8024 5636
rect 7432 5596 8024 5624
rect 7432 5584 7438 5596
rect 8018 5584 8024 5596
rect 8076 5624 8082 5636
rect 8266 5624 8294 5800
rect 10796 5760 10824 5800
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 12066 5828 12072 5840
rect 11112 5800 12072 5828
rect 11112 5788 11118 5800
rect 12066 5788 12072 5800
rect 12124 5828 12130 5840
rect 12406 5828 12434 5868
rect 12124 5800 12434 5828
rect 12124 5788 12130 5800
rect 10796 5732 11284 5760
rect 8478 5652 8484 5704
rect 8536 5692 8542 5704
rect 9861 5695 9919 5701
rect 9861 5692 9873 5695
rect 8536 5664 9873 5692
rect 8536 5652 8542 5664
rect 9861 5661 9873 5664
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 10284 5664 10425 5692
rect 10284 5652 10290 5664
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 8076 5596 8294 5624
rect 10428 5624 10456 5655
rect 10594 5652 10600 5704
rect 10652 5692 10658 5704
rect 11256 5701 11284 5732
rect 11057 5695 11115 5701
rect 11057 5692 11069 5695
rect 10652 5664 10697 5692
rect 10888 5664 11069 5692
rect 10652 5652 10658 5664
rect 10888 5624 10916 5664
rect 11057 5661 11069 5664
rect 11103 5692 11115 5695
rect 11241 5695 11299 5701
rect 11103 5664 11192 5692
rect 11103 5661 11115 5664
rect 11057 5655 11115 5661
rect 10428 5596 10916 5624
rect 11164 5624 11192 5664
rect 11241 5661 11253 5695
rect 11287 5692 11299 5695
rect 12342 5692 12348 5704
rect 11287 5664 12348 5692
rect 11287 5661 11299 5664
rect 11241 5655 11299 5661
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 12912 5692 12940 5868
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 14829 5899 14887 5905
rect 14829 5865 14841 5899
rect 14875 5896 14887 5899
rect 15010 5896 15016 5908
rect 14875 5868 15016 5896
rect 14875 5865 14887 5868
rect 14829 5859 14887 5865
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 16390 5896 16396 5908
rect 16351 5868 16396 5896
rect 16390 5856 16396 5868
rect 16448 5856 16454 5908
rect 16574 5856 16580 5908
rect 16632 5896 16638 5908
rect 16945 5899 17003 5905
rect 16945 5896 16957 5899
rect 16632 5868 16957 5896
rect 16632 5856 16638 5868
rect 16945 5865 16957 5868
rect 16991 5865 17003 5899
rect 16945 5859 17003 5865
rect 18141 5899 18199 5905
rect 18141 5865 18153 5899
rect 18187 5896 18199 5899
rect 18322 5896 18328 5908
rect 18187 5868 18328 5896
rect 18187 5865 18199 5868
rect 18141 5859 18199 5865
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 18693 5899 18751 5905
rect 18693 5865 18705 5899
rect 18739 5896 18751 5899
rect 18782 5896 18788 5908
rect 18739 5868 18788 5896
rect 18739 5865 18751 5868
rect 18693 5859 18751 5865
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 19337 5899 19395 5905
rect 19337 5896 19349 5899
rect 19300 5868 19349 5896
rect 19300 5856 19306 5868
rect 19337 5865 19349 5868
rect 19383 5865 19395 5899
rect 19886 5896 19892 5908
rect 19847 5868 19892 5896
rect 19337 5859 19395 5865
rect 19886 5856 19892 5868
rect 19944 5856 19950 5908
rect 20993 5899 21051 5905
rect 20993 5865 21005 5899
rect 21039 5896 21051 5899
rect 21174 5896 21180 5908
rect 21039 5868 21180 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 21174 5856 21180 5868
rect 21232 5856 21238 5908
rect 23106 5896 23112 5908
rect 23067 5868 23112 5896
rect 23106 5856 23112 5868
rect 23164 5856 23170 5908
rect 23290 5856 23296 5908
rect 23348 5896 23354 5908
rect 26605 5899 26663 5905
rect 26605 5896 26617 5899
rect 23348 5868 26617 5896
rect 23348 5856 23354 5868
rect 26605 5865 26617 5868
rect 26651 5865 26663 5899
rect 27154 5896 27160 5908
rect 27115 5868 27160 5896
rect 26605 5859 26663 5865
rect 27154 5856 27160 5868
rect 27212 5856 27218 5908
rect 27798 5896 27804 5908
rect 27759 5868 27804 5896
rect 27798 5856 27804 5868
rect 27856 5856 27862 5908
rect 27890 5856 27896 5908
rect 27948 5896 27954 5908
rect 34514 5896 34520 5908
rect 27948 5868 34520 5896
rect 27948 5856 27954 5868
rect 34514 5856 34520 5868
rect 34572 5856 34578 5908
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 13872 5800 18092 5828
rect 13872 5788 13878 5800
rect 12989 5763 13047 5769
rect 12989 5729 13001 5763
rect 13035 5760 13047 5763
rect 13170 5760 13176 5772
rect 13035 5732 13176 5760
rect 13035 5729 13047 5732
rect 12989 5723 13047 5729
rect 13170 5720 13176 5732
rect 13228 5760 13234 5772
rect 14185 5763 14243 5769
rect 14185 5760 14197 5763
rect 13228 5732 14197 5760
rect 13228 5720 13234 5732
rect 14185 5729 14197 5732
rect 14231 5729 14243 5763
rect 15286 5760 15292 5772
rect 14185 5723 14243 5729
rect 14292 5732 15292 5760
rect 14292 5692 14320 5732
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 16022 5720 16028 5772
rect 16080 5760 16086 5772
rect 18064 5760 18092 5800
rect 18966 5788 18972 5840
rect 19024 5828 19030 5840
rect 26053 5831 26111 5837
rect 26053 5828 26065 5831
rect 19024 5800 26065 5828
rect 19024 5788 19030 5800
rect 26053 5797 26065 5800
rect 26099 5797 26111 5831
rect 26053 5791 26111 5797
rect 20346 5760 20352 5772
rect 16080 5732 18000 5760
rect 18064 5732 20352 5760
rect 16080 5720 16086 5732
rect 12912 5664 14320 5692
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5692 14519 5695
rect 15654 5692 15660 5704
rect 14507 5664 15660 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 17034 5692 17040 5704
rect 16816 5664 17040 5692
rect 16816 5652 16822 5664
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 17586 5692 17592 5704
rect 17547 5664 17592 5692
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 17972 5692 18000 5732
rect 20346 5720 20352 5732
rect 20404 5720 20410 5772
rect 23198 5720 23204 5772
rect 23256 5760 23262 5772
rect 24949 5763 25007 5769
rect 24949 5760 24961 5763
rect 23256 5732 24961 5760
rect 23256 5720 23262 5732
rect 24949 5729 24961 5732
rect 24995 5729 25007 5763
rect 24949 5723 25007 5729
rect 24578 5692 24584 5704
rect 17972 5664 24584 5692
rect 24578 5652 24584 5664
rect 24636 5652 24642 5704
rect 42702 5652 42708 5704
rect 42760 5692 42766 5704
rect 43901 5695 43959 5701
rect 43901 5692 43913 5695
rect 42760 5664 43913 5692
rect 42760 5652 42766 5664
rect 43901 5661 43913 5664
rect 43947 5661 43959 5695
rect 43901 5655 43959 5661
rect 11606 5624 11612 5636
rect 11164 5596 11612 5624
rect 8076 5584 8082 5596
rect 11606 5584 11612 5596
rect 11664 5584 11670 5636
rect 14366 5624 14372 5636
rect 14327 5596 14372 5624
rect 14366 5584 14372 5596
rect 14424 5584 14430 5636
rect 15841 5627 15899 5633
rect 15841 5624 15853 5627
rect 14476 5596 15853 5624
rect 14476 5568 14504 5596
rect 15841 5593 15853 5596
rect 15887 5624 15899 5627
rect 16117 5627 16175 5633
rect 15887 5596 16068 5624
rect 15887 5593 15899 5596
rect 15841 5587 15899 5593
rect 5445 5559 5503 5565
rect 5445 5525 5457 5559
rect 5491 5556 5503 5559
rect 5626 5556 5632 5568
rect 5491 5528 5632 5556
rect 5491 5525 5503 5528
rect 5445 5519 5503 5525
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 5902 5556 5908 5568
rect 5863 5528 5908 5556
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 6086 5516 6092 5568
rect 6144 5556 6150 5568
rect 7006 5556 7012 5568
rect 6144 5528 7012 5556
rect 6144 5516 6150 5528
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 9766 5556 9772 5568
rect 9723 5528 9772 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 11790 5556 11796 5568
rect 11751 5528 11796 5556
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 11882 5516 11888 5568
rect 11940 5556 11946 5568
rect 13081 5559 13139 5565
rect 13081 5556 13093 5559
rect 11940 5528 13093 5556
rect 11940 5516 11946 5528
rect 13081 5525 13093 5528
rect 13127 5525 13139 5559
rect 13081 5519 13139 5525
rect 13170 5516 13176 5568
rect 13228 5556 13234 5568
rect 13228 5528 13273 5556
rect 13228 5516 13234 5528
rect 14458 5516 14464 5568
rect 14516 5516 14522 5568
rect 15930 5556 15936 5568
rect 15891 5528 15936 5556
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 16040 5556 16068 5596
rect 16117 5593 16129 5627
rect 16163 5624 16175 5627
rect 19334 5624 19340 5636
rect 16163 5596 19340 5624
rect 16163 5593 16175 5596
rect 16117 5587 16175 5593
rect 19334 5584 19340 5596
rect 19392 5584 19398 5636
rect 22186 5584 22192 5636
rect 22244 5624 22250 5636
rect 22557 5627 22615 5633
rect 22557 5624 22569 5627
rect 22244 5596 22569 5624
rect 22244 5584 22250 5596
rect 22557 5593 22569 5596
rect 22603 5593 22615 5627
rect 22557 5587 22615 5593
rect 23014 5584 23020 5636
rect 23072 5624 23078 5636
rect 24397 5627 24455 5633
rect 24397 5624 24409 5627
rect 23072 5596 24409 5624
rect 23072 5584 23078 5596
rect 24397 5593 24409 5596
rect 24443 5593 24455 5627
rect 24397 5587 24455 5593
rect 18506 5556 18512 5568
rect 16040 5528 18512 5556
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 21545 5559 21603 5565
rect 21545 5525 21557 5559
rect 21591 5556 21603 5559
rect 22002 5556 22008 5568
rect 21591 5528 22008 5556
rect 21591 5525 21603 5528
rect 21545 5519 21603 5525
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 22097 5559 22155 5565
rect 22097 5525 22109 5559
rect 22143 5556 22155 5559
rect 22462 5556 22468 5568
rect 22143 5528 22468 5556
rect 22143 5525 22155 5528
rect 22097 5519 22155 5525
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 23658 5556 23664 5568
rect 23619 5528 23664 5556
rect 23658 5516 23664 5528
rect 23716 5516 23722 5568
rect 24854 5516 24860 5568
rect 24912 5556 24918 5568
rect 25501 5559 25559 5565
rect 25501 5556 25513 5559
rect 24912 5528 25513 5556
rect 24912 5516 24918 5528
rect 25501 5525 25513 5528
rect 25547 5525 25559 5559
rect 25501 5519 25559 5525
rect 26142 5516 26148 5568
rect 26200 5556 26206 5568
rect 30190 5556 30196 5568
rect 26200 5528 30196 5556
rect 26200 5516 26206 5528
rect 30190 5516 30196 5528
rect 30248 5516 30254 5568
rect 41690 5556 41696 5568
rect 41651 5528 41696 5556
rect 41690 5516 41696 5528
rect 41748 5516 41754 5568
rect 42150 5516 42156 5568
rect 42208 5556 42214 5568
rect 42245 5559 42303 5565
rect 42245 5556 42257 5559
rect 42208 5528 42257 5556
rect 42208 5516 42214 5528
rect 42245 5525 42257 5528
rect 42291 5556 42303 5559
rect 42334 5556 42340 5568
rect 42291 5528 42340 5556
rect 42291 5525 42303 5528
rect 42245 5519 42303 5525
rect 42334 5516 42340 5528
rect 42392 5516 42398 5568
rect 42886 5556 42892 5568
rect 42847 5528 42892 5556
rect 42886 5516 42892 5528
rect 42944 5516 42950 5568
rect 43441 5559 43499 5565
rect 43441 5525 43453 5559
rect 43487 5556 43499 5559
rect 43530 5556 43536 5568
rect 43487 5528 43536 5556
rect 43487 5525 43499 5528
rect 43441 5519 43499 5525
rect 43530 5516 43536 5528
rect 43588 5516 43594 5568
rect 44085 5559 44143 5565
rect 44085 5525 44097 5559
rect 44131 5556 44143 5559
rect 45094 5556 45100 5568
rect 44131 5528 45100 5556
rect 44131 5525 44143 5528
rect 44085 5519 44143 5525
rect 45094 5516 45100 5528
rect 45152 5516 45158 5568
rect 1104 5466 44896 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 44896 5466
rect 1104 5392 44896 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 1670 5352 1676 5364
rect 1627 5324 1676 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 1670 5312 1676 5324
rect 1728 5312 1734 5364
rect 2130 5352 2136 5364
rect 2091 5324 2136 5352
rect 2130 5312 2136 5324
rect 2188 5312 2194 5364
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 5902 5352 5908 5364
rect 4203 5324 5908 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 6362 5352 6368 5364
rect 6323 5324 6368 5352
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 8018 5352 8024 5364
rect 7979 5324 8024 5352
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 9858 5352 9864 5364
rect 9815 5324 9864 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 10134 5312 10140 5364
rect 10192 5352 10198 5364
rect 10321 5355 10379 5361
rect 10321 5352 10333 5355
rect 10192 5324 10333 5352
rect 10192 5312 10198 5324
rect 10321 5321 10333 5324
rect 10367 5321 10379 5355
rect 10321 5315 10379 5321
rect 10778 5312 10784 5364
rect 10836 5352 10842 5364
rect 11517 5355 11575 5361
rect 11517 5352 11529 5355
rect 10836 5324 11529 5352
rect 10836 5312 10842 5324
rect 11517 5321 11529 5324
rect 11563 5321 11575 5355
rect 11517 5315 11575 5321
rect 842 5244 848 5296
rect 900 5284 906 5296
rect 2777 5287 2835 5293
rect 2777 5284 2789 5287
rect 900 5256 2789 5284
rect 900 5244 906 5256
rect 2777 5253 2789 5256
rect 2823 5253 2835 5287
rect 2777 5247 2835 5253
rect 4062 5244 4068 5296
rect 4120 5284 4126 5296
rect 5442 5284 5448 5296
rect 4120 5256 5448 5284
rect 4120 5244 4126 5256
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 7006 5244 7012 5296
rect 7064 5284 7070 5296
rect 8573 5287 8631 5293
rect 8573 5284 8585 5287
rect 7064 5256 8585 5284
rect 7064 5244 7070 5256
rect 8573 5253 8585 5256
rect 8619 5284 8631 5287
rect 10226 5284 10232 5296
rect 8619 5256 10232 5284
rect 8619 5253 8631 5256
rect 8573 5247 8631 5253
rect 10226 5244 10232 5256
rect 10284 5244 10290 5296
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5176 1458 5228
rect 8386 5176 8392 5228
rect 8444 5216 8450 5228
rect 9585 5219 9643 5225
rect 9585 5216 9597 5219
rect 8444 5188 9597 5216
rect 8444 5176 8450 5188
rect 9585 5185 9597 5188
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 8846 5148 8852 5160
rect 4028 5120 8852 5148
rect 4028 5108 4034 5120
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 10778 5148 10784 5160
rect 10739 5120 10784 5148
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 11532 5148 11560 5315
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 15565 5355 15623 5361
rect 11848 5324 15516 5352
rect 11848 5312 11854 5324
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 14461 5287 14519 5293
rect 14461 5284 14473 5287
rect 12308 5256 14473 5284
rect 12308 5244 12314 5256
rect 14461 5253 14473 5256
rect 14507 5253 14519 5287
rect 15488 5284 15516 5324
rect 15565 5321 15577 5355
rect 15611 5352 15623 5355
rect 15654 5352 15660 5364
rect 15611 5324 15660 5352
rect 15611 5321 15623 5324
rect 15565 5315 15623 5321
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 16114 5352 16120 5364
rect 16075 5324 16120 5352
rect 16114 5312 16120 5324
rect 16172 5312 16178 5364
rect 16761 5355 16819 5361
rect 16761 5321 16773 5355
rect 16807 5352 16819 5355
rect 16850 5352 16856 5364
rect 16807 5324 16856 5352
rect 16807 5321 16819 5324
rect 16761 5315 16819 5321
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17862 5352 17868 5364
rect 17823 5324 17868 5352
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 18414 5352 18420 5364
rect 18196 5324 18420 5352
rect 18196 5312 18202 5324
rect 18414 5312 18420 5324
rect 18472 5352 18478 5364
rect 18877 5355 18935 5361
rect 18877 5352 18889 5355
rect 18472 5324 18889 5352
rect 18472 5312 18478 5324
rect 18877 5321 18889 5324
rect 18923 5321 18935 5355
rect 18877 5315 18935 5321
rect 20622 5312 20628 5364
rect 20680 5352 20686 5364
rect 23658 5352 23664 5364
rect 20680 5324 23664 5352
rect 20680 5312 20686 5324
rect 23658 5312 23664 5324
rect 23716 5312 23722 5364
rect 28074 5352 28080 5364
rect 28035 5324 28080 5352
rect 28074 5312 28080 5324
rect 28132 5352 28138 5364
rect 28258 5352 28264 5364
rect 28132 5324 28264 5352
rect 28132 5312 28138 5324
rect 28258 5312 28264 5324
rect 28316 5312 28322 5364
rect 41414 5352 41420 5364
rect 41375 5324 41420 5352
rect 41414 5312 41420 5324
rect 41472 5312 41478 5364
rect 16666 5284 16672 5296
rect 15488 5256 16672 5284
rect 14461 5247 14519 5253
rect 16666 5244 16672 5256
rect 16724 5244 16730 5296
rect 18322 5284 18328 5296
rect 18283 5256 18328 5284
rect 18322 5244 18328 5256
rect 18380 5244 18386 5296
rect 19518 5284 19524 5296
rect 19431 5256 19524 5284
rect 19518 5244 19524 5256
rect 19576 5284 19582 5296
rect 26602 5284 26608 5296
rect 19576 5256 26608 5284
rect 19576 5244 19582 5256
rect 26602 5244 26608 5256
rect 26660 5244 26666 5296
rect 42242 5244 42248 5296
rect 42300 5284 42306 5296
rect 43901 5287 43959 5293
rect 43901 5284 43913 5287
rect 42300 5256 43913 5284
rect 42300 5244 42306 5256
rect 43901 5253 43913 5256
rect 43947 5253 43959 5287
rect 43901 5247 43959 5253
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5216 12495 5219
rect 12710 5216 12716 5228
rect 12483 5188 12716 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 12710 5176 12716 5188
rect 12768 5216 12774 5228
rect 14642 5216 14648 5228
rect 12768 5188 14504 5216
rect 14603 5188 14648 5216
rect 12768 5176 12774 5188
rect 14182 5148 14188 5160
rect 11532 5120 14188 5148
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 14366 5148 14372 5160
rect 14327 5120 14372 5148
rect 14366 5108 14372 5120
rect 14424 5108 14430 5160
rect 14476 5148 14504 5188
rect 14642 5176 14648 5188
rect 14700 5176 14706 5228
rect 16298 5176 16304 5228
rect 16356 5216 16362 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 16356 5188 21833 5216
rect 16356 5176 16362 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 22186 5176 22192 5228
rect 22244 5216 22250 5228
rect 24581 5219 24639 5225
rect 24581 5216 24593 5219
rect 22244 5188 24593 5216
rect 22244 5176 22250 5188
rect 24581 5185 24593 5188
rect 24627 5185 24639 5219
rect 24581 5179 24639 5185
rect 42886 5176 42892 5228
rect 42944 5216 42950 5228
rect 44085 5219 44143 5225
rect 44085 5216 44097 5219
rect 42944 5188 44097 5216
rect 42944 5176 42950 5188
rect 44085 5185 44097 5188
rect 44131 5216 44143 5219
rect 45738 5216 45744 5228
rect 44131 5188 45744 5216
rect 44131 5185 44143 5188
rect 44085 5179 44143 5185
rect 45738 5176 45744 5188
rect 45796 5176 45802 5228
rect 14918 5148 14924 5160
rect 14476 5120 14924 5148
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 15010 5108 15016 5160
rect 15068 5148 15074 5160
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 15068 5120 20545 5148
rect 15068 5108 15074 5120
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 21910 5108 21916 5160
rect 21968 5148 21974 5160
rect 23477 5151 23535 5157
rect 23477 5148 23489 5151
rect 21968 5120 23489 5148
rect 21968 5108 21974 5120
rect 23477 5117 23489 5120
rect 23523 5117 23535 5151
rect 23477 5111 23535 5117
rect 23934 5108 23940 5160
rect 23992 5148 23998 5160
rect 27525 5151 27583 5157
rect 27525 5148 27537 5151
rect 23992 5120 27537 5148
rect 23992 5108 23998 5120
rect 27525 5117 27537 5120
rect 27571 5117 27583 5151
rect 27525 5111 27583 5117
rect 3421 5083 3479 5089
rect 3421 5049 3433 5083
rect 3467 5080 3479 5083
rect 4522 5080 4528 5092
rect 3467 5052 4528 5080
rect 3467 5049 3479 5052
rect 3421 5043 3479 5049
rect 4522 5040 4528 5052
rect 4580 5080 4586 5092
rect 11054 5080 11060 5092
rect 4580 5052 5304 5080
rect 4580 5040 4586 5052
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 5276 5021 5304 5052
rect 5828 5052 11060 5080
rect 5828 5024 5856 5052
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 11330 5040 11336 5092
rect 11388 5080 11394 5092
rect 21085 5083 21143 5089
rect 21085 5080 21097 5083
rect 11388 5052 21097 5080
rect 11388 5040 11394 5052
rect 21085 5049 21097 5052
rect 21131 5049 21143 5083
rect 22922 5080 22928 5092
rect 22883 5052 22928 5080
rect 21085 5043 21143 5049
rect 22922 5040 22928 5052
rect 22980 5040 22986 5092
rect 23382 5040 23388 5092
rect 23440 5080 23446 5092
rect 27890 5080 27896 5092
rect 23440 5052 27896 5080
rect 23440 5040 23446 5052
rect 27890 5040 27896 5052
rect 27948 5040 27954 5092
rect 5261 5015 5319 5021
rect 5261 4981 5273 5015
rect 5307 5012 5319 5015
rect 5442 5012 5448 5024
rect 5307 4984 5448 5012
rect 5307 4981 5319 4984
rect 5261 4975 5319 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 5810 5012 5816 5024
rect 5771 4984 5816 5012
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 7098 4972 7104 5024
rect 7156 5012 7162 5024
rect 7374 5012 7380 5024
rect 7156 4984 7380 5012
rect 7156 4972 7162 4984
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 9030 5012 9036 5024
rect 8991 4984 9036 5012
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 12989 5015 13047 5021
rect 12989 4981 13001 5015
rect 13035 5012 13047 5015
rect 13078 5012 13084 5024
rect 13035 4984 13084 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 13541 5015 13599 5021
rect 13541 4981 13553 5015
rect 13587 5012 13599 5015
rect 13722 5012 13728 5024
rect 13587 4984 13728 5012
rect 13587 4981 13599 4984
rect 13541 4975 13599 4981
rect 13722 4972 13728 4984
rect 13780 4972 13786 5024
rect 14921 5015 14979 5021
rect 14921 4981 14933 5015
rect 14967 5012 14979 5015
rect 15102 5012 15108 5024
rect 14967 4984 15108 5012
rect 14967 4981 14979 4984
rect 14921 4975 14979 4981
rect 15102 4972 15108 4984
rect 15160 4972 15166 5024
rect 17034 4972 17040 5024
rect 17092 5012 17098 5024
rect 17221 5015 17279 5021
rect 17221 5012 17233 5015
rect 17092 4984 17233 5012
rect 17092 4972 17098 4984
rect 17221 4981 17233 4984
rect 17267 4981 17279 5015
rect 17221 4975 17279 4981
rect 17954 4972 17960 5024
rect 18012 5012 18018 5024
rect 19981 5015 20039 5021
rect 19981 5012 19993 5015
rect 18012 4984 19993 5012
rect 18012 4972 18018 4984
rect 19981 4981 19993 4984
rect 20027 4981 20039 5015
rect 19981 4975 20039 4981
rect 22278 4972 22284 5024
rect 22336 5012 22342 5024
rect 22373 5015 22431 5021
rect 22373 5012 22385 5015
rect 22336 4984 22385 5012
rect 22336 4972 22342 4984
rect 22373 4981 22385 4984
rect 22419 4981 22431 5015
rect 24026 5012 24032 5024
rect 23987 4984 24032 5012
rect 22373 4975 22431 4981
rect 24026 4972 24032 4984
rect 24084 4972 24090 5024
rect 24670 4972 24676 5024
rect 24728 5012 24734 5024
rect 25133 5015 25191 5021
rect 25133 5012 25145 5015
rect 24728 4984 25145 5012
rect 24728 4972 24734 4984
rect 25133 4981 25145 4984
rect 25179 4981 25191 5015
rect 25133 4975 25191 4981
rect 25590 4972 25596 5024
rect 25648 5012 25654 5024
rect 25685 5015 25743 5021
rect 25685 5012 25697 5015
rect 25648 4984 25697 5012
rect 25648 4972 25654 4984
rect 25685 4981 25697 4984
rect 25731 4981 25743 5015
rect 26326 5012 26332 5024
rect 26287 4984 26332 5012
rect 25685 4975 25743 4981
rect 26326 4972 26332 4984
rect 26384 4972 26390 5024
rect 26970 5012 26976 5024
rect 26931 4984 26976 5012
rect 26970 4972 26976 4984
rect 27028 4972 27034 5024
rect 42610 5012 42616 5024
rect 42571 4984 42616 5012
rect 42610 4972 42616 4984
rect 42668 4972 42674 5024
rect 43438 5012 43444 5024
rect 43399 4984 43444 5012
rect 43438 4972 43444 4984
rect 43496 4972 43502 5024
rect 1104 4922 44896 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 44896 4922
rect 1104 4848 44896 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 2685 4811 2743 4817
rect 2685 4808 2697 4811
rect 1360 4780 2697 4808
rect 1360 4768 1366 4780
rect 2685 4777 2697 4780
rect 2731 4777 2743 4811
rect 4614 4808 4620 4820
rect 4575 4780 4620 4808
rect 2685 4771 2743 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 5169 4811 5227 4817
rect 5169 4777 5181 4811
rect 5215 4808 5227 4811
rect 8938 4808 8944 4820
rect 5215 4780 8944 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9122 4808 9128 4820
rect 9083 4780 9128 4808
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 9677 4811 9735 4817
rect 9677 4808 9689 4811
rect 9364 4780 9689 4808
rect 9364 4768 9370 4780
rect 9677 4777 9689 4780
rect 9723 4777 9735 4811
rect 10502 4808 10508 4820
rect 10463 4780 10508 4808
rect 9677 4771 9735 4777
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 11238 4808 11244 4820
rect 11199 4780 11244 4808
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 13173 4811 13231 4817
rect 13173 4808 13185 4811
rect 12676 4780 13185 4808
rect 12676 4768 12682 4780
rect 13173 4777 13185 4780
rect 13219 4777 13231 4811
rect 14734 4808 14740 4820
rect 14695 4780 14740 4808
rect 13173 4771 13231 4777
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 14918 4768 14924 4820
rect 14976 4808 14982 4820
rect 15197 4811 15255 4817
rect 15197 4808 15209 4811
rect 14976 4780 15209 4808
rect 14976 4768 14982 4780
rect 15197 4777 15209 4780
rect 15243 4777 15255 4811
rect 16666 4808 16672 4820
rect 16627 4780 16672 4808
rect 15197 4771 15255 4777
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 17310 4768 17316 4820
rect 17368 4808 17374 4820
rect 17773 4811 17831 4817
rect 17773 4808 17785 4811
rect 17368 4780 17785 4808
rect 17368 4768 17374 4780
rect 17773 4777 17785 4780
rect 17819 4777 17831 4811
rect 17773 4771 17831 4777
rect 18230 4768 18236 4820
rect 18288 4808 18294 4820
rect 18325 4811 18383 4817
rect 18325 4808 18337 4811
rect 18288 4780 18337 4808
rect 18288 4768 18294 4780
rect 18325 4777 18337 4780
rect 18371 4777 18383 4811
rect 18325 4771 18383 4777
rect 19337 4811 19395 4817
rect 19337 4777 19349 4811
rect 19383 4808 19395 4811
rect 19978 4808 19984 4820
rect 19383 4780 19984 4808
rect 19383 4777 19395 4780
rect 19337 4771 19395 4777
rect 19978 4768 19984 4780
rect 20036 4768 20042 4820
rect 23658 4808 23664 4820
rect 23619 4780 23664 4808
rect 23658 4768 23664 4780
rect 23716 4768 23722 4820
rect 28810 4808 28816 4820
rect 28771 4780 28816 4808
rect 28810 4768 28816 4780
rect 28868 4768 28874 4820
rect 35894 4768 35900 4820
rect 35952 4808 35958 4820
rect 37918 4808 37924 4820
rect 35952 4780 35997 4808
rect 37879 4780 37924 4808
rect 35952 4768 35958 4780
rect 37918 4768 37924 4780
rect 37976 4768 37982 4820
rect 40770 4808 40776 4820
rect 40731 4780 40776 4808
rect 40770 4768 40776 4780
rect 40828 4768 40834 4820
rect 1578 4740 1584 4752
rect 1539 4712 1584 4740
rect 1578 4700 1584 4712
rect 1636 4700 1642 4752
rect 2225 4743 2283 4749
rect 2225 4709 2237 4743
rect 2271 4740 2283 4743
rect 10410 4740 10416 4752
rect 2271 4712 10416 4740
rect 2271 4709 2283 4712
rect 2225 4703 2283 4709
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 12713 4743 12771 4749
rect 12713 4709 12725 4743
rect 12759 4740 12771 4743
rect 13446 4740 13452 4752
rect 12759 4712 13452 4740
rect 12759 4709 12771 4712
rect 12713 4703 12771 4709
rect 13446 4700 13452 4712
rect 13504 4700 13510 4752
rect 13538 4700 13544 4752
rect 13596 4740 13602 4752
rect 16206 4740 16212 4752
rect 13596 4712 16212 4740
rect 13596 4700 13602 4712
rect 16206 4700 16212 4712
rect 16264 4700 16270 4752
rect 22094 4700 22100 4752
rect 22152 4740 22158 4752
rect 28261 4743 28319 4749
rect 28261 4740 28273 4743
rect 22152 4712 22197 4740
rect 23492 4712 28273 4740
rect 22152 4700 22158 4712
rect 3881 4675 3939 4681
rect 3881 4641 3893 4675
rect 3927 4672 3939 4675
rect 6546 4672 6552 4684
rect 3927 4644 6552 4672
rect 3927 4641 3939 4644
rect 3881 4635 3939 4641
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 6730 4632 6736 4684
rect 6788 4672 6794 4684
rect 7285 4675 7343 4681
rect 7285 4672 7297 4675
rect 6788 4644 7297 4672
rect 6788 4632 6794 4644
rect 7285 4641 7297 4644
rect 7331 4641 7343 4675
rect 7285 4635 7343 4641
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 9490 4672 9496 4684
rect 8435 4644 9496 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 9490 4632 9496 4644
rect 9548 4672 9554 4684
rect 13630 4672 13636 4684
rect 9548 4644 13636 4672
rect 9548 4632 9554 4644
rect 13630 4632 13636 4644
rect 13688 4672 13694 4684
rect 14734 4672 14740 4684
rect 13688 4644 14740 4672
rect 13688 4632 13694 4644
rect 14734 4632 14740 4644
rect 14792 4672 14798 4684
rect 19518 4672 19524 4684
rect 14792 4644 19524 4672
rect 14792 4632 14798 4644
rect 19518 4632 19524 4644
rect 19576 4632 19582 4684
rect 21266 4632 21272 4684
rect 21324 4672 21330 4684
rect 23492 4672 23520 4712
rect 28261 4709 28273 4712
rect 28307 4709 28319 4743
rect 28261 4703 28319 4709
rect 28626 4700 28632 4752
rect 28684 4740 28690 4752
rect 37090 4740 37096 4752
rect 28684 4712 37096 4740
rect 28684 4700 28690 4712
rect 37090 4700 37096 4712
rect 37148 4700 37154 4752
rect 42518 4700 42524 4752
rect 42576 4740 42582 4752
rect 43901 4743 43959 4749
rect 43901 4740 43913 4743
rect 42576 4712 43913 4740
rect 42576 4700 42582 4712
rect 43901 4709 43913 4712
rect 43947 4709 43959 4743
rect 43901 4703 43959 4709
rect 21324 4644 23520 4672
rect 21324 4632 21330 4644
rect 23566 4632 23572 4684
rect 23624 4672 23630 4684
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 23624 4644 24409 4672
rect 23624 4632 23630 4644
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 24397 4635 24455 4641
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 1412 4536 1440 4567
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 2038 4604 2044 4616
rect 1728 4576 2044 4604
rect 1728 4564 1734 4576
rect 2038 4564 2044 4576
rect 2096 4564 2102 4616
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 5684 4576 6837 4604
rect 5684 4564 5690 4576
rect 6825 4573 6837 4576
rect 6871 4604 6883 4607
rect 9030 4604 9036 4616
rect 6871 4576 9036 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 9030 4564 9036 4576
rect 9088 4604 9094 4616
rect 11701 4607 11759 4613
rect 11701 4604 11713 4607
rect 9088 4576 11713 4604
rect 9088 4564 9094 4576
rect 11701 4573 11713 4576
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 14182 4564 14188 4616
rect 14240 4604 14246 4616
rect 15194 4604 15200 4616
rect 14240 4576 15200 4604
rect 14240 4564 14246 4576
rect 15194 4564 15200 4576
rect 15252 4604 15258 4616
rect 16117 4607 16175 4613
rect 16117 4604 16129 4607
rect 15252 4576 16129 4604
rect 15252 4564 15258 4576
rect 16117 4573 16129 4576
rect 16163 4573 16175 4607
rect 16117 4567 16175 4573
rect 3050 4536 3056 4548
rect 1412 4508 3056 4536
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 4706 4496 4712 4548
rect 4764 4536 4770 4548
rect 5721 4539 5779 4545
rect 5721 4536 5733 4539
rect 4764 4508 5733 4536
rect 4764 4496 4770 4508
rect 5721 4505 5733 4508
rect 5767 4536 5779 4539
rect 12710 4536 12716 4548
rect 5767 4508 12716 4536
rect 5767 4505 5779 4508
rect 5721 4499 5779 4505
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 16132 4536 16160 4567
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 19797 4607 19855 4613
rect 19797 4604 19809 4607
rect 16448 4576 19809 4604
rect 16448 4564 16454 4576
rect 19797 4573 19809 4576
rect 19843 4573 19855 4607
rect 19797 4567 19855 4573
rect 20346 4564 20352 4616
rect 20404 4604 20410 4616
rect 26970 4604 26976 4616
rect 20404 4576 26976 4604
rect 20404 4564 20410 4576
rect 26970 4564 26976 4576
rect 27028 4564 27034 4616
rect 39114 4604 39120 4616
rect 27724 4576 39120 4604
rect 17221 4539 17279 4545
rect 17221 4536 17233 4539
rect 16132 4508 17233 4536
rect 17221 4505 17233 4508
rect 17267 4505 17279 4539
rect 17221 4499 17279 4505
rect 18506 4496 18512 4548
rect 18564 4536 18570 4548
rect 20901 4539 20959 4545
rect 20901 4536 20913 4539
rect 18564 4508 20913 4536
rect 18564 4496 18570 4508
rect 20901 4505 20913 4508
rect 20947 4505 20959 4539
rect 22557 4539 22615 4545
rect 22557 4536 22569 4539
rect 20901 4499 20959 4505
rect 22066 4508 22569 4536
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 6273 4471 6331 4477
rect 6273 4468 6285 4471
rect 5500 4440 6285 4468
rect 5500 4428 5506 4440
rect 6273 4437 6285 4440
rect 6319 4468 6331 4471
rect 7926 4468 7932 4480
rect 6319 4440 7932 4468
rect 6319 4437 6331 4440
rect 6273 4431 6331 4437
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 13170 4428 13176 4480
rect 13228 4468 13234 4480
rect 14182 4468 14188 4480
rect 13228 4440 14188 4468
rect 13228 4428 13234 4440
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 19978 4428 19984 4480
rect 20036 4468 20042 4480
rect 20349 4471 20407 4477
rect 20349 4468 20361 4471
rect 20036 4440 20361 4468
rect 20036 4428 20042 4440
rect 20349 4437 20361 4440
rect 20395 4437 20407 4471
rect 21450 4468 21456 4480
rect 21411 4440 21456 4468
rect 20349 4431 20407 4437
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 21542 4428 21548 4480
rect 21600 4468 21606 4480
rect 22066 4468 22094 4508
rect 22557 4505 22569 4508
rect 22603 4505 22615 4539
rect 22557 4499 22615 4505
rect 24118 4496 24124 4548
rect 24176 4536 24182 4548
rect 27724 4536 27752 4576
rect 39114 4564 39120 4576
rect 39172 4564 39178 4616
rect 43162 4604 43168 4616
rect 43123 4576 43168 4604
rect 43162 4564 43168 4576
rect 43220 4564 43226 4616
rect 24176 4508 27752 4536
rect 24176 4496 24182 4508
rect 27890 4496 27896 4548
rect 27948 4536 27954 4548
rect 42153 4539 42211 4545
rect 27948 4508 36584 4536
rect 27948 4496 27954 4508
rect 23106 4468 23112 4480
rect 21600 4440 22094 4468
rect 23067 4440 23112 4468
rect 21600 4428 21606 4440
rect 23106 4428 23112 4440
rect 23164 4428 23170 4480
rect 24946 4468 24952 4480
rect 24907 4440 24952 4468
rect 24946 4428 24952 4440
rect 25004 4428 25010 4480
rect 25038 4428 25044 4480
rect 25096 4468 25102 4480
rect 25501 4471 25559 4477
rect 25501 4468 25513 4471
rect 25096 4440 25513 4468
rect 25096 4428 25102 4440
rect 25501 4437 25513 4440
rect 25547 4437 25559 4471
rect 25501 4431 25559 4437
rect 26145 4471 26203 4477
rect 26145 4437 26157 4471
rect 26191 4468 26203 4471
rect 26418 4468 26424 4480
rect 26191 4440 26424 4468
rect 26191 4437 26203 4440
rect 26145 4431 26203 4437
rect 26418 4428 26424 4440
rect 26476 4428 26482 4480
rect 26602 4468 26608 4480
rect 26563 4440 26608 4468
rect 26602 4428 26608 4440
rect 26660 4428 26666 4480
rect 27246 4468 27252 4480
rect 27207 4440 27252 4468
rect 27246 4428 27252 4440
rect 27304 4428 27310 4480
rect 27706 4468 27712 4480
rect 27667 4440 27712 4468
rect 27706 4428 27712 4440
rect 27764 4428 27770 4480
rect 33502 4428 33508 4480
rect 33560 4468 33566 4480
rect 33781 4471 33839 4477
rect 33781 4468 33793 4471
rect 33560 4440 33793 4468
rect 33560 4428 33566 4440
rect 33781 4437 33793 4440
rect 33827 4437 33839 4471
rect 34790 4468 34796 4480
rect 34751 4440 34796 4468
rect 33781 4431 33839 4437
rect 34790 4428 34796 4440
rect 34848 4428 34854 4480
rect 35342 4468 35348 4480
rect 35303 4440 35348 4468
rect 35342 4428 35348 4440
rect 35400 4428 35406 4480
rect 36556 4477 36584 4508
rect 42153 4505 42165 4539
rect 42199 4536 42211 4539
rect 42978 4536 42984 4548
rect 42199 4508 42984 4536
rect 42199 4505 42211 4508
rect 42153 4499 42211 4505
rect 42978 4496 42984 4508
rect 43036 4496 43042 4548
rect 44085 4539 44143 4545
rect 44085 4505 44097 4539
rect 44131 4536 44143 4539
rect 44174 4536 44180 4548
rect 44131 4508 44180 4536
rect 44131 4505 44143 4508
rect 44085 4499 44143 4505
rect 44174 4496 44180 4508
rect 44232 4536 44238 4548
rect 44818 4536 44824 4548
rect 44232 4508 44824 4536
rect 44232 4496 44238 4508
rect 44818 4496 44824 4508
rect 44876 4496 44882 4548
rect 36541 4471 36599 4477
rect 36541 4437 36553 4471
rect 36587 4468 36599 4471
rect 36630 4468 36636 4480
rect 36587 4440 36636 4468
rect 36587 4437 36599 4440
rect 36541 4431 36599 4437
rect 36630 4428 36636 4440
rect 36688 4428 36694 4480
rect 37274 4468 37280 4480
rect 37235 4440 37280 4468
rect 37274 4428 37280 4440
rect 37332 4428 37338 4480
rect 38654 4468 38660 4480
rect 38615 4440 38660 4468
rect 38654 4428 38660 4440
rect 38712 4428 38718 4480
rect 39850 4468 39856 4480
rect 39811 4440 39856 4468
rect 39850 4428 39856 4440
rect 39908 4428 39914 4480
rect 41417 4471 41475 4477
rect 41417 4437 41429 4471
rect 41463 4468 41475 4471
rect 41506 4468 41512 4480
rect 41463 4440 41512 4468
rect 41463 4437 41475 4440
rect 41417 4431 41475 4437
rect 41506 4428 41512 4440
rect 41564 4428 41570 4480
rect 42705 4471 42763 4477
rect 42705 4437 42717 4471
rect 42751 4468 42763 4471
rect 43162 4468 43168 4480
rect 42751 4440 43168 4468
rect 42751 4437 42763 4440
rect 42705 4431 42763 4437
rect 43162 4428 43168 4440
rect 43220 4428 43226 4480
rect 43346 4468 43352 4480
rect 43307 4440 43352 4468
rect 43346 4428 43352 4440
rect 43404 4428 43410 4480
rect 1104 4378 44896 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 44896 4378
rect 1104 4304 44896 4326
rect 5810 4264 5816 4276
rect 5771 4236 5816 4264
rect 5810 4224 5816 4236
rect 5868 4224 5874 4276
rect 9490 4264 9496 4276
rect 9451 4236 9496 4264
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 21450 4264 21456 4276
rect 9732 4236 21456 4264
rect 9732 4224 9738 4236
rect 21450 4224 21456 4236
rect 21508 4224 21514 4276
rect 43530 4224 43536 4276
rect 43588 4264 43594 4276
rect 43588 4236 44128 4264
rect 43588 4224 43594 4236
rect 1394 4156 1400 4208
rect 1452 4196 1458 4208
rect 3973 4199 4031 4205
rect 3973 4196 3985 4199
rect 1452 4168 3985 4196
rect 1452 4156 1458 4168
rect 3973 4165 3985 4168
rect 4019 4165 4031 4199
rect 3973 4159 4031 4165
rect 10045 4199 10103 4205
rect 10045 4165 10057 4199
rect 10091 4196 10103 4199
rect 10410 4196 10416 4208
rect 10091 4168 10416 4196
rect 10091 4165 10103 4168
rect 10045 4159 10103 4165
rect 10410 4156 10416 4168
rect 10468 4156 10474 4208
rect 10686 4196 10692 4208
rect 10647 4168 10692 4196
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 11422 4156 11428 4208
rect 11480 4156 11486 4208
rect 11606 4196 11612 4208
rect 11567 4168 11612 4196
rect 11606 4156 11612 4168
rect 11664 4196 11670 4208
rect 12621 4199 12679 4205
rect 12621 4196 12633 4199
rect 11664 4168 12633 4196
rect 11664 4156 11670 4168
rect 12621 4165 12633 4168
rect 12667 4196 12679 4199
rect 13354 4196 13360 4208
rect 12667 4168 13360 4196
rect 12667 4165 12679 4168
rect 12621 4159 12679 4165
rect 13354 4156 13360 4168
rect 13412 4156 13418 4208
rect 14182 4156 14188 4208
rect 14240 4196 14246 4208
rect 14369 4199 14427 4205
rect 14369 4196 14381 4199
rect 14240 4168 14381 4196
rect 14240 4156 14246 4168
rect 14369 4165 14381 4168
rect 14415 4165 14427 4199
rect 14369 4159 14427 4165
rect 19444 4168 19656 4196
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 7374 4128 7380 4140
rect 3936 4100 7380 4128
rect 3936 4088 3942 4100
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7742 4128 7748 4140
rect 7703 4100 7748 4128
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 8018 4088 8024 4140
rect 8076 4128 8082 4140
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8076 4100 8401 4128
rect 8076 4088 8082 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 11440 4128 11468 4156
rect 8389 4091 8447 4097
rect 10796 4100 11468 4128
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4060 7343 4063
rect 7926 4060 7932 4072
rect 7331 4032 7932 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 1302 3952 1308 4004
rect 1360 3992 1366 4004
rect 2041 3995 2099 4001
rect 2041 3992 2053 3995
rect 1360 3964 2053 3992
rect 1360 3952 1366 3964
rect 2041 3961 2053 3964
rect 2087 3961 2099 3995
rect 2041 3955 2099 3961
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3992 4767 3995
rect 8478 3992 8484 4004
rect 4755 3964 8484 3992
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 8478 3952 8484 3964
rect 8536 3952 8542 4004
rect 8573 3995 8631 4001
rect 8573 3961 8585 3995
rect 8619 3992 8631 3995
rect 9214 3992 9220 4004
rect 8619 3964 9220 3992
rect 8619 3961 8631 3964
rect 8573 3955 8631 3961
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 106 3884 112 3936
rect 164 3924 170 3936
rect 1397 3927 1455 3933
rect 1397 3924 1409 3927
rect 164 3896 1409 3924
rect 164 3884 170 3896
rect 1397 3893 1409 3896
rect 1443 3893 1455 3927
rect 1397 3887 1455 3893
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2685 3927 2743 3933
rect 2685 3924 2697 3927
rect 2004 3896 2697 3924
rect 2004 3884 2010 3896
rect 2685 3893 2697 3896
rect 2731 3893 2743 3927
rect 2685 3887 2743 3893
rect 3234 3884 3240 3936
rect 3292 3924 3298 3936
rect 3329 3927 3387 3933
rect 3329 3924 3341 3927
rect 3292 3896 3341 3924
rect 3292 3884 3298 3896
rect 3329 3893 3341 3896
rect 3375 3893 3387 3927
rect 3329 3887 3387 3893
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 5169 3927 5227 3933
rect 5169 3924 5181 3927
rect 5132 3896 5181 3924
rect 5132 3884 5138 3896
rect 5169 3893 5181 3896
rect 5215 3893 5227 3927
rect 5169 3887 5227 3893
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 6730 3924 6736 3936
rect 5776 3896 6736 3924
rect 5776 3884 5782 3896
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7929 3927 7987 3933
rect 7929 3893 7941 3927
rect 7975 3924 7987 3927
rect 10796 3924 10824 4100
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 13173 4131 13231 4137
rect 13173 4128 13185 4131
rect 12860 4100 13185 4128
rect 12860 4088 12866 4100
rect 13173 4097 13185 4100
rect 13219 4097 13231 4131
rect 13173 4091 13231 4097
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4128 13875 4131
rect 14274 4128 14280 4140
rect 13863 4100 14280 4128
rect 13863 4097 13875 4100
rect 13817 4091 13875 4097
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 15838 4128 15844 4140
rect 14384 4100 15844 4128
rect 11422 4020 11428 4072
rect 11480 4060 11486 4072
rect 14384 4060 14412 4100
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 16574 4088 16580 4140
rect 16632 4128 16638 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16632 4100 16681 4128
rect 16632 4088 16638 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 17402 4128 17408 4140
rect 17363 4100 17408 4128
rect 16669 4091 16727 4097
rect 15378 4060 15384 4072
rect 11480 4032 14136 4060
rect 11480 4020 11486 4032
rect 12158 3992 12164 4004
rect 12071 3964 12164 3992
rect 12158 3952 12164 3964
rect 12216 3992 12222 4004
rect 13538 3992 13544 4004
rect 12216 3964 13544 3992
rect 12216 3952 12222 3964
rect 13538 3952 13544 3964
rect 13596 3952 13602 4004
rect 14108 3992 14136 4032
rect 14292 4032 14412 4060
rect 15339 4032 15384 4060
rect 14292 3992 14320 4032
rect 15378 4020 15384 4032
rect 15436 4020 15442 4072
rect 16684 4060 16712 4091
rect 17402 4088 17408 4100
rect 17460 4128 17466 4140
rect 18230 4128 18236 4140
rect 17460 4100 18236 4128
rect 17460 4088 17466 4100
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 18417 4131 18475 4137
rect 18417 4128 18429 4131
rect 18380 4100 18429 4128
rect 18380 4088 18386 4100
rect 18417 4097 18429 4100
rect 18463 4128 18475 4131
rect 18506 4128 18512 4140
rect 18463 4100 18512 4128
rect 18463 4097 18475 4100
rect 18417 4091 18475 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 19444 4128 19472 4168
rect 18616 4100 19472 4128
rect 19521 4131 19579 4137
rect 17586 4060 17592 4072
rect 16684 4032 17592 4060
rect 17586 4020 17592 4032
rect 17644 4020 17650 4072
rect 14108 3964 14320 3992
rect 14366 3952 14372 4004
rect 14424 3992 14430 4004
rect 18616 3992 18644 4100
rect 19521 4097 19533 4131
rect 19567 4097 19579 4131
rect 19628 4128 19656 4168
rect 22738 4156 22744 4208
rect 22796 4196 22802 4208
rect 25130 4196 25136 4208
rect 22796 4168 25136 4196
rect 22796 4156 22802 4168
rect 25130 4156 25136 4168
rect 25188 4156 25194 4208
rect 43349 4199 43407 4205
rect 43349 4165 43361 4199
rect 43395 4196 43407 4199
rect 43806 4196 43812 4208
rect 43395 4168 43812 4196
rect 43395 4165 43407 4168
rect 43349 4159 43407 4165
rect 43806 4156 43812 4168
rect 43864 4156 43870 4208
rect 44100 4205 44128 4236
rect 44085 4199 44143 4205
rect 44085 4165 44097 4199
rect 44131 4196 44143 4199
rect 45462 4196 45468 4208
rect 44131 4168 45468 4196
rect 44131 4165 44143 4168
rect 44085 4159 44143 4165
rect 45462 4156 45468 4168
rect 45520 4156 45526 4208
rect 19981 4131 20039 4137
rect 19981 4128 19993 4131
rect 19628 4100 19993 4128
rect 19521 4091 19579 4097
rect 19981 4097 19993 4100
rect 20027 4097 20039 4131
rect 19981 4091 20039 4097
rect 19150 4020 19156 4072
rect 19208 4060 19214 4072
rect 19536 4060 19564 4091
rect 21634 4088 21640 4140
rect 21692 4128 21698 4140
rect 21692 4100 21956 4128
rect 21692 4088 21698 4100
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 19208 4032 21833 4060
rect 19208 4020 19214 4032
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 21928 4060 21956 4100
rect 22370 4088 22376 4140
rect 22428 4128 22434 4140
rect 26237 4131 26295 4137
rect 26237 4128 26249 4131
rect 22428 4100 26249 4128
rect 22428 4088 22434 4100
rect 26237 4097 26249 4100
rect 26283 4097 26295 4131
rect 26237 4091 26295 4097
rect 27525 4131 27583 4137
rect 27525 4097 27537 4131
rect 27571 4128 27583 4131
rect 27982 4128 27988 4140
rect 27571 4100 27988 4128
rect 27571 4097 27583 4100
rect 27525 4091 27583 4097
rect 27982 4088 27988 4100
rect 28040 4088 28046 4140
rect 41690 4088 41696 4140
rect 41748 4128 41754 4140
rect 42429 4131 42487 4137
rect 42429 4128 42441 4131
rect 41748 4100 42441 4128
rect 41748 4088 41754 4100
rect 42429 4097 42441 4100
rect 42475 4097 42487 4131
rect 42429 4091 42487 4097
rect 43165 4131 43223 4137
rect 43165 4097 43177 4131
rect 43211 4128 43223 4131
rect 43254 4128 43260 4140
rect 43211 4100 43260 4128
rect 43211 4097 43223 4100
rect 43165 4091 43223 4097
rect 43254 4088 43260 4100
rect 43312 4088 43318 4140
rect 43901 4131 43959 4137
rect 43901 4097 43913 4131
rect 43947 4128 43959 4131
rect 43990 4128 43996 4140
rect 43947 4100 43996 4128
rect 43947 4097 43959 4100
rect 43901 4091 43959 4097
rect 43990 4088 43996 4100
rect 44048 4088 44054 4140
rect 21928 4032 31754 4060
rect 21821 4023 21879 4029
rect 19334 3992 19340 4004
rect 14424 3964 18644 3992
rect 19295 3964 19340 3992
rect 14424 3952 14430 3964
rect 19334 3952 19340 3964
rect 19392 3952 19398 4004
rect 20254 3952 20260 4004
rect 20312 3992 20318 4004
rect 22373 3995 22431 4001
rect 22373 3992 22385 3995
rect 20312 3964 22385 3992
rect 20312 3952 20318 3964
rect 22373 3961 22385 3964
rect 22419 3961 22431 3995
rect 22373 3955 22431 3961
rect 23569 3995 23627 4001
rect 23569 3961 23581 3995
rect 23615 3992 23627 3995
rect 24118 3992 24124 4004
rect 23615 3964 24124 3992
rect 23615 3961 23627 3964
rect 23569 3955 23627 3961
rect 24118 3952 24124 3964
rect 24176 3952 24182 4004
rect 31726 3992 31754 4032
rect 33042 4020 33048 4072
rect 33100 4060 33106 4072
rect 33597 4063 33655 4069
rect 33597 4060 33609 4063
rect 33100 4032 33609 4060
rect 33100 4020 33106 4032
rect 33597 4029 33609 4032
rect 33643 4029 33655 4063
rect 33597 4023 33655 4029
rect 36906 4020 36912 4072
rect 36964 4060 36970 4072
rect 37829 4063 37887 4069
rect 37829 4060 37841 4063
rect 36964 4032 37841 4060
rect 36964 4020 36970 4032
rect 37829 4029 37841 4032
rect 37875 4029 37887 4063
rect 37829 4023 37887 4029
rect 37366 3992 37372 4004
rect 31726 3964 37372 3992
rect 37366 3952 37372 3964
rect 37424 3952 37430 4004
rect 41877 3995 41935 4001
rect 41877 3961 41889 3995
rect 41923 3992 41935 3995
rect 44450 3992 44456 4004
rect 41923 3964 44456 3992
rect 41923 3961 41935 3964
rect 41877 3955 41935 3961
rect 44450 3952 44456 3964
rect 44508 3952 44514 4004
rect 7975 3896 10824 3924
rect 7975 3893 7987 3896
rect 7929 3887 7987 3893
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 14090 3924 14096 3936
rect 13872 3896 14096 3924
rect 13872 3884 13878 3896
rect 14090 3884 14096 3896
rect 14148 3924 14154 3936
rect 14829 3927 14887 3933
rect 14829 3924 14841 3927
rect 14148 3896 14841 3924
rect 14148 3884 14154 3896
rect 14829 3893 14841 3896
rect 14875 3893 14887 3927
rect 14829 3887 14887 3893
rect 15286 3884 15292 3936
rect 15344 3924 15350 3936
rect 15933 3927 15991 3933
rect 15933 3924 15945 3927
rect 15344 3896 15945 3924
rect 15344 3884 15350 3896
rect 15933 3893 15945 3896
rect 15979 3893 15991 3927
rect 15933 3887 15991 3893
rect 18601 3927 18659 3933
rect 18601 3893 18613 3927
rect 18647 3924 18659 3927
rect 19242 3924 19248 3936
rect 18647 3896 19248 3924
rect 18647 3893 18659 3896
rect 18601 3887 18659 3893
rect 19242 3884 19248 3896
rect 19300 3884 19306 3936
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 20533 3927 20591 3933
rect 20533 3924 20545 3927
rect 20496 3896 20545 3924
rect 20496 3884 20502 3896
rect 20533 3893 20545 3896
rect 20579 3893 20591 3927
rect 21082 3924 21088 3936
rect 21043 3896 21088 3924
rect 20533 3887 20591 3893
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 22922 3924 22928 3936
rect 22883 3896 22928 3924
rect 22922 3884 22928 3896
rect 22980 3884 22986 3936
rect 23934 3884 23940 3936
rect 23992 3924 23998 3936
rect 24029 3927 24087 3933
rect 24029 3924 24041 3927
rect 23992 3896 24041 3924
rect 23992 3884 23998 3896
rect 24029 3893 24041 3896
rect 24075 3893 24087 3927
rect 24578 3924 24584 3936
rect 24539 3896 24584 3924
rect 24029 3887 24087 3893
rect 24578 3884 24584 3896
rect 24636 3884 24642 3936
rect 25130 3924 25136 3936
rect 25091 3896 25136 3924
rect 25130 3884 25136 3896
rect 25188 3884 25194 3936
rect 25314 3884 25320 3936
rect 25372 3924 25378 3936
rect 25685 3927 25743 3933
rect 25685 3924 25697 3927
rect 25372 3896 25697 3924
rect 25372 3884 25378 3896
rect 25685 3893 25697 3896
rect 25731 3893 25743 3927
rect 25685 3887 25743 3893
rect 27154 3884 27160 3936
rect 27212 3924 27218 3936
rect 27341 3927 27399 3933
rect 27341 3924 27353 3927
rect 27212 3896 27353 3924
rect 27212 3884 27218 3896
rect 27341 3893 27353 3896
rect 27387 3893 27399 3927
rect 27982 3924 27988 3936
rect 27943 3896 27988 3924
rect 27341 3887 27399 3893
rect 27982 3884 27988 3896
rect 28040 3884 28046 3936
rect 28718 3924 28724 3936
rect 28679 3896 28724 3924
rect 28718 3884 28724 3896
rect 28776 3884 28782 3936
rect 29362 3924 29368 3936
rect 29323 3896 29368 3924
rect 29362 3884 29368 3896
rect 29420 3884 29426 3936
rect 30009 3927 30067 3933
rect 30009 3893 30021 3927
rect 30055 3924 30067 3927
rect 30282 3924 30288 3936
rect 30055 3896 30288 3924
rect 30055 3893 30067 3896
rect 30009 3887 30067 3893
rect 30282 3884 30288 3896
rect 30340 3884 30346 3936
rect 30742 3924 30748 3936
rect 30703 3896 30748 3924
rect 30742 3884 30748 3896
rect 30800 3884 30806 3936
rect 31202 3924 31208 3936
rect 31163 3896 31208 3924
rect 31202 3884 31208 3896
rect 31260 3884 31266 3936
rect 31662 3884 31668 3936
rect 31720 3924 31726 3936
rect 32309 3927 32367 3933
rect 32309 3924 32321 3927
rect 31720 3896 32321 3924
rect 31720 3884 31726 3896
rect 32309 3893 32321 3896
rect 32355 3893 32367 3927
rect 32309 3887 32367 3893
rect 33137 3927 33195 3933
rect 33137 3893 33149 3927
rect 33183 3924 33195 3927
rect 33318 3924 33324 3936
rect 33183 3896 33324 3924
rect 33183 3893 33195 3896
rect 33137 3887 33195 3893
rect 33318 3884 33324 3896
rect 33376 3884 33382 3936
rect 34606 3924 34612 3936
rect 34567 3896 34612 3924
rect 34606 3884 34612 3896
rect 34664 3884 34670 3936
rect 35345 3927 35403 3933
rect 35345 3893 35357 3927
rect 35391 3924 35403 3927
rect 35434 3924 35440 3936
rect 35391 3896 35440 3924
rect 35391 3893 35403 3896
rect 35345 3887 35403 3893
rect 35434 3884 35440 3896
rect 35492 3884 35498 3936
rect 36078 3924 36084 3936
rect 36039 3896 36084 3924
rect 36078 3884 36084 3896
rect 36136 3884 36142 3936
rect 36262 3884 36268 3936
rect 36320 3924 36326 3936
rect 36541 3927 36599 3933
rect 36541 3924 36553 3927
rect 36320 3896 36553 3924
rect 36320 3884 36326 3896
rect 36541 3893 36553 3896
rect 36587 3893 36599 3927
rect 36541 3887 36599 3893
rect 37182 3884 37188 3936
rect 37240 3924 37246 3936
rect 37277 3927 37335 3933
rect 37277 3924 37289 3927
rect 37240 3896 37289 3924
rect 37240 3884 37246 3896
rect 37277 3893 37289 3896
rect 37323 3893 37335 3927
rect 38838 3924 38844 3936
rect 38799 3896 38844 3924
rect 37277 3887 37335 3893
rect 38838 3884 38844 3896
rect 38896 3884 38902 3936
rect 39758 3924 39764 3936
rect 39719 3896 39764 3924
rect 39758 3884 39764 3896
rect 39816 3884 39822 3936
rect 39942 3884 39948 3936
rect 40000 3924 40006 3936
rect 40221 3927 40279 3933
rect 40221 3924 40233 3927
rect 40000 3896 40233 3924
rect 40000 3884 40006 3896
rect 40221 3893 40233 3896
rect 40267 3893 40279 3927
rect 40221 3887 40279 3893
rect 40402 3884 40408 3936
rect 40460 3924 40466 3936
rect 40773 3927 40831 3933
rect 40773 3924 40785 3927
rect 40460 3896 40785 3924
rect 40460 3884 40466 3896
rect 40773 3893 40785 3896
rect 40819 3893 40831 3927
rect 40773 3887 40831 3893
rect 42613 3927 42671 3933
rect 42613 3893 42625 3927
rect 42659 3924 42671 3927
rect 44174 3924 44180 3936
rect 42659 3896 44180 3924
rect 42659 3893 42671 3896
rect 42613 3887 42671 3893
rect 44174 3884 44180 3896
rect 44232 3884 44238 3936
rect 1104 3834 44896 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 44896 3834
rect 1104 3760 44896 3782
rect 6638 3720 6644 3732
rect 6599 3692 6644 3720
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 9490 3720 9496 3732
rect 9451 3692 9496 3720
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 9950 3720 9956 3732
rect 9911 3692 9956 3720
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10781 3723 10839 3729
rect 10781 3689 10793 3723
rect 10827 3720 10839 3723
rect 10870 3720 10876 3732
rect 10827 3692 10876 3720
rect 10827 3689 10839 3692
rect 10781 3683 10839 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 11422 3720 11428 3732
rect 11383 3692 11428 3720
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 11514 3680 11520 3732
rect 11572 3720 11578 3732
rect 11885 3723 11943 3729
rect 11885 3720 11897 3723
rect 11572 3692 11897 3720
rect 11572 3680 11578 3692
rect 11885 3689 11897 3692
rect 11931 3689 11943 3723
rect 13354 3720 13360 3732
rect 13315 3692 13360 3720
rect 11885 3683 11943 3689
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 13964 3692 14105 3720
rect 13964 3680 13970 3692
rect 14093 3689 14105 3692
rect 14139 3689 14151 3723
rect 14093 3683 14151 3689
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 16577 3723 16635 3729
rect 16577 3720 16589 3723
rect 14700 3692 16589 3720
rect 14700 3680 14706 3692
rect 16577 3689 16589 3692
rect 16623 3689 16635 3723
rect 16577 3683 16635 3689
rect 18325 3723 18383 3729
rect 18325 3689 18337 3723
rect 18371 3720 18383 3723
rect 18874 3720 18880 3732
rect 18371 3692 18880 3720
rect 18371 3689 18383 3692
rect 18325 3683 18383 3689
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 19429 3723 19487 3729
rect 19429 3689 19441 3723
rect 19475 3720 19487 3723
rect 20162 3720 20168 3732
rect 19475 3692 20168 3720
rect 19475 3689 19487 3692
rect 19429 3683 19487 3689
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20533 3723 20591 3729
rect 20533 3689 20545 3723
rect 20579 3720 20591 3723
rect 20990 3720 20996 3732
rect 20579 3692 20996 3720
rect 20579 3689 20591 3692
rect 20533 3683 20591 3689
rect 20990 3680 20996 3692
rect 21048 3680 21054 3732
rect 21269 3723 21327 3729
rect 21269 3689 21281 3723
rect 21315 3720 21327 3723
rect 21358 3720 21364 3732
rect 21315 3692 21364 3720
rect 21315 3689 21327 3692
rect 21269 3683 21327 3689
rect 21358 3680 21364 3692
rect 21416 3680 21422 3732
rect 27522 3720 27528 3732
rect 22066 3692 27528 3720
rect 658 3612 664 3664
rect 716 3652 722 3664
rect 2685 3655 2743 3661
rect 2685 3652 2697 3655
rect 716 3624 2697 3652
rect 716 3612 722 3624
rect 2685 3621 2697 3624
rect 2731 3621 2743 3655
rect 3970 3652 3976 3664
rect 3931 3624 3976 3652
rect 2685 3615 2743 3621
rect 3970 3612 3976 3624
rect 4028 3612 4034 3664
rect 5997 3655 6055 3661
rect 5997 3621 6009 3655
rect 6043 3652 6055 3655
rect 10042 3652 10048 3664
rect 6043 3624 10048 3652
rect 6043 3621 6055 3624
rect 5997 3615 6055 3621
rect 10042 3612 10048 3624
rect 10100 3612 10106 3664
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 12713 3655 12771 3661
rect 12713 3652 12725 3655
rect 11756 3624 12725 3652
rect 11756 3612 11762 3624
rect 12713 3621 12725 3624
rect 12759 3621 12771 3655
rect 14734 3652 14740 3664
rect 14695 3624 14740 3652
rect 12713 3615 12771 3621
rect 14734 3612 14740 3624
rect 14792 3612 14798 3664
rect 14826 3612 14832 3664
rect 14884 3652 14890 3664
rect 15565 3655 15623 3661
rect 15565 3652 15577 3655
rect 14884 3624 15577 3652
rect 14884 3612 14890 3624
rect 15565 3621 15577 3624
rect 15611 3621 15623 3655
rect 20438 3652 20444 3664
rect 15565 3615 15623 3621
rect 15764 3624 20444 3652
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 7466 3584 7472 3596
rect 1995 3556 7472 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 7650 3584 7656 3596
rect 7611 3556 7656 3584
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 15010 3584 15016 3596
rect 8352 3556 15016 3584
rect 8352 3544 8358 3556
rect 15010 3544 15016 3556
rect 15068 3544 15074 3596
rect 1026 3476 1032 3528
rect 1084 3516 1090 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 1084 3488 2237 3516
rect 1084 3476 1090 3488
rect 2225 3485 2237 3488
rect 2271 3516 2283 3519
rect 2271 3488 2774 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2746 3448 2774 3488
rect 2958 3476 2964 3528
rect 3016 3516 3022 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3016 3488 3801 3516
rect 3016 3476 3022 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 4212 3488 4445 3516
rect 4212 3476 4218 3488
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5776 3488 5825 3516
rect 5776 3476 5782 3488
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 6144 3488 6469 3516
rect 6144 3476 6150 3488
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 7926 3516 7932 3528
rect 7887 3488 7932 3516
rect 6457 3479 6515 3485
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 9306 3516 9312 3528
rect 9267 3488 9312 3516
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 10594 3516 10600 3528
rect 10555 3488 10600 3516
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 11238 3516 11244 3528
rect 11199 3488 11244 3516
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 12069 3519 12127 3525
rect 12069 3485 12081 3519
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3485 12955 3519
rect 12897 3479 12955 3485
rect 5166 3448 5172 3460
rect 2746 3420 5172 3448
rect 5166 3408 5172 3420
rect 5224 3408 5230 3460
rect 5353 3451 5411 3457
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 11698 3448 11704 3460
rect 5399 3420 11704 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 11698 3408 11704 3420
rect 11756 3448 11762 3460
rect 12084 3448 12112 3479
rect 11756 3420 12112 3448
rect 11756 3408 11762 3420
rect 12618 3408 12624 3460
rect 12676 3448 12682 3460
rect 12912 3448 12940 3479
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13688 3488 14289 3516
rect 13688 3476 13694 3488
rect 14277 3485 14289 3488
rect 14323 3516 14335 3519
rect 14366 3516 14372 3528
rect 14323 3488 14372 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 15654 3476 15660 3528
rect 15712 3516 15718 3528
rect 15764 3525 15792 3624
rect 20438 3612 20444 3624
rect 20496 3612 20502 3664
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 22066 3652 22094 3692
rect 27522 3680 27528 3692
rect 27580 3680 27586 3732
rect 37458 3720 37464 3732
rect 27632 3692 35894 3720
rect 37419 3692 37464 3720
rect 20772 3624 22094 3652
rect 20772 3612 20778 3624
rect 22646 3612 22652 3664
rect 22704 3652 22710 3664
rect 25041 3655 25099 3661
rect 25041 3652 25053 3655
rect 22704 3624 25053 3652
rect 22704 3612 22710 3624
rect 25041 3621 25053 3624
rect 25087 3621 25099 3655
rect 25041 3615 25099 3621
rect 27249 3655 27307 3661
rect 27249 3621 27261 3655
rect 27295 3652 27307 3655
rect 27338 3652 27344 3664
rect 27295 3624 27344 3652
rect 27295 3621 27307 3624
rect 27249 3615 27307 3621
rect 27338 3612 27344 3624
rect 27396 3612 27402 3664
rect 27430 3612 27436 3664
rect 27488 3652 27494 3664
rect 27632 3652 27660 3692
rect 27488 3624 27660 3652
rect 28169 3655 28227 3661
rect 27488 3612 27494 3624
rect 28169 3621 28181 3655
rect 28215 3652 28227 3655
rect 30098 3652 30104 3664
rect 28215 3624 30104 3652
rect 28215 3621 28227 3624
rect 28169 3615 28227 3621
rect 30098 3612 30104 3624
rect 30156 3612 30162 3664
rect 19978 3584 19984 3596
rect 16776 3556 19984 3584
rect 15749 3519 15807 3525
rect 15749 3516 15761 3519
rect 15712 3488 15761 3516
rect 15712 3476 15718 3488
rect 15749 3485 15761 3488
rect 15795 3485 15807 3519
rect 15749 3479 15807 3485
rect 16482 3476 16488 3528
rect 16540 3516 16546 3528
rect 16776 3525 16804 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 20070 3544 20076 3596
rect 20128 3584 20134 3596
rect 20128 3556 23336 3584
rect 20128 3544 20134 3556
rect 16761 3519 16819 3525
rect 16761 3516 16773 3519
rect 16540 3488 16773 3516
rect 16540 3476 16546 3488
rect 16761 3485 16773 3488
rect 16807 3485 16819 3519
rect 18138 3516 18144 3528
rect 18099 3488 18144 3516
rect 16761 3479 16819 3485
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 18966 3476 18972 3528
rect 19024 3516 19030 3528
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 19024 3488 19257 3516
rect 19024 3476 19030 3488
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 20346 3516 20352 3528
rect 20307 3488 20352 3516
rect 19245 3479 19303 3485
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 21266 3476 21272 3528
rect 21324 3516 21330 3528
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 21324 3488 21465 3516
rect 21324 3476 21330 3488
rect 21453 3485 21465 3488
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 22094 3476 22100 3528
rect 22152 3516 22158 3528
rect 22373 3519 22431 3525
rect 22373 3516 22385 3519
rect 22152 3488 22385 3516
rect 22152 3476 22158 3488
rect 22373 3485 22385 3488
rect 22419 3516 22431 3519
rect 22738 3516 22744 3528
rect 22419 3488 22744 3516
rect 22419 3485 22431 3488
rect 22373 3479 22431 3485
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 17954 3448 17960 3460
rect 12676 3420 17960 3448
rect 12676 3408 12682 3420
rect 17954 3408 17960 3420
rect 18012 3408 18018 3460
rect 19334 3448 19340 3460
rect 18064 3420 19340 3448
rect 4614 3380 4620 3392
rect 4575 3352 4620 3380
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 16574 3340 16580 3392
rect 16632 3380 16638 3392
rect 17221 3383 17279 3389
rect 17221 3380 17233 3383
rect 16632 3352 17233 3380
rect 16632 3340 16638 3352
rect 17221 3349 17233 3352
rect 17267 3349 17279 3383
rect 17221 3343 17279 3349
rect 17862 3340 17868 3392
rect 17920 3380 17926 3392
rect 18064 3380 18092 3420
rect 19334 3408 19340 3420
rect 19392 3408 19398 3460
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 19484 3420 23244 3448
rect 19484 3408 19490 3420
rect 17920 3352 18092 3380
rect 17920 3340 17926 3352
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 23216 3389 23244 3420
rect 22189 3383 22247 3389
rect 22189 3380 22201 3383
rect 18656 3352 22201 3380
rect 18656 3340 18662 3352
rect 22189 3349 22201 3352
rect 22235 3349 22247 3383
rect 22189 3343 22247 3349
rect 23201 3383 23259 3389
rect 23201 3349 23213 3383
rect 23247 3349 23259 3383
rect 23308 3380 23336 3556
rect 23566 3544 23572 3596
rect 23624 3584 23630 3596
rect 25682 3584 25688 3596
rect 23624 3556 25688 3584
rect 23624 3544 23630 3556
rect 25682 3544 25688 3556
rect 25740 3544 25746 3596
rect 28350 3544 28356 3596
rect 28408 3584 28414 3596
rect 35866 3584 35894 3692
rect 37458 3680 37464 3692
rect 37516 3680 37522 3732
rect 43070 3612 43076 3664
rect 43128 3652 43134 3664
rect 43165 3655 43223 3661
rect 43165 3652 43177 3655
rect 43128 3624 43177 3652
rect 43128 3612 43134 3624
rect 43165 3621 43177 3624
rect 43211 3621 43223 3655
rect 43898 3652 43904 3664
rect 43859 3624 43904 3652
rect 43165 3615 43223 3621
rect 43898 3612 43904 3624
rect 43956 3612 43962 3664
rect 43990 3584 43996 3596
rect 28408 3556 30328 3584
rect 35866 3556 43996 3584
rect 28408 3544 28414 3556
rect 23382 3476 23388 3528
rect 23440 3516 23446 3528
rect 23440 3488 23485 3516
rect 23440 3476 23446 3488
rect 24026 3476 24032 3528
rect 24084 3516 24090 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 24084 3488 24593 3516
rect 24084 3476 24090 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 24946 3476 24952 3528
rect 25004 3516 25010 3528
rect 25222 3516 25228 3528
rect 25004 3488 25228 3516
rect 25004 3476 25010 3488
rect 25222 3476 25228 3488
rect 25280 3476 25286 3528
rect 26513 3519 26571 3525
rect 26513 3485 26525 3519
rect 26559 3516 26571 3519
rect 27614 3516 27620 3528
rect 26559 3488 27620 3516
rect 26559 3485 26571 3488
rect 26513 3479 26571 3485
rect 27614 3476 27620 3488
rect 27672 3476 27678 3528
rect 27982 3516 27988 3528
rect 27943 3488 27988 3516
rect 27982 3476 27988 3488
rect 28040 3476 28046 3528
rect 28810 3476 28816 3528
rect 28868 3516 28874 3528
rect 28905 3519 28963 3525
rect 28905 3516 28917 3519
rect 28868 3488 28917 3516
rect 28868 3476 28874 3488
rect 28905 3485 28917 3488
rect 28951 3485 28963 3519
rect 29546 3516 29552 3528
rect 29507 3488 29552 3516
rect 28905 3479 28963 3485
rect 29546 3476 29552 3488
rect 29604 3476 29610 3528
rect 30300 3525 30328 3556
rect 43990 3544 43996 3556
rect 44048 3544 44054 3596
rect 30285 3519 30343 3525
rect 30285 3485 30297 3519
rect 30331 3485 30343 3519
rect 31018 3516 31024 3528
rect 30979 3488 31024 3516
rect 30285 3479 30343 3485
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 31938 3516 31944 3528
rect 31899 3488 31944 3516
rect 31938 3476 31944 3488
rect 31996 3476 32002 3528
rect 32950 3516 32956 3528
rect 32911 3488 32956 3516
rect 32950 3476 32956 3488
rect 33008 3476 33014 3528
rect 33870 3516 33876 3528
rect 33831 3488 33876 3516
rect 33870 3476 33876 3488
rect 33928 3476 33934 3528
rect 34514 3476 34520 3528
rect 34572 3516 34578 3528
rect 34793 3519 34851 3525
rect 34793 3516 34805 3519
rect 34572 3488 34805 3516
rect 34572 3476 34578 3488
rect 34793 3485 34805 3488
rect 34839 3485 34851 3519
rect 34793 3479 34851 3485
rect 35713 3519 35771 3525
rect 35713 3485 35725 3519
rect 35759 3516 35771 3519
rect 35894 3516 35900 3528
rect 35759 3488 35900 3516
rect 35759 3485 35771 3488
rect 35713 3479 35771 3485
rect 35894 3476 35900 3488
rect 35952 3476 35958 3528
rect 36630 3516 36636 3528
rect 36591 3488 36636 3516
rect 36630 3476 36636 3488
rect 36688 3476 36694 3528
rect 37918 3476 37924 3528
rect 37976 3516 37982 3528
rect 38105 3519 38163 3525
rect 38105 3516 38117 3519
rect 37976 3488 38117 3516
rect 37976 3476 37982 3488
rect 38105 3485 38117 3488
rect 38151 3485 38163 3519
rect 39114 3516 39120 3528
rect 39075 3488 39120 3516
rect 38105 3479 38163 3485
rect 39114 3476 39120 3488
rect 39172 3476 39178 3528
rect 39850 3516 39856 3528
rect 39811 3488 39856 3516
rect 39850 3476 39856 3488
rect 39908 3476 39914 3528
rect 41414 3476 41420 3528
rect 41472 3516 41478 3528
rect 41601 3519 41659 3525
rect 41601 3516 41613 3519
rect 41472 3488 41613 3516
rect 41472 3476 41478 3488
rect 41601 3485 41613 3488
rect 41647 3485 41659 3519
rect 42334 3516 42340 3528
rect 42295 3488 42340 3516
rect 41601 3479 41659 3485
rect 42334 3476 42340 3488
rect 42392 3476 42398 3528
rect 27062 3448 27068 3460
rect 27023 3420 27068 3448
rect 27062 3408 27068 3420
rect 27120 3408 27126 3460
rect 27338 3408 27344 3460
rect 27396 3448 27402 3460
rect 32398 3448 32404 3460
rect 27396 3420 32404 3448
rect 27396 3408 27402 3420
rect 32398 3408 32404 3420
rect 32456 3408 32462 3460
rect 37274 3408 37280 3460
rect 37332 3448 37338 3460
rect 37553 3451 37611 3457
rect 37553 3448 37565 3451
rect 37332 3420 37565 3448
rect 37332 3408 37338 3420
rect 37553 3417 37565 3420
rect 37599 3417 37611 3451
rect 37553 3411 37611 3417
rect 42978 3408 42984 3460
rect 43036 3448 43042 3460
rect 43349 3451 43407 3457
rect 43349 3448 43361 3451
rect 43036 3420 43361 3448
rect 43036 3408 43042 3420
rect 43349 3417 43361 3420
rect 43395 3417 43407 3451
rect 43349 3411 43407 3417
rect 44085 3451 44143 3457
rect 44085 3417 44097 3451
rect 44131 3448 44143 3451
rect 44450 3448 44456 3460
rect 44131 3420 44456 3448
rect 44131 3417 44143 3420
rect 44085 3411 44143 3417
rect 44450 3408 44456 3420
rect 44508 3408 44514 3460
rect 24397 3383 24455 3389
rect 24397 3380 24409 3383
rect 23308 3352 24409 3380
rect 23201 3343 23259 3349
rect 24397 3349 24409 3352
rect 24443 3349 24455 3383
rect 24397 3343 24455 3349
rect 24578 3340 24584 3392
rect 24636 3380 24642 3392
rect 24854 3380 24860 3392
rect 24636 3352 24860 3380
rect 24636 3340 24642 3352
rect 24854 3340 24860 3352
rect 24912 3340 24918 3392
rect 25682 3380 25688 3392
rect 25643 3352 25688 3380
rect 25682 3340 25688 3352
rect 25740 3340 25746 3392
rect 26234 3340 26240 3392
rect 26292 3380 26298 3392
rect 26329 3383 26387 3389
rect 26329 3380 26341 3383
rect 26292 3352 26341 3380
rect 26292 3340 26298 3352
rect 26329 3349 26341 3352
rect 26375 3349 26387 3383
rect 26329 3343 26387 3349
rect 28166 3340 28172 3392
rect 28224 3380 28230 3392
rect 28721 3383 28779 3389
rect 28721 3380 28733 3383
rect 28224 3352 28733 3380
rect 28224 3340 28230 3352
rect 28721 3349 28733 3352
rect 28767 3349 28779 3383
rect 28721 3343 28779 3349
rect 29086 3340 29092 3392
rect 29144 3380 29150 3392
rect 29733 3383 29791 3389
rect 29733 3380 29745 3383
rect 29144 3352 29745 3380
rect 29144 3340 29150 3352
rect 29733 3349 29745 3352
rect 29779 3349 29791 3383
rect 29733 3343 29791 3349
rect 30006 3340 30012 3392
rect 30064 3380 30070 3392
rect 30469 3383 30527 3389
rect 30469 3380 30481 3383
rect 30064 3352 30481 3380
rect 30064 3340 30070 3352
rect 30469 3349 30481 3352
rect 30515 3349 30527 3383
rect 30469 3343 30527 3349
rect 30926 3340 30932 3392
rect 30984 3380 30990 3392
rect 31205 3383 31263 3389
rect 31205 3380 31217 3383
rect 30984 3352 31217 3380
rect 30984 3340 30990 3352
rect 31205 3349 31217 3352
rect 31251 3349 31263 3383
rect 31205 3343 31263 3349
rect 31846 3340 31852 3392
rect 31904 3380 31910 3392
rect 32125 3383 32183 3389
rect 32125 3380 32137 3383
rect 31904 3352 32137 3380
rect 31904 3340 31910 3352
rect 32125 3349 32137 3352
rect 32171 3349 32183 3383
rect 32125 3343 32183 3349
rect 32858 3340 32864 3392
rect 32916 3380 32922 3392
rect 33137 3383 33195 3389
rect 33137 3380 33149 3383
rect 32916 3352 33149 3380
rect 32916 3340 32922 3352
rect 33137 3349 33149 3352
rect 33183 3349 33195 3383
rect 33137 3343 33195 3349
rect 33778 3340 33784 3392
rect 33836 3380 33842 3392
rect 34057 3383 34115 3389
rect 34057 3380 34069 3383
rect 33836 3352 34069 3380
rect 33836 3340 33842 3352
rect 34057 3349 34069 3352
rect 34103 3349 34115 3383
rect 34057 3343 34115 3349
rect 34698 3340 34704 3392
rect 34756 3380 34762 3392
rect 34977 3383 35035 3389
rect 34977 3380 34989 3383
rect 34756 3352 34989 3380
rect 34756 3340 34762 3352
rect 34977 3349 34989 3352
rect 35023 3349 35035 3383
rect 34977 3343 35035 3349
rect 35618 3340 35624 3392
rect 35676 3380 35682 3392
rect 35897 3383 35955 3389
rect 35897 3380 35909 3383
rect 35676 3352 35909 3380
rect 35676 3340 35682 3352
rect 35897 3349 35909 3352
rect 35943 3349 35955 3383
rect 35897 3343 35955 3349
rect 36630 3340 36636 3392
rect 36688 3380 36694 3392
rect 36817 3383 36875 3389
rect 36817 3380 36829 3383
rect 36688 3352 36829 3380
rect 36688 3340 36694 3352
rect 36817 3349 36829 3352
rect 36863 3349 36875 3383
rect 36817 3343 36875 3349
rect 37642 3340 37648 3392
rect 37700 3380 37706 3392
rect 38289 3383 38347 3389
rect 38289 3380 38301 3383
rect 37700 3352 38301 3380
rect 37700 3340 37706 3352
rect 38289 3349 38301 3352
rect 38335 3349 38347 3383
rect 38289 3343 38347 3349
rect 38470 3340 38476 3392
rect 38528 3380 38534 3392
rect 38933 3383 38991 3389
rect 38933 3380 38945 3383
rect 38528 3352 38945 3380
rect 38528 3340 38534 3352
rect 38933 3349 38945 3352
rect 38979 3349 38991 3383
rect 38933 3343 38991 3349
rect 39482 3340 39488 3392
rect 39540 3380 39546 3392
rect 40037 3383 40095 3389
rect 40037 3380 40049 3383
rect 39540 3352 40049 3380
rect 39540 3340 39546 3352
rect 40037 3349 40049 3352
rect 40083 3349 40095 3383
rect 40678 3380 40684 3392
rect 40639 3352 40684 3380
rect 40037 3343 40095 3349
rect 40678 3340 40684 3352
rect 40736 3340 40742 3392
rect 41322 3340 41328 3392
rect 41380 3380 41386 3392
rect 41785 3383 41843 3389
rect 41785 3380 41797 3383
rect 41380 3352 41797 3380
rect 41380 3340 41386 3352
rect 41785 3349 41797 3352
rect 41831 3349 41843 3383
rect 41785 3343 41843 3349
rect 42242 3340 42248 3392
rect 42300 3380 42306 3392
rect 42521 3383 42579 3389
rect 42521 3380 42533 3383
rect 42300 3352 42533 3380
rect 42300 3340 42306 3352
rect 42521 3349 42533 3352
rect 42567 3349 42579 3383
rect 42521 3343 42579 3349
rect 1104 3290 44896 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 44896 3290
rect 1104 3216 44896 3238
rect 4062 3176 4068 3188
rect 2746 3148 4068 3176
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 2746 3040 2774 3148
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 11882 3176 11888 3188
rect 4203 3148 11888 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 12250 3136 12256 3188
rect 12308 3136 12314 3188
rect 14366 3176 14372 3188
rect 14327 3148 14372 3176
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 14550 3136 14556 3188
rect 14608 3176 14614 3188
rect 15013 3179 15071 3185
rect 15013 3176 15025 3179
rect 14608 3148 15025 3176
rect 14608 3136 14614 3148
rect 15013 3145 15025 3148
rect 15059 3145 15071 3179
rect 17770 3176 17776 3188
rect 15013 3139 15071 3145
rect 15120 3148 16528 3176
rect 17731 3148 17776 3176
rect 4706 3108 4712 3120
rect 3528 3080 4712 3108
rect 1995 3012 2774 3040
rect 3237 3043 3295 3049
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 3237 3009 3249 3043
rect 3283 3040 3295 3043
rect 3418 3040 3424 3052
rect 3283 3012 3424 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 3418 3000 3424 3012
rect 3476 3000 3482 3052
rect 382 2932 388 2984
rect 440 2972 446 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 440 2944 2237 2972
rect 440 2932 446 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 2240 2836 2268 2935
rect 2314 2932 2320 2984
rect 2372 2972 2378 2984
rect 3528 2981 3556 3080
rect 4706 3068 4712 3080
rect 4764 3068 4770 3120
rect 12268 3108 12296 3136
rect 5644 3080 12296 3108
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 2372 2944 3525 2972
rect 2372 2932 2378 2944
rect 3513 2941 3525 2944
rect 3559 2941 3571 2975
rect 3513 2935 3571 2941
rect 3988 2972 4016 3003
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 4120 3012 4629 3040
rect 4120 3000 4126 3012
rect 4617 3009 4629 3012
rect 4663 3040 4675 3043
rect 4890 3040 4896 3052
rect 4663 3012 4896 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 5537 3043 5595 3049
rect 5537 3040 5549 3043
rect 5500 3012 5549 3040
rect 5500 3000 5506 3012
rect 5537 3009 5549 3012
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 4706 2972 4712 2984
rect 3988 2944 4712 2972
rect 2590 2864 2596 2916
rect 2648 2904 2654 2916
rect 3988 2904 4016 2944
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 5534 2904 5540 2916
rect 2648 2876 4016 2904
rect 4080 2876 5540 2904
rect 2648 2864 2654 2876
rect 4080 2836 4108 2876
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 2240 2808 4108 2836
rect 4801 2839 4859 2845
rect 4801 2805 4813 2839
rect 4847 2836 4859 2839
rect 5644 2836 5672 3080
rect 13078 3068 13084 3120
rect 13136 3108 13142 3120
rect 15120 3108 15148 3148
rect 16390 3108 16396 3120
rect 13136 3080 15148 3108
rect 15212 3080 16396 3108
rect 13136 3068 13142 3080
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 6788 3012 7573 3040
rect 6788 3000 6794 3012
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 8570 3040 8576 3052
rect 8531 3012 8576 3040
rect 7561 3003 7619 3009
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 8938 3000 8944 3052
rect 8996 3040 9002 3052
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 8996 3012 9321 3040
rect 8996 3000 9002 3012
rect 9309 3009 9321 3012
rect 9355 3040 9367 3043
rect 9674 3040 9680 3052
rect 9355 3012 9680 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 10502 3040 10508 3052
rect 10463 3012 10508 3040
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 10778 3040 10784 3052
rect 10739 3012 10784 3040
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 12250 3040 12256 3052
rect 12211 3012 12256 3040
rect 11793 3003 11851 3009
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2941 7343 2975
rect 8846 2972 8852 2984
rect 8807 2944 8852 2972
rect 7285 2935 7343 2941
rect 5721 2907 5779 2913
rect 5721 2873 5733 2907
rect 5767 2904 5779 2907
rect 6914 2904 6920 2916
rect 5767 2876 6920 2904
rect 5767 2873 5779 2876
rect 5721 2867 5779 2873
rect 6914 2864 6920 2876
rect 6972 2864 6978 2916
rect 7300 2904 7328 2935
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 10796 2972 10824 3000
rect 9916 2944 10824 2972
rect 9916 2932 9922 2944
rect 11808 2904 11836 3003
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 12912 2972 12940 3003
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 13541 3043 13599 3049
rect 13541 3040 13553 3043
rect 13320 3012 13553 3040
rect 13320 3000 13326 3012
rect 13541 3009 13553 3012
rect 13587 3009 13599 3043
rect 13541 3003 13599 3009
rect 14274 3000 14280 3052
rect 14332 3040 14338 3052
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 14332 3012 14565 3040
rect 14332 3000 14338 3012
rect 14553 3009 14565 3012
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 14642 3000 14648 3052
rect 14700 3040 14706 3052
rect 15212 3049 15240 3080
rect 16390 3068 16396 3080
rect 16448 3068 16454 3120
rect 16500 3108 16528 3148
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18233 3179 18291 3185
rect 18233 3176 18245 3179
rect 18012 3148 18245 3176
rect 18012 3136 18018 3148
rect 18233 3145 18245 3148
rect 18279 3145 18291 3179
rect 20165 3179 20223 3185
rect 18233 3139 18291 3145
rect 18340 3148 19564 3176
rect 16500 3080 17954 3108
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 14700 3012 15209 3040
rect 14700 3000 14706 3012
rect 15197 3009 15209 3012
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 16114 3040 16120 3052
rect 15979 3012 16120 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3009 17647 3043
rect 17926 3040 17954 3080
rect 18340 3040 18368 3148
rect 19536 3108 19564 3148
rect 20165 3145 20177 3179
rect 20211 3176 20223 3179
rect 20530 3176 20536 3188
rect 20211 3148 20536 3176
rect 20211 3145 20223 3148
rect 20165 3139 20223 3145
rect 20530 3136 20536 3148
rect 20588 3136 20594 3188
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 20993 3179 21051 3185
rect 20993 3176 21005 3179
rect 20956 3148 21005 3176
rect 20956 3136 20962 3148
rect 20993 3145 21005 3148
rect 21039 3145 21051 3179
rect 20993 3139 21051 3145
rect 21818 3136 21824 3188
rect 21876 3176 21882 3188
rect 21913 3179 21971 3185
rect 21913 3176 21925 3179
rect 21876 3148 21925 3176
rect 21876 3136 21882 3148
rect 21913 3145 21925 3148
rect 21959 3145 21971 3179
rect 22830 3176 22836 3188
rect 22791 3148 22836 3176
rect 21913 3139 21971 3145
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 23106 3136 23112 3188
rect 23164 3176 23170 3188
rect 23290 3176 23296 3188
rect 23164 3148 23296 3176
rect 23164 3136 23170 3148
rect 23290 3136 23296 3148
rect 23348 3136 23354 3188
rect 23753 3179 23811 3185
rect 23753 3145 23765 3179
rect 23799 3176 23811 3179
rect 23842 3176 23848 3188
rect 23799 3148 23848 3176
rect 23799 3145 23811 3148
rect 23753 3139 23811 3145
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 24210 3136 24216 3188
rect 24268 3176 24274 3188
rect 24581 3179 24639 3185
rect 24581 3176 24593 3179
rect 24268 3148 24593 3176
rect 24268 3136 24274 3148
rect 24581 3145 24593 3148
rect 24627 3145 24639 3179
rect 24581 3139 24639 3145
rect 26878 3136 26884 3188
rect 26936 3176 26942 3188
rect 27062 3176 27068 3188
rect 26936 3148 27068 3176
rect 26936 3136 26942 3148
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 27522 3136 27528 3188
rect 27580 3176 27586 3188
rect 32585 3179 32643 3185
rect 32585 3176 32597 3179
rect 27580 3148 32597 3176
rect 27580 3136 27586 3148
rect 32585 3145 32597 3148
rect 32631 3145 32643 3179
rect 32585 3139 32643 3145
rect 32766 3136 32772 3188
rect 32824 3176 32830 3188
rect 34057 3179 34115 3185
rect 34057 3176 34069 3179
rect 32824 3148 34069 3176
rect 32824 3136 32830 3148
rect 34057 3145 34069 3148
rect 34103 3145 34115 3179
rect 35526 3176 35532 3188
rect 35487 3148 35532 3176
rect 34057 3139 34115 3145
rect 35526 3136 35532 3148
rect 35584 3136 35590 3188
rect 37366 3176 37372 3188
rect 37327 3148 37372 3176
rect 37366 3136 37372 3148
rect 37424 3136 37430 3188
rect 43990 3176 43996 3188
rect 43951 3148 43996 3176
rect 43990 3136 43996 3148
rect 44048 3136 44054 3188
rect 20714 3108 20720 3120
rect 19536 3080 20720 3108
rect 20714 3068 20720 3080
rect 20772 3068 20778 3120
rect 22370 3108 22376 3120
rect 21192 3080 22376 3108
rect 19058 3040 19064 3052
rect 17926 3012 18368 3040
rect 19019 3012 19064 3040
rect 17589 3003 17647 3009
rect 13814 2972 13820 2984
rect 12400 2944 13820 2972
rect 12400 2932 12406 2944
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 17034 2932 17040 2984
rect 17092 2972 17098 2984
rect 17604 2972 17632 3003
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 19978 3040 19984 3052
rect 19891 3012 19984 3040
rect 19978 3000 19984 3012
rect 20036 3040 20042 3052
rect 20622 3040 20628 3052
rect 20036 3012 20628 3040
rect 20036 3000 20042 3012
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 20898 3000 20904 3052
rect 20956 3040 20962 3052
rect 21192 3049 21220 3080
rect 22370 3068 22376 3080
rect 22428 3068 22434 3120
rect 25038 3108 25044 3120
rect 23952 3080 25044 3108
rect 21177 3043 21235 3049
rect 21177 3040 21189 3043
rect 20956 3012 21189 3040
rect 20956 3000 20962 3012
rect 21177 3009 21189 3012
rect 21223 3009 21235 3043
rect 21177 3003 21235 3009
rect 21818 3000 21824 3052
rect 21876 3040 21882 3052
rect 22097 3043 22155 3049
rect 22097 3040 22109 3043
rect 21876 3012 22109 3040
rect 21876 3000 21882 3012
rect 22097 3009 22109 3012
rect 22143 3040 22155 3043
rect 22186 3040 22192 3052
rect 22143 3012 22192 3040
rect 22143 3009 22155 3012
rect 22097 3003 22155 3009
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 22738 3000 22744 3052
rect 22796 3040 22802 3052
rect 23014 3040 23020 3052
rect 22796 3012 23020 3040
rect 22796 3000 22802 3012
rect 23014 3000 23020 3012
rect 23072 3000 23078 3052
rect 23658 3000 23664 3052
rect 23716 3040 23722 3052
rect 23952 3049 23980 3080
rect 25038 3068 25044 3080
rect 25096 3068 25102 3120
rect 25866 3068 25872 3120
rect 25924 3108 25930 3120
rect 26053 3111 26111 3117
rect 26053 3108 26065 3111
rect 25924 3080 26065 3108
rect 25924 3068 25930 3080
rect 26053 3077 26065 3080
rect 26099 3108 26111 3111
rect 26142 3108 26148 3120
rect 26099 3080 26148 3108
rect 26099 3077 26111 3080
rect 26053 3071 26111 3077
rect 26142 3068 26148 3080
rect 26200 3068 26206 3120
rect 26237 3111 26295 3117
rect 26237 3077 26249 3111
rect 26283 3108 26295 3111
rect 27338 3108 27344 3120
rect 26283 3080 27344 3108
rect 26283 3077 26295 3080
rect 26237 3071 26295 3077
rect 27338 3068 27344 3080
rect 27396 3068 27402 3120
rect 27430 3068 27436 3120
rect 27488 3108 27494 3120
rect 27617 3111 27675 3117
rect 27617 3108 27629 3111
rect 27488 3080 27629 3108
rect 27488 3068 27494 3080
rect 27617 3077 27629 3080
rect 27663 3108 27675 3111
rect 27706 3108 27712 3120
rect 27663 3080 27712 3108
rect 27663 3077 27675 3080
rect 27617 3071 27675 3077
rect 27706 3068 27712 3080
rect 27764 3068 27770 3120
rect 27801 3111 27859 3117
rect 27801 3077 27813 3111
rect 27847 3108 27859 3111
rect 28442 3108 28448 3120
rect 27847 3080 28448 3108
rect 27847 3077 27859 3080
rect 27801 3071 27859 3077
rect 28442 3068 28448 3080
rect 28500 3068 28506 3120
rect 29638 3068 29644 3120
rect 29696 3108 29702 3120
rect 30282 3108 30288 3120
rect 29696 3080 30288 3108
rect 29696 3068 29702 3080
rect 30282 3068 30288 3080
rect 30340 3068 30346 3120
rect 30650 3068 30656 3120
rect 30708 3108 30714 3120
rect 31021 3111 31079 3117
rect 31021 3108 31033 3111
rect 30708 3080 31033 3108
rect 30708 3068 30714 3080
rect 31021 3077 31033 3080
rect 31067 3108 31079 3111
rect 31202 3108 31208 3120
rect 31067 3080 31208 3108
rect 31067 3077 31079 3080
rect 31021 3071 31079 3077
rect 31202 3068 31208 3080
rect 31260 3068 31266 3120
rect 32490 3068 32496 3120
rect 32548 3108 32554 3120
rect 33042 3108 33048 3120
rect 32548 3080 33048 3108
rect 32548 3068 32554 3080
rect 33042 3068 33048 3080
rect 33100 3108 33106 3120
rect 33413 3111 33471 3117
rect 33413 3108 33425 3111
rect 33100 3080 33425 3108
rect 33100 3068 33106 3080
rect 33413 3077 33425 3080
rect 33459 3077 33471 3111
rect 33413 3071 33471 3077
rect 34514 3068 34520 3120
rect 34572 3108 34578 3120
rect 34701 3111 34759 3117
rect 34701 3108 34713 3111
rect 34572 3080 34713 3108
rect 34572 3068 34578 3080
rect 34701 3077 34713 3080
rect 34747 3077 34759 3111
rect 34701 3071 34759 3077
rect 35986 3068 35992 3120
rect 36044 3108 36050 3120
rect 37182 3108 37188 3120
rect 36044 3080 37188 3108
rect 36044 3068 36050 3080
rect 37182 3068 37188 3080
rect 37240 3108 37246 3120
rect 37461 3111 37519 3117
rect 37461 3108 37473 3111
rect 37240 3080 37473 3108
rect 37240 3068 37246 3080
rect 37461 3077 37473 3080
rect 37507 3077 37519 3111
rect 38010 3108 38016 3120
rect 37971 3080 38016 3108
rect 37461 3071 37519 3077
rect 38010 3068 38016 3080
rect 38068 3068 38074 3120
rect 39390 3068 39396 3120
rect 39448 3108 39454 3120
rect 39485 3111 39543 3117
rect 39485 3108 39497 3111
rect 39448 3080 39497 3108
rect 39448 3068 39454 3080
rect 39485 3077 39497 3080
rect 39531 3077 39543 3111
rect 40218 3108 40224 3120
rect 40179 3080 40224 3108
rect 39485 3071 39543 3077
rect 40218 3068 40224 3080
rect 40276 3068 40282 3120
rect 42794 3108 42800 3120
rect 42755 3080 42800 3108
rect 42794 3068 42800 3080
rect 42852 3068 42858 3120
rect 43162 3068 43168 3120
rect 43220 3108 43226 3120
rect 43530 3108 43536 3120
rect 43220 3080 43536 3108
rect 43220 3068 43226 3080
rect 43530 3068 43536 3080
rect 43588 3108 43594 3120
rect 44085 3111 44143 3117
rect 44085 3108 44097 3111
rect 43588 3080 44097 3108
rect 43588 3068 43594 3080
rect 44085 3077 44097 3080
rect 44131 3077 44143 3111
rect 44085 3071 44143 3077
rect 23937 3043 23995 3049
rect 23937 3040 23949 3043
rect 23716 3012 23949 3040
rect 23716 3000 23722 3012
rect 23937 3009 23949 3012
rect 23983 3009 23995 3043
rect 23937 3003 23995 3009
rect 24765 3043 24823 3049
rect 24765 3009 24777 3043
rect 24811 3009 24823 3043
rect 24765 3003 24823 3009
rect 25501 3043 25559 3049
rect 25501 3009 25513 3043
rect 25547 3040 25559 3043
rect 25774 3040 25780 3052
rect 25547 3012 25780 3040
rect 25547 3009 25559 3012
rect 25501 3003 25559 3009
rect 24578 2972 24584 2984
rect 17092 2944 24584 2972
rect 17092 2932 17098 2944
rect 24578 2932 24584 2944
rect 24636 2932 24642 2984
rect 24670 2932 24676 2984
rect 24728 2972 24734 2984
rect 24780 2972 24808 3003
rect 25774 3000 25780 3012
rect 25832 3000 25838 3052
rect 26694 3000 26700 3052
rect 26752 3040 26758 3052
rect 26752 3012 27476 3040
rect 26752 3000 26758 3012
rect 24728 2944 24808 2972
rect 24728 2932 24734 2944
rect 26786 2932 26792 2984
rect 26844 2972 26850 2984
rect 27338 2972 27344 2984
rect 26844 2944 27344 2972
rect 26844 2932 26850 2944
rect 27338 2932 27344 2944
rect 27396 2932 27402 2984
rect 27448 2972 27476 3012
rect 28718 3000 28724 3052
rect 28776 3040 28782 3052
rect 28813 3043 28871 3049
rect 28813 3040 28825 3043
rect 28776 3012 28825 3040
rect 28776 3000 28782 3012
rect 28813 3009 28825 3012
rect 28859 3009 28871 3043
rect 28813 3003 28871 3009
rect 28902 3000 28908 3052
rect 28960 3040 28966 3052
rect 30101 3043 30159 3049
rect 30101 3040 30113 3043
rect 28960 3012 30113 3040
rect 28960 3000 28966 3012
rect 30101 3009 30113 3012
rect 30147 3009 30159 3043
rect 30101 3003 30159 3009
rect 30190 3000 30196 3052
rect 30248 3040 30254 3052
rect 30837 3043 30895 3049
rect 30837 3040 30849 3043
rect 30248 3012 30849 3040
rect 30248 3000 30254 3012
rect 30837 3009 30849 3012
rect 30883 3009 30895 3043
rect 30837 3003 30895 3009
rect 31662 3000 31668 3052
rect 31720 3040 31726 3052
rect 32677 3043 32735 3049
rect 32677 3040 32689 3043
rect 31720 3012 32689 3040
rect 31720 3000 31726 3012
rect 32677 3009 32689 3012
rect 32723 3009 32735 3043
rect 32677 3003 32735 3009
rect 33502 3000 33508 3052
rect 33560 3040 33566 3052
rect 34149 3043 34207 3049
rect 34149 3040 34161 3043
rect 33560 3012 34161 3040
rect 33560 3000 33566 3012
rect 34149 3009 34161 3012
rect 34195 3009 34207 3043
rect 34149 3003 34207 3009
rect 34422 3000 34428 3052
rect 34480 3040 34486 3052
rect 34790 3040 34796 3052
rect 34480 3012 34796 3040
rect 34480 3000 34486 3012
rect 34790 3000 34796 3012
rect 34848 3040 34854 3052
rect 34885 3043 34943 3049
rect 34885 3040 34897 3043
rect 34848 3012 34897 3040
rect 34848 3000 34854 3012
rect 34885 3009 34897 3012
rect 34931 3009 34943 3043
rect 34885 3003 34943 3009
rect 35342 3000 35348 3052
rect 35400 3040 35406 3052
rect 35621 3043 35679 3049
rect 35621 3040 35633 3043
rect 35400 3012 35633 3040
rect 35400 3000 35406 3012
rect 35621 3009 35633 3012
rect 35667 3009 35679 3043
rect 35621 3003 35679 3009
rect 36262 3000 36268 3052
rect 36320 3040 36326 3052
rect 36541 3043 36599 3049
rect 36541 3040 36553 3043
rect 36320 3012 36553 3040
rect 36320 3000 36326 3012
rect 36541 3009 36553 3012
rect 36587 3009 36599 3043
rect 36541 3003 36599 3009
rect 38197 3043 38255 3049
rect 38197 3009 38209 3043
rect 38243 3009 38255 3043
rect 38197 3003 38255 3009
rect 36357 2975 36415 2981
rect 36357 2972 36369 2975
rect 27448 2944 36369 2972
rect 36357 2941 36369 2944
rect 36403 2941 36415 2975
rect 36357 2935 36415 2941
rect 36906 2932 36912 2984
rect 36964 2972 36970 2984
rect 38212 2972 38240 3003
rect 38286 3000 38292 3052
rect 38344 3040 38350 3052
rect 38654 3040 38660 3052
rect 38344 3012 38660 3040
rect 38344 3000 38350 3012
rect 38654 3000 38660 3012
rect 38712 3040 38718 3052
rect 38933 3043 38991 3049
rect 38933 3040 38945 3043
rect 38712 3012 38945 3040
rect 38712 3000 38718 3012
rect 38933 3009 38945 3012
rect 38979 3009 38991 3043
rect 38933 3003 38991 3009
rect 39114 3000 39120 3052
rect 39172 3040 39178 3052
rect 39669 3043 39727 3049
rect 39669 3040 39681 3043
rect 39172 3012 39681 3040
rect 39172 3000 39178 3012
rect 39669 3009 39681 3012
rect 39715 3040 39727 3043
rect 39942 3040 39948 3052
rect 39715 3012 39948 3040
rect 39715 3009 39727 3012
rect 39669 3003 39727 3009
rect 39942 3000 39948 3012
rect 40000 3000 40006 3052
rect 40034 3000 40040 3052
rect 40092 3040 40098 3052
rect 40402 3040 40408 3052
rect 40092 3012 40408 3040
rect 40092 3000 40098 3012
rect 40402 3000 40408 3012
rect 40460 3000 40466 3052
rect 40770 3000 40776 3052
rect 40828 3040 40834 3052
rect 40957 3043 41015 3049
rect 40957 3040 40969 3043
rect 40828 3012 40969 3040
rect 40828 3000 40834 3012
rect 40957 3009 40969 3012
rect 41003 3009 41015 3043
rect 40957 3003 41015 3009
rect 41966 3000 41972 3052
rect 42024 3040 42030 3052
rect 42610 3040 42616 3052
rect 42024 3012 42616 3040
rect 42024 3000 42030 3012
rect 42610 3000 42616 3012
rect 42668 3040 42674 3052
rect 42981 3043 43039 3049
rect 42981 3040 42993 3043
rect 42668 3012 42993 3040
rect 42668 3000 42674 3012
rect 42981 3009 42993 3012
rect 43027 3009 43039 3043
rect 42981 3003 43039 3009
rect 36964 2944 38240 2972
rect 36964 2932 36970 2944
rect 7300 2876 11744 2904
rect 11808 2876 12572 2904
rect 4847 2808 5672 2836
rect 9493 2839 9551 2845
rect 4847 2805 4859 2808
rect 4801 2799 4859 2805
rect 9493 2805 9505 2839
rect 9539 2836 9551 2839
rect 9582 2836 9588 2848
rect 9539 2808 9588 2836
rect 9539 2805 9551 2808
rect 9493 2799 9551 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 11609 2839 11667 2845
rect 11609 2836 11621 2839
rect 11112 2808 11621 2836
rect 11112 2796 11118 2808
rect 11609 2805 11621 2808
rect 11655 2805 11667 2839
rect 11716 2836 11744 2876
rect 11882 2836 11888 2848
rect 11716 2808 11888 2836
rect 11609 2799 11667 2805
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 12434 2836 12440 2848
rect 12395 2808 12440 2836
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 12544 2836 12572 2876
rect 12710 2864 12716 2916
rect 12768 2904 12774 2916
rect 13081 2907 13139 2913
rect 13081 2904 13093 2907
rect 12768 2876 13093 2904
rect 12768 2864 12774 2876
rect 13081 2873 13093 2876
rect 13127 2873 13139 2907
rect 15746 2904 15752 2916
rect 13081 2867 13139 2873
rect 13188 2876 15752 2904
rect 13188 2836 13216 2876
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 16117 2907 16175 2913
rect 16117 2873 16129 2907
rect 16163 2904 16175 2907
rect 18046 2904 18052 2916
rect 16163 2876 18052 2904
rect 16163 2873 16175 2876
rect 16117 2867 16175 2873
rect 18046 2864 18052 2876
rect 18104 2864 18110 2916
rect 19886 2904 19892 2916
rect 18616 2876 19892 2904
rect 12544 2808 13216 2836
rect 13725 2839 13783 2845
rect 13725 2805 13737 2839
rect 13771 2836 13783 2839
rect 16666 2836 16672 2848
rect 13771 2808 16672 2836
rect 13771 2805 13783 2808
rect 13725 2799 13783 2805
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 16945 2839 17003 2845
rect 16945 2836 16957 2839
rect 16816 2808 16957 2836
rect 16816 2796 16822 2808
rect 16945 2805 16957 2808
rect 16991 2805 17003 2839
rect 16945 2799 17003 2805
rect 17586 2796 17592 2848
rect 17644 2836 17650 2848
rect 18616 2836 18644 2876
rect 19886 2864 19892 2876
rect 19944 2864 19950 2916
rect 22554 2864 22560 2916
rect 22612 2904 22618 2916
rect 33226 2904 33232 2916
rect 22612 2876 28488 2904
rect 33187 2876 33232 2904
rect 22612 2864 22618 2876
rect 17644 2808 18644 2836
rect 17644 2796 17650 2808
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 18877 2839 18935 2845
rect 18877 2836 18889 2839
rect 18748 2808 18889 2836
rect 18748 2796 18754 2808
rect 18877 2805 18889 2808
rect 18923 2805 18935 2839
rect 18877 2799 18935 2805
rect 25222 2796 25228 2848
rect 25280 2836 25286 2848
rect 25317 2839 25375 2845
rect 25317 2836 25329 2839
rect 25280 2808 25329 2836
rect 25280 2796 25286 2808
rect 25317 2805 25329 2808
rect 25363 2805 25375 2839
rect 25317 2799 25375 2805
rect 25774 2796 25780 2848
rect 25832 2836 25838 2848
rect 26418 2836 26424 2848
rect 25832 2808 26424 2836
rect 25832 2796 25838 2808
rect 26418 2796 26424 2808
rect 26476 2796 26482 2848
rect 28350 2836 28356 2848
rect 28311 2808 28356 2836
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 28460 2836 28488 2876
rect 33226 2864 33232 2876
rect 33284 2864 33290 2916
rect 34146 2864 34152 2916
rect 34204 2904 34210 2916
rect 38749 2907 38807 2913
rect 38749 2904 38761 2907
rect 34204 2876 38761 2904
rect 34204 2864 34210 2876
rect 38749 2873 38761 2876
rect 38795 2873 38807 2907
rect 38749 2867 38807 2873
rect 29043 2839 29101 2845
rect 29043 2836 29055 2839
rect 28460 2808 29055 2836
rect 29043 2805 29055 2808
rect 29089 2805 29101 2839
rect 29043 2799 29101 2805
rect 40402 2796 40408 2848
rect 40460 2836 40466 2848
rect 41141 2839 41199 2845
rect 41141 2836 41153 2839
rect 40460 2808 41153 2836
rect 40460 2796 40466 2808
rect 41141 2805 41153 2808
rect 41187 2805 41199 2839
rect 41141 2799 41199 2805
rect 41690 2796 41696 2848
rect 41748 2836 41754 2848
rect 41785 2839 41843 2845
rect 41785 2836 41797 2839
rect 41748 2808 41797 2836
rect 41748 2796 41754 2808
rect 41785 2805 41797 2808
rect 41831 2836 41843 2839
rect 42794 2836 42800 2848
rect 41831 2808 42800 2836
rect 41831 2805 41843 2808
rect 41785 2799 41843 2805
rect 42794 2796 42800 2808
rect 42852 2796 42858 2848
rect 1104 2746 44896 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 44896 2746
rect 1104 2672 44896 2694
rect 4249 2635 4307 2641
rect 4249 2601 4261 2635
rect 4295 2632 4307 2635
rect 5258 2632 5264 2644
rect 4295 2604 5264 2632
rect 4295 2601 4307 2604
rect 4249 2595 4307 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8570 2632 8576 2644
rect 8352 2604 8576 2632
rect 8352 2592 8358 2604
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9490 2632 9496 2644
rect 9171 2604 9496 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 19886 2592 19892 2644
rect 19944 2632 19950 2644
rect 32585 2635 32643 2641
rect 32585 2632 32597 2635
rect 19944 2604 32597 2632
rect 19944 2592 19950 2604
rect 32585 2601 32597 2604
rect 32631 2601 32643 2635
rect 32585 2595 32643 2601
rect 33686 2592 33692 2644
rect 33744 2632 33750 2644
rect 38013 2635 38071 2641
rect 38013 2632 38025 2635
rect 33744 2604 38025 2632
rect 33744 2592 33750 2604
rect 38013 2601 38025 2604
rect 38059 2601 38071 2635
rect 38013 2595 38071 2601
rect 2682 2564 2688 2576
rect 2643 2536 2688 2564
rect 2682 2524 2688 2536
rect 2740 2524 2746 2576
rect 5721 2567 5779 2573
rect 5721 2533 5733 2567
rect 5767 2564 5779 2567
rect 8110 2564 8116 2576
rect 5767 2536 8116 2564
rect 5767 2533 5779 2536
rect 5721 2527 5779 2533
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 8389 2567 8447 2573
rect 8389 2533 8401 2567
rect 8435 2564 8447 2567
rect 11146 2564 11152 2576
rect 8435 2536 11152 2564
rect 8435 2533 8447 2536
rect 8389 2527 8447 2533
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 17770 2564 17776 2576
rect 17731 2536 17776 2564
rect 17770 2524 17776 2536
rect 17828 2524 17834 2576
rect 19996 2536 26234 2564
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 5350 2496 5356 2508
rect 1995 2468 5356 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 5350 2456 5356 2468
rect 5408 2456 5414 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6886 2468 7297 2496
rect 6886 2440 6914 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 9582 2496 9588 2508
rect 7285 2459 7343 2465
rect 8128 2468 9588 2496
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2774 2428 2780 2440
rect 2271 2400 2780 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 4430 2388 4436 2440
rect 4488 2428 4494 2440
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4488 2400 4905 2428
rect 4488 2388 4494 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5074 2388 5080 2440
rect 5132 2428 5138 2440
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 5132 2400 5549 2428
rect 5132 2388 5138 2400
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 6822 2388 6828 2440
rect 6880 2400 6914 2440
rect 6880 2388 6886 2400
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7064 2400 7109 2428
rect 7064 2388 7070 2400
rect 2866 2360 2872 2372
rect 2827 2332 2872 2360
rect 2866 2320 2872 2332
rect 2924 2320 2930 2372
rect 4062 2320 4068 2372
rect 4120 2360 4126 2372
rect 4341 2363 4399 2369
rect 4341 2360 4353 2363
rect 4120 2332 4353 2360
rect 4120 2320 4126 2332
rect 4341 2329 4353 2332
rect 4387 2360 4399 2363
rect 8128 2360 8156 2468
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 10134 2496 10140 2508
rect 10095 2468 10140 2496
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 10413 2499 10471 2505
rect 10413 2465 10425 2499
rect 10459 2496 10471 2499
rect 11422 2496 11428 2508
rect 10459 2468 11428 2496
rect 10459 2465 10471 2468
rect 10413 2459 10471 2465
rect 8202 2388 8208 2440
rect 8260 2428 8266 2440
rect 8260 2400 8305 2428
rect 8260 2388 8266 2400
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8536 2400 8953 2428
rect 8536 2388 8542 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9490 2388 9496 2440
rect 9548 2428 9554 2440
rect 10428 2428 10456 2459
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 11882 2456 11888 2508
rect 11940 2496 11946 2508
rect 17494 2496 17500 2508
rect 11940 2468 17500 2496
rect 11940 2456 11946 2468
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 9548 2400 10456 2428
rect 11793 2431 11851 2437
rect 9548 2388 9554 2400
rect 11793 2397 11805 2431
rect 11839 2428 11851 2431
rect 12434 2428 12440 2440
rect 11839 2400 12440 2428
rect 11839 2397 11851 2400
rect 11793 2391 11851 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12986 2428 12992 2440
rect 12575 2400 12992 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2428 13415 2431
rect 13998 2428 14004 2440
rect 13403 2400 14004 2428
rect 13403 2397 13415 2400
rect 13357 2391 13415 2397
rect 13998 2388 14004 2400
rect 14056 2388 14062 2440
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2428 15255 2431
rect 15562 2428 15568 2440
rect 15243 2400 15568 2428
rect 15243 2397 15255 2400
rect 15197 2391 15255 2397
rect 10873 2363 10931 2369
rect 10873 2360 10885 2363
rect 4387 2332 8156 2360
rect 8312 2332 10885 2360
rect 4387 2329 4399 2332
rect 4341 2323 4399 2329
rect 6362 2252 6368 2304
rect 6420 2292 6426 2304
rect 8312 2292 8340 2332
rect 10873 2329 10885 2332
rect 10919 2329 10931 2363
rect 14384 2360 14412 2391
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2428 15715 2431
rect 15930 2428 15936 2440
rect 15703 2400 15936 2428
rect 15703 2397 15715 2400
rect 15657 2391 15715 2397
rect 15470 2360 15476 2372
rect 14384 2332 15476 2360
rect 10873 2323 10931 2329
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 6420 2264 8340 2292
rect 6420 2252 6426 2264
rect 10134 2252 10140 2304
rect 10192 2292 10198 2304
rect 11609 2295 11667 2301
rect 11609 2292 11621 2295
rect 10192 2264 11621 2292
rect 10192 2252 10198 2264
rect 11609 2261 11621 2264
rect 11655 2261 11667 2295
rect 11609 2255 11667 2261
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 12124 2264 12357 2292
rect 12124 2252 12130 2264
rect 12345 2261 12357 2264
rect 12391 2261 12403 2295
rect 12345 2255 12403 2261
rect 12986 2252 12992 2304
rect 13044 2292 13050 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 13044 2264 13185 2292
rect 13044 2252 13050 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 13906 2252 13912 2304
rect 13964 2292 13970 2304
rect 14185 2295 14243 2301
rect 14185 2292 14197 2295
rect 13964 2264 14197 2292
rect 13964 2252 13970 2264
rect 14185 2261 14197 2264
rect 14231 2261 14243 2295
rect 14185 2255 14243 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14884 2264 15025 2292
rect 14884 2252 14890 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 15672 2292 15700 2391
rect 15930 2388 15936 2400
rect 15988 2388 15994 2440
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2428 17003 2431
rect 17218 2428 17224 2440
rect 16991 2400 17224 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 18506 2428 18512 2440
rect 18467 2400 18512 2428
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 19996 2437 20024 2536
rect 25958 2496 25964 2508
rect 25919 2468 25964 2496
rect 25958 2456 25964 2468
rect 26016 2456 26022 2508
rect 19981 2431 20039 2437
rect 19981 2397 19993 2431
rect 20027 2397 20039 2431
rect 19981 2391 20039 2397
rect 20806 2388 20812 2440
rect 20864 2428 20870 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20864 2400 20913 2428
rect 20864 2388 20870 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 21726 2388 21732 2440
rect 21784 2428 21790 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 21784 2400 21833 2428
rect 21784 2388 21790 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2428 22891 2431
rect 23474 2428 23480 2440
rect 22879 2400 23480 2428
rect 22879 2397 22891 2400
rect 22833 2391 22891 2397
rect 23474 2388 23480 2400
rect 23532 2388 23538 2440
rect 23750 2428 23756 2440
rect 23711 2400 23756 2428
rect 23750 2388 23756 2400
rect 23808 2388 23814 2440
rect 24302 2388 24308 2440
rect 24360 2428 24366 2440
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 24360 2400 24409 2428
rect 24360 2388 24366 2400
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 25590 2388 25596 2440
rect 25648 2428 25654 2440
rect 25774 2428 25780 2440
rect 25648 2400 25780 2428
rect 25648 2388 25654 2400
rect 25774 2388 25780 2400
rect 25832 2388 25838 2440
rect 17402 2320 17408 2372
rect 17460 2360 17466 2372
rect 17589 2363 17647 2369
rect 17589 2360 17601 2363
rect 17460 2332 17601 2360
rect 17460 2320 17466 2332
rect 17589 2329 17601 2332
rect 17635 2360 17647 2363
rect 21082 2360 21088 2372
rect 17635 2332 21088 2360
rect 17635 2329 17647 2332
rect 17589 2323 17647 2329
rect 21082 2320 21088 2332
rect 21140 2320 21146 2372
rect 15838 2292 15844 2304
rect 15252 2264 15700 2292
rect 15799 2264 15844 2292
rect 15252 2252 15258 2264
rect 15838 2252 15844 2264
rect 15896 2252 15902 2304
rect 15930 2252 15936 2304
rect 15988 2292 15994 2304
rect 16761 2295 16819 2301
rect 16761 2292 16773 2295
rect 15988 2264 16773 2292
rect 15988 2252 15994 2264
rect 16761 2261 16773 2264
rect 16807 2261 16819 2295
rect 16761 2255 16819 2261
rect 17770 2252 17776 2304
rect 17828 2292 17834 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 17828 2264 18337 2292
rect 17828 2252 17834 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 19426 2252 19432 2304
rect 19484 2292 19490 2304
rect 19797 2295 19855 2301
rect 19797 2292 19809 2295
rect 19484 2264 19809 2292
rect 19484 2252 19490 2264
rect 19797 2261 19809 2264
rect 19843 2261 19855 2295
rect 19797 2255 19855 2261
rect 20530 2252 20536 2304
rect 20588 2292 20594 2304
rect 20717 2295 20775 2301
rect 20717 2292 20729 2295
rect 20588 2264 20729 2292
rect 20588 2252 20594 2264
rect 20717 2261 20729 2264
rect 20763 2261 20775 2295
rect 20717 2255 20775 2261
rect 21450 2252 21456 2304
rect 21508 2292 21514 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21508 2264 22017 2292
rect 21508 2252 21514 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 22462 2252 22468 2304
rect 22520 2292 22526 2304
rect 22649 2295 22707 2301
rect 22649 2292 22661 2295
rect 22520 2264 22661 2292
rect 22520 2252 22526 2264
rect 22649 2261 22661 2264
rect 22695 2261 22707 2295
rect 22649 2255 22707 2261
rect 23382 2252 23388 2304
rect 23440 2292 23446 2304
rect 23569 2295 23627 2301
rect 23569 2292 23581 2295
rect 23440 2264 23581 2292
rect 23440 2252 23446 2264
rect 23569 2261 23581 2264
rect 23615 2261 23627 2295
rect 23569 2255 23627 2261
rect 24302 2252 24308 2304
rect 24360 2292 24366 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24360 2264 24593 2292
rect 24360 2252 24366 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 25130 2292 25136 2304
rect 25091 2264 25136 2292
rect 24581 2255 24639 2261
rect 25130 2252 25136 2264
rect 25188 2252 25194 2304
rect 26206 2292 26234 2536
rect 27338 2524 27344 2576
rect 27396 2564 27402 2576
rect 28399 2567 28457 2573
rect 28399 2564 28411 2567
rect 27396 2536 28411 2564
rect 27396 2524 27402 2536
rect 28399 2533 28411 2536
rect 28445 2533 28457 2567
rect 28399 2527 28457 2533
rect 28534 2524 28540 2576
rect 28592 2564 28598 2576
rect 29779 2567 29837 2573
rect 29779 2564 29791 2567
rect 28592 2536 29791 2564
rect 28592 2524 28598 2536
rect 29779 2533 29791 2536
rect 29825 2533 29837 2567
rect 29779 2527 29837 2533
rect 32674 2524 32680 2576
rect 32732 2564 32738 2576
rect 34701 2567 34759 2573
rect 34701 2564 34713 2567
rect 32732 2536 34713 2564
rect 32732 2524 32738 2536
rect 34701 2533 34713 2536
rect 34747 2533 34759 2567
rect 34701 2527 34759 2533
rect 35066 2524 35072 2576
rect 35124 2564 35130 2576
rect 36173 2567 36231 2573
rect 36173 2564 36185 2567
rect 35124 2536 36185 2564
rect 35124 2524 35130 2536
rect 36173 2533 36185 2536
rect 36219 2533 36231 2567
rect 36173 2527 36231 2533
rect 37090 2524 37096 2576
rect 37148 2564 37154 2576
rect 38933 2567 38991 2573
rect 38933 2564 38945 2567
rect 37148 2536 38945 2564
rect 37148 2524 37154 2536
rect 38933 2533 38945 2536
rect 38979 2533 38991 2567
rect 38933 2527 38991 2533
rect 27522 2456 27528 2508
rect 27580 2496 27586 2508
rect 30837 2499 30895 2505
rect 30837 2496 30849 2499
rect 27580 2468 30849 2496
rect 27580 2456 27586 2468
rect 30837 2465 30849 2468
rect 30883 2465 30895 2499
rect 30837 2459 30895 2465
rect 32214 2456 32220 2508
rect 32272 2496 32278 2508
rect 33318 2496 33324 2508
rect 32272 2468 33324 2496
rect 32272 2456 32278 2468
rect 33318 2456 33324 2468
rect 33376 2496 33382 2508
rect 33376 2468 33456 2496
rect 33376 2456 33382 2468
rect 28169 2431 28227 2437
rect 28169 2397 28181 2431
rect 28215 2428 28227 2431
rect 28350 2428 28356 2440
rect 28215 2400 28356 2428
rect 28215 2397 28227 2400
rect 28169 2391 28227 2397
rect 28350 2388 28356 2400
rect 28408 2388 28414 2440
rect 29362 2388 29368 2440
rect 29420 2428 29426 2440
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29420 2400 29561 2428
rect 29420 2388 29426 2400
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 33428 2437 33456 2468
rect 34974 2456 34980 2508
rect 35032 2496 35038 2508
rect 43533 2499 43591 2505
rect 43533 2496 43545 2499
rect 35032 2468 43545 2496
rect 35032 2456 35038 2468
rect 43533 2465 43545 2468
rect 43579 2465 43591 2499
rect 43533 2459 43591 2465
rect 33229 2431 33287 2437
rect 33229 2428 33241 2431
rect 30432 2400 33241 2428
rect 30432 2388 30438 2400
rect 33229 2397 33241 2400
rect 33275 2397 33287 2431
rect 33229 2391 33287 2397
rect 33413 2431 33471 2437
rect 33413 2397 33425 2431
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 34054 2388 34060 2440
rect 34112 2428 34118 2440
rect 34112 2400 35020 2428
rect 34112 2388 34118 2400
rect 26510 2320 26516 2372
rect 26568 2360 26574 2372
rect 27246 2360 27252 2372
rect 26568 2332 27252 2360
rect 26568 2320 26574 2332
rect 27246 2320 27252 2332
rect 27304 2360 27310 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 27304 2332 27445 2360
rect 27304 2320 27310 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 27617 2363 27675 2369
rect 27617 2329 27629 2363
rect 27663 2360 27675 2363
rect 29914 2360 29920 2372
rect 27663 2332 29920 2360
rect 27663 2329 27675 2332
rect 27617 2323 27675 2329
rect 29914 2320 29920 2332
rect 29972 2320 29978 2372
rect 30282 2320 30288 2372
rect 30340 2360 30346 2372
rect 30742 2360 30748 2372
rect 30340 2332 30748 2360
rect 30340 2320 30346 2332
rect 30742 2320 30748 2332
rect 30800 2360 30806 2372
rect 31021 2363 31079 2369
rect 31021 2360 31033 2363
rect 30800 2332 31033 2360
rect 30800 2320 30806 2332
rect 31021 2329 31033 2332
rect 31067 2329 31079 2363
rect 31021 2323 31079 2329
rect 31294 2320 31300 2372
rect 31352 2360 31358 2372
rect 32677 2363 32735 2369
rect 32677 2360 32689 2363
rect 31352 2332 32689 2360
rect 31352 2320 31358 2332
rect 32677 2329 32689 2332
rect 32723 2329 32735 2363
rect 32677 2323 32735 2329
rect 28258 2292 28264 2304
rect 26206 2264 28264 2292
rect 28258 2252 28264 2264
rect 28316 2252 28322 2304
rect 32692 2292 32720 2323
rect 33134 2320 33140 2372
rect 33192 2360 33198 2372
rect 34606 2360 34612 2372
rect 33192 2332 34612 2360
rect 33192 2320 33198 2332
rect 34606 2320 34612 2332
rect 34664 2360 34670 2372
rect 34885 2363 34943 2369
rect 34885 2360 34897 2363
rect 34664 2332 34897 2360
rect 34664 2320 34670 2332
rect 34885 2329 34897 2332
rect 34931 2329 34943 2363
rect 34992 2360 35020 2400
rect 35066 2388 35072 2440
rect 35124 2428 35130 2440
rect 36078 2428 36084 2440
rect 35124 2400 36084 2428
rect 35124 2388 35130 2400
rect 36078 2388 36084 2400
rect 36136 2428 36142 2440
rect 36357 2431 36415 2437
rect 36357 2428 36369 2431
rect 36136 2400 36369 2428
rect 36136 2388 36142 2400
rect 36357 2397 36369 2400
rect 36403 2397 36415 2431
rect 36357 2391 36415 2397
rect 39758 2388 39764 2440
rect 39816 2428 39822 2440
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 39816 2400 39865 2428
rect 39816 2388 39822 2400
rect 39853 2397 39865 2400
rect 39899 2397 39911 2431
rect 39853 2391 39911 2397
rect 42794 2388 42800 2440
rect 42852 2428 42858 2440
rect 42981 2431 43039 2437
rect 42981 2428 42993 2431
rect 42852 2400 42993 2428
rect 42852 2388 42858 2400
rect 42981 2397 42993 2400
rect 43027 2397 43039 2431
rect 42981 2391 43039 2397
rect 35434 2360 35440 2372
rect 34992 2332 35440 2360
rect 34885 2323 34943 2329
rect 35434 2320 35440 2332
rect 35492 2360 35498 2372
rect 35621 2363 35679 2369
rect 35621 2360 35633 2363
rect 35492 2332 35633 2360
rect 35492 2320 35498 2332
rect 35621 2329 35633 2332
rect 35667 2329 35679 2363
rect 35621 2323 35679 2329
rect 37461 2363 37519 2369
rect 37461 2329 37473 2363
rect 37507 2360 37519 2363
rect 37826 2360 37832 2372
rect 37507 2332 37832 2360
rect 37507 2329 37519 2332
rect 37461 2323 37519 2329
rect 37826 2320 37832 2332
rect 37884 2360 37890 2372
rect 38105 2363 38163 2369
rect 38105 2360 38117 2363
rect 37884 2332 38117 2360
rect 37884 2320 37890 2332
rect 38105 2329 38117 2332
rect 38151 2329 38163 2363
rect 38105 2323 38163 2329
rect 38838 2320 38844 2372
rect 38896 2360 38902 2372
rect 39117 2363 39175 2369
rect 39117 2360 39129 2363
rect 38896 2332 39129 2360
rect 38896 2320 38902 2332
rect 39117 2329 39129 2332
rect 39163 2329 39175 2363
rect 39117 2323 39175 2329
rect 40678 2320 40684 2372
rect 40736 2360 40742 2372
rect 40957 2363 41015 2369
rect 40957 2360 40969 2363
rect 40736 2332 40969 2360
rect 40736 2320 40742 2332
rect 40957 2329 40969 2332
rect 41003 2329 41015 2363
rect 40957 2323 41015 2329
rect 41046 2320 41052 2372
rect 41104 2360 41110 2372
rect 41506 2360 41512 2372
rect 41104 2332 41512 2360
rect 41104 2320 41110 2332
rect 41506 2320 41512 2332
rect 41564 2360 41570 2372
rect 41693 2363 41751 2369
rect 41693 2360 41705 2363
rect 41564 2332 41705 2360
rect 41564 2320 41570 2332
rect 41693 2329 41705 2332
rect 41739 2329 41751 2363
rect 41693 2323 41751 2329
rect 42610 2320 42616 2372
rect 42668 2360 42674 2372
rect 43438 2360 43444 2372
rect 42668 2332 43444 2360
rect 42668 2320 42674 2332
rect 43438 2320 43444 2332
rect 43496 2360 43502 2372
rect 43717 2363 43775 2369
rect 43717 2360 43729 2363
rect 43496 2332 43729 2360
rect 43496 2320 43502 2332
rect 43717 2329 43729 2332
rect 43763 2329 43775 2363
rect 43717 2323 43775 2329
rect 33965 2295 34023 2301
rect 33965 2292 33977 2295
rect 32692 2264 33977 2292
rect 33965 2261 33977 2264
rect 34011 2261 34023 2295
rect 35526 2292 35532 2304
rect 35487 2264 35532 2292
rect 33965 2255 34023 2261
rect 35526 2252 35532 2264
rect 35584 2252 35590 2304
rect 40034 2292 40040 2304
rect 39995 2264 40040 2292
rect 40034 2252 40040 2264
rect 40092 2252 40098 2304
rect 40126 2252 40132 2304
rect 40184 2292 40190 2304
rect 40865 2295 40923 2301
rect 40865 2292 40877 2295
rect 40184 2264 40877 2292
rect 40184 2252 40190 2264
rect 40865 2261 40877 2264
rect 40911 2261 40923 2295
rect 41598 2292 41604 2304
rect 41559 2264 41604 2292
rect 40865 2255 40923 2261
rect 41598 2252 41604 2264
rect 41656 2252 41662 2304
rect 42886 2292 42892 2304
rect 42847 2264 42892 2292
rect 42886 2252 42892 2264
rect 42944 2252 42950 2304
rect 1104 2202 44896 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 44896 2202
rect 1104 2128 44896 2150
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 17310 2088 17316 2100
rect 7708 2060 17316 2088
rect 7708 2048 7714 2060
rect 17310 2048 17316 2060
rect 17368 2048 17374 2100
rect 20714 2048 20720 2100
rect 20772 2088 20778 2100
rect 41598 2088 41604 2100
rect 20772 2060 41604 2088
rect 20772 2048 20778 2060
rect 41598 2048 41604 2060
rect 41656 2048 41662 2100
rect 5534 1980 5540 2032
rect 5592 2020 5598 2032
rect 25682 2020 25688 2032
rect 5592 1992 25688 2020
rect 5592 1980 5598 1992
rect 25682 1980 25688 1992
rect 25740 1980 25746 2032
rect 31110 1980 31116 2032
rect 31168 2020 31174 2032
rect 34974 2020 34980 2032
rect 31168 1992 34980 2020
rect 31168 1980 31174 1992
rect 34974 1980 34980 1992
rect 35032 1980 35038 2032
rect 5718 1912 5724 1964
rect 5776 1952 5782 1964
rect 22922 1952 22928 1964
rect 5776 1924 22928 1952
rect 5776 1912 5782 1924
rect 22922 1912 22928 1924
rect 22980 1912 22986 1964
rect 27062 1912 27068 1964
rect 27120 1952 27126 1964
rect 40034 1952 40040 1964
rect 27120 1924 40040 1952
rect 27120 1912 27126 1924
rect 40034 1912 40040 1924
rect 40092 1912 40098 1964
rect 6362 1844 6368 1896
rect 6420 1884 6426 1896
rect 6822 1884 6828 1896
rect 6420 1856 6828 1884
rect 6420 1844 6426 1856
rect 6822 1844 6828 1856
rect 6880 1884 6886 1896
rect 25130 1884 25136 1896
rect 6880 1856 25136 1884
rect 6880 1844 6886 1856
rect 25130 1844 25136 1856
rect 25188 1844 25194 1896
rect 2866 1776 2872 1828
rect 2924 1816 2930 1828
rect 11606 1816 11612 1828
rect 2924 1788 11612 1816
rect 2924 1776 2930 1788
rect 11606 1776 11612 1788
rect 11664 1776 11670 1828
rect 13814 1776 13820 1828
rect 13872 1816 13878 1828
rect 24486 1816 24492 1828
rect 13872 1788 24492 1816
rect 13872 1776 13878 1788
rect 24486 1776 24492 1788
rect 24544 1776 24550 1828
rect 8110 1708 8116 1760
rect 8168 1748 8174 1760
rect 11974 1748 11980 1760
rect 8168 1720 11980 1748
rect 8168 1708 8174 1720
rect 11974 1708 11980 1720
rect 12032 1708 12038 1760
rect 18414 1708 18420 1760
rect 18472 1748 18478 1760
rect 35526 1748 35532 1760
rect 18472 1720 35532 1748
rect 18472 1708 18478 1720
rect 35526 1708 35532 1720
rect 35584 1708 35590 1760
rect 8018 1640 8024 1692
rect 8076 1680 8082 1692
rect 23934 1680 23940 1692
rect 8076 1652 23940 1680
rect 8076 1640 8082 1652
rect 23934 1640 23940 1652
rect 23992 1640 23998 1692
rect 7006 1572 7012 1624
rect 7064 1612 7070 1624
rect 7926 1612 7932 1624
rect 7064 1584 7932 1612
rect 7064 1572 7070 1584
rect 7926 1572 7932 1584
rect 7984 1612 7990 1624
rect 22002 1612 22008 1624
rect 7984 1584 22008 1612
rect 7984 1572 7990 1584
rect 22002 1572 22008 1584
rect 22060 1572 22066 1624
rect 17862 1504 17868 1556
rect 17920 1544 17926 1556
rect 20254 1544 20260 1556
rect 17920 1516 20260 1544
rect 17920 1504 17926 1516
rect 20254 1504 20260 1516
rect 20312 1504 20318 1556
rect 11790 1368 11796 1420
rect 11848 1408 11854 1420
rect 20438 1408 20444 1420
rect 11848 1380 20444 1408
rect 11848 1368 11854 1380
rect 20438 1368 20444 1380
rect 20496 1368 20502 1420
rect 14 1300 20 1352
rect 72 1340 78 1352
rect 934 1340 940 1352
rect 72 1312 940 1340
rect 72 1300 78 1312
rect 934 1300 940 1312
rect 992 1300 998 1352
rect 15378 1300 15384 1352
rect 15436 1340 15442 1352
rect 27522 1340 27528 1352
rect 15436 1312 27528 1340
rect 15436 1300 15442 1312
rect 27522 1300 27528 1312
rect 27580 1300 27586 1352
rect 17310 1232 17316 1284
rect 17368 1272 17374 1284
rect 20162 1272 20168 1284
rect 17368 1244 20168 1272
rect 17368 1232 17374 1244
rect 20162 1232 20168 1244
rect 20220 1232 20226 1284
rect 20438 1232 20444 1284
rect 20496 1272 20502 1284
rect 22186 1272 22192 1284
rect 20496 1244 22192 1272
rect 20496 1232 20502 1244
rect 22186 1232 22192 1244
rect 22244 1232 22250 1284
rect 6914 1164 6920 1216
rect 6972 1204 6978 1216
rect 24118 1204 24124 1216
rect 6972 1176 24124 1204
rect 6972 1164 6978 1176
rect 24118 1164 24124 1176
rect 24176 1164 24182 1216
rect 10778 1096 10784 1148
rect 10836 1136 10842 1148
rect 11238 1136 11244 1148
rect 10836 1108 11244 1136
rect 10836 1096 10842 1108
rect 11238 1096 11244 1108
rect 11296 1136 11302 1148
rect 17954 1136 17960 1148
rect 11296 1108 17960 1136
rect 11296 1096 11302 1108
rect 17954 1096 17960 1108
rect 18012 1096 18018 1148
rect 18138 1096 18144 1148
rect 18196 1136 18202 1148
rect 25406 1136 25412 1148
rect 18196 1108 25412 1136
rect 18196 1096 18202 1108
rect 25406 1096 25412 1108
rect 25464 1096 25470 1148
rect 7282 1028 7288 1080
rect 7340 1068 7346 1080
rect 8846 1068 8852 1080
rect 7340 1040 8852 1068
rect 7340 1028 7346 1040
rect 8846 1028 8852 1040
rect 8904 1068 8910 1080
rect 22278 1068 22284 1080
rect 8904 1040 22284 1068
rect 8904 1028 8910 1040
rect 22278 1028 22284 1040
rect 22336 1028 22342 1080
rect 2774 960 2780 1012
rect 2832 1000 2838 1012
rect 22554 1000 22560 1012
rect 2832 972 22560 1000
rect 2832 960 2838 972
rect 22554 960 22560 972
rect 22612 960 22618 1012
rect 7558 892 7564 944
rect 7616 932 7622 944
rect 7616 904 16574 932
rect 7616 892 7622 904
rect 5534 824 5540 876
rect 5592 864 5598 876
rect 16298 864 16304 876
rect 5592 836 16304 864
rect 5592 824 5598 836
rect 16298 824 16304 836
rect 16356 824 16362 876
rect 16546 864 16574 904
rect 17954 892 17960 944
rect 18012 932 18018 944
rect 23566 932 23572 944
rect 18012 904 23572 932
rect 18012 892 18018 904
rect 23566 892 23572 904
rect 23624 892 23630 944
rect 24762 864 24768 876
rect 16546 836 24768 864
rect 24762 824 24768 836
rect 24820 824 24826 876
rect 3786 756 3792 808
rect 3844 796 3850 808
rect 15102 796 15108 808
rect 3844 768 15108 796
rect 3844 756 3850 768
rect 15102 756 15108 768
rect 15160 756 15166 808
rect 4706 688 4712 740
rect 4764 728 4770 740
rect 16850 728 16856 740
rect 4764 700 16856 728
rect 4764 688 4770 700
rect 16850 688 16856 700
rect 16908 688 16914 740
rect 9398 348 9404 400
rect 9456 388 9462 400
rect 17862 388 17868 400
rect 9456 360 17868 388
rect 9456 348 9462 360
rect 17862 348 17868 360
rect 17920 348 17926 400
rect 13354 280 13360 332
rect 13412 320 13418 332
rect 23198 320 23204 332
rect 13412 292 23204 320
rect 13412 280 13418 292
rect 23198 280 23204 292
rect 23256 280 23262 332
rect 16206 212 16212 264
rect 16264 252 16270 264
rect 26326 252 26332 264
rect 16264 224 26332 252
rect 16264 212 16270 224
rect 26326 212 26332 224
rect 26384 212 26390 264
rect 11606 144 11612 196
rect 11664 184 11670 196
rect 12250 184 12256 196
rect 11664 156 12256 184
rect 11664 144 11670 156
rect 12250 144 12256 156
rect 12308 184 12314 196
rect 25498 184 25504 196
rect 12308 156 25504 184
rect 12308 144 12314 156
rect 25498 144 25504 156
rect 25556 144 25562 196
rect 14366 76 14372 128
rect 14424 116 14430 128
rect 26602 116 26608 128
rect 14424 88 26608 116
rect 14424 76 14430 88
rect 26602 76 26608 88
rect 26660 76 26666 128
rect 10686 8 10692 60
rect 10744 48 10750 60
rect 25314 48 25320 60
rect 10744 20 25320 48
rect 10744 8 10750 20
rect 25314 8 25320 20
rect 25372 8 25378 60
<< via1 >>
rect 21824 38020 21876 38072
rect 30012 38020 30064 38072
rect 12716 37952 12768 38004
rect 24952 37952 25004 38004
rect 9496 37884 9548 37936
rect 20260 37884 20312 37936
rect 20904 37884 20956 37936
rect 28172 37884 28224 37936
rect 2780 37816 2832 37868
rect 11152 37816 11204 37868
rect 18052 37816 18104 37868
rect 27436 37816 27488 37868
rect 27712 37816 27764 37868
rect 35808 37816 35860 37868
rect 3056 37748 3108 37800
rect 10324 37748 10376 37800
rect 10416 37748 10468 37800
rect 23848 37748 23900 37800
rect 29828 37748 29880 37800
rect 37832 37748 37884 37800
rect 3976 37680 4028 37732
rect 12440 37680 12492 37732
rect 17776 37680 17828 37732
rect 22560 37680 22612 37732
rect 25320 37680 25372 37732
rect 33324 37680 33376 37732
rect 7656 37612 7708 37664
rect 21456 37612 21508 37664
rect 24308 37612 24360 37664
rect 34704 37612 34756 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2780 37408 2832 37460
rect 3056 37451 3108 37460
rect 3056 37417 3065 37451
rect 3065 37417 3099 37451
rect 3099 37417 3108 37451
rect 3056 37408 3108 37417
rect 3516 37408 3568 37460
rect 5172 37408 5224 37460
rect 7656 37451 7708 37460
rect 7656 37417 7665 37451
rect 7665 37417 7699 37451
rect 7699 37417 7708 37451
rect 7656 37408 7708 37417
rect 9496 37451 9548 37460
rect 9496 37417 9505 37451
rect 9505 37417 9539 37451
rect 9539 37417 9548 37451
rect 9496 37408 9548 37417
rect 10416 37408 10468 37460
rect 4712 37340 4764 37392
rect 5356 37383 5408 37392
rect 5356 37349 5365 37383
rect 5365 37349 5399 37383
rect 5399 37349 5408 37383
rect 5356 37340 5408 37349
rect 8116 37340 8168 37392
rect 12716 37340 12768 37392
rect 21088 37383 21140 37392
rect 21088 37349 21097 37383
rect 21097 37349 21131 37383
rect 21131 37349 21140 37383
rect 21088 37340 21140 37349
rect 27436 37451 27488 37460
rect 22468 37340 22520 37392
rect 22560 37340 22612 37392
rect 27436 37417 27445 37451
rect 27445 37417 27479 37451
rect 27479 37417 27488 37451
rect 27436 37408 27488 37417
rect 28172 37451 28224 37460
rect 28172 37417 28181 37451
rect 28181 37417 28215 37451
rect 28215 37417 28224 37451
rect 28172 37408 28224 37417
rect 30012 37451 30064 37460
rect 30012 37417 30021 37451
rect 30021 37417 30055 37451
rect 30055 37417 30064 37451
rect 30012 37408 30064 37417
rect 33324 37451 33376 37460
rect 33324 37417 33333 37451
rect 33333 37417 33367 37451
rect 33367 37417 33376 37451
rect 33324 37408 33376 37417
rect 34704 37408 34756 37460
rect 37832 37451 37884 37460
rect 37832 37417 37841 37451
rect 37841 37417 37875 37451
rect 37875 37417 37884 37451
rect 37832 37408 37884 37417
rect 40408 37451 40460 37460
rect 40408 37417 40417 37451
rect 40417 37417 40451 37451
rect 40451 37417 40460 37451
rect 40408 37408 40460 37417
rect 41236 37451 41288 37460
rect 41236 37417 41245 37451
rect 41245 37417 41279 37451
rect 41279 37417 41288 37451
rect 41236 37408 41288 37417
rect 29736 37340 29788 37392
rect 3700 37272 3752 37324
rect 5080 37272 5132 37324
rect 204 37204 256 37256
rect 1492 37204 1544 37256
rect 2228 37247 2280 37256
rect 2228 37213 2237 37247
rect 2237 37213 2271 37247
rect 2271 37213 2280 37247
rect 2228 37204 2280 37213
rect 2780 37204 2832 37256
rect 3792 37204 3844 37256
rect 4804 37204 4856 37256
rect 4988 37204 5040 37256
rect 6184 37204 6236 37256
rect 12256 37272 12308 37324
rect 7380 37204 7432 37256
rect 8668 37204 8720 37256
rect 9588 37204 9640 37256
rect 9864 37204 9916 37256
rect 11060 37204 11112 37256
rect 13452 37272 13504 37324
rect 18328 37272 18380 37324
rect 19064 37272 19116 37324
rect 20076 37272 20128 37324
rect 24768 37315 24820 37324
rect 24768 37281 24777 37315
rect 24777 37281 24811 37315
rect 24811 37281 24820 37315
rect 24768 37272 24820 37281
rect 26884 37272 26936 37324
rect 35808 37383 35860 37392
rect 35808 37349 35817 37383
rect 35817 37349 35851 37383
rect 35851 37349 35860 37383
rect 35808 37340 35860 37349
rect 13360 37247 13412 37256
rect 13360 37213 13369 37247
rect 13369 37213 13403 37247
rect 13403 37213 13412 37247
rect 13360 37204 13412 37213
rect 15384 37247 15436 37256
rect 2412 37136 2464 37188
rect 15384 37213 15393 37247
rect 15393 37213 15427 37247
rect 15427 37213 15436 37247
rect 15384 37204 15436 37213
rect 15936 37204 15988 37256
rect 16672 37247 16724 37256
rect 16672 37213 16681 37247
rect 16681 37213 16715 37247
rect 16715 37213 16724 37247
rect 16672 37204 16724 37213
rect 16120 37136 16172 37188
rect 16580 37136 16632 37188
rect 17040 37204 17092 37256
rect 18604 37136 18656 37188
rect 20720 37204 20772 37256
rect 23204 37204 23256 37256
rect 23388 37204 23440 37256
rect 24400 37204 24452 37256
rect 25596 37204 25648 37256
rect 26792 37204 26844 37256
rect 27528 37247 27580 37256
rect 27528 37213 27537 37247
rect 27537 37213 27571 37247
rect 27571 37213 27580 37247
rect 27528 37204 27580 37213
rect 27988 37204 28040 37256
rect 29184 37204 29236 37256
rect 30380 37204 30432 37256
rect 31760 37204 31812 37256
rect 32864 37204 32916 37256
rect 33140 37204 33192 37256
rect 34060 37204 34112 37256
rect 35348 37204 35400 37256
rect 35716 37204 35768 37256
rect 37648 37204 37700 37256
rect 38384 37204 38436 37256
rect 38568 37204 38620 37256
rect 38936 37204 38988 37256
rect 40132 37204 40184 37256
rect 42340 37204 42392 37256
rect 43076 37204 43128 37256
rect 43444 37204 43496 37256
rect 22100 37136 22152 37188
rect 40224 37136 40276 37188
rect 41512 37179 41564 37188
rect 41512 37145 41521 37179
rect 41521 37145 41555 37179
rect 41555 37145 41564 37179
rect 41512 37136 41564 37145
rect 2596 37068 2648 37120
rect 12624 37068 12676 37120
rect 15200 37068 15252 37120
rect 16304 37068 16356 37120
rect 30748 37111 30800 37120
rect 30748 37077 30757 37111
rect 30757 37077 30791 37111
rect 30791 37077 30800 37111
rect 30748 37068 30800 37077
rect 38844 37111 38896 37120
rect 38844 37077 38853 37111
rect 38853 37077 38887 37111
rect 38887 37077 38896 37111
rect 38844 37068 38896 37077
rect 41696 37068 41748 37120
rect 42892 37068 42944 37120
rect 44180 37068 44232 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 572 36864 624 36916
rect 1768 36864 1820 36916
rect 2964 36864 3016 36916
rect 4160 36864 4212 36916
rect 4804 36864 4856 36916
rect 5540 36864 5592 36916
rect 6644 36864 6696 36916
rect 7840 36864 7892 36916
rect 9036 36864 9088 36916
rect 9404 36864 9456 36916
rect 10692 36864 10744 36916
rect 11428 36864 11480 36916
rect 13084 36864 13136 36916
rect 13912 36864 13964 36916
rect 16672 36907 16724 36916
rect 16672 36873 16681 36907
rect 16681 36873 16715 36907
rect 16715 36873 16724 36907
rect 16672 36864 16724 36873
rect 18696 36864 18748 36916
rect 20352 36864 20404 36916
rect 21180 36864 21232 36916
rect 22376 36864 22428 36916
rect 23572 36864 23624 36916
rect 24860 36864 24912 36916
rect 25964 36864 26016 36916
rect 27160 36864 27212 36916
rect 27528 36864 27580 36916
rect 28448 36864 28500 36916
rect 29644 36864 29696 36916
rect 30380 36864 30432 36916
rect 30840 36864 30892 36916
rect 32036 36864 32088 36916
rect 32404 36864 32456 36916
rect 33232 36864 33284 36916
rect 34520 36864 34572 36916
rect 35624 36864 35676 36916
rect 36084 36864 36136 36916
rect 37280 36864 37332 36916
rect 38384 36864 38436 36916
rect 39304 36864 39356 36916
rect 40500 36864 40552 36916
rect 42156 36864 42208 36916
rect 43352 36907 43404 36916
rect 43352 36873 43361 36907
rect 43361 36873 43395 36907
rect 43395 36873 43404 36907
rect 43352 36864 43404 36873
rect 45376 36864 45428 36916
rect 1308 36796 1360 36848
rect 3884 36728 3936 36780
rect 4712 36728 4764 36780
rect 6460 36728 6512 36780
rect 2504 36660 2556 36712
rect 8668 36728 8720 36780
rect 9496 36728 9548 36780
rect 10968 36771 11020 36780
rect 10968 36737 10977 36771
rect 10977 36737 11011 36771
rect 11011 36737 11020 36771
rect 10968 36728 11020 36737
rect 11980 36728 12032 36780
rect 12624 36728 12676 36780
rect 13728 36728 13780 36780
rect 14464 36728 14516 36780
rect 15660 36728 15712 36780
rect 17132 36728 17184 36780
rect 18236 36728 18288 36780
rect 19432 36728 19484 36780
rect 20628 36728 20680 36780
rect 22652 36728 22704 36780
rect 23204 36728 23256 36780
rect 23664 36771 23716 36780
rect 23664 36737 23673 36771
rect 23673 36737 23707 36771
rect 23707 36737 23716 36771
rect 23664 36728 23716 36737
rect 25228 36728 25280 36780
rect 26056 36771 26108 36780
rect 26056 36737 26065 36771
rect 26065 36737 26099 36771
rect 26099 36737 26108 36771
rect 26056 36728 26108 36737
rect 27068 36728 27120 36780
rect 28540 36771 28592 36780
rect 28540 36737 28549 36771
rect 28549 36737 28583 36771
rect 28583 36737 28592 36771
rect 28540 36728 28592 36737
rect 29552 36728 29604 36780
rect 30380 36728 30432 36780
rect 31024 36728 31076 36780
rect 32128 36771 32180 36780
rect 32128 36737 32137 36771
rect 32137 36737 32171 36771
rect 32171 36737 32180 36771
rect 32128 36728 32180 36737
rect 32680 36728 32732 36780
rect 33508 36728 33560 36780
rect 34244 36728 34296 36780
rect 35992 36771 36044 36780
rect 35992 36737 36001 36771
rect 36001 36737 36035 36771
rect 36035 36737 36044 36771
rect 35992 36728 36044 36737
rect 36268 36728 36320 36780
rect 36544 36728 36596 36780
rect 37096 36728 37148 36780
rect 37832 36728 37884 36780
rect 39212 36728 39264 36780
rect 40592 36771 40644 36780
rect 40592 36737 40601 36771
rect 40601 36737 40635 36771
rect 40635 36737 40644 36771
rect 40592 36728 40644 36737
rect 41420 36728 41472 36780
rect 42432 36771 42484 36780
rect 42432 36737 42441 36771
rect 42441 36737 42475 36771
rect 42475 36737 42484 36771
rect 42432 36728 42484 36737
rect 43168 36771 43220 36780
rect 43168 36737 43177 36771
rect 43177 36737 43211 36771
rect 43211 36737 43220 36771
rect 43168 36728 43220 36737
rect 43536 36728 43588 36780
rect 10876 36660 10928 36712
rect 15200 36660 15252 36712
rect 17500 36703 17552 36712
rect 17500 36669 17509 36703
rect 17509 36669 17543 36703
rect 17543 36669 17552 36703
rect 17500 36660 17552 36669
rect 19892 36703 19944 36712
rect 19892 36669 19901 36703
rect 19901 36669 19935 36703
rect 19935 36669 19944 36703
rect 19892 36660 19944 36669
rect 10232 36592 10284 36644
rect 37280 36635 37332 36644
rect 37280 36601 37289 36635
rect 37289 36601 37323 36635
rect 37323 36601 37332 36635
rect 37280 36592 37332 36601
rect 10784 36524 10836 36576
rect 41604 36524 41656 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 940 36320 992 36372
rect 2136 36320 2188 36372
rect 3424 36320 3476 36372
rect 4620 36320 4672 36372
rect 5816 36320 5868 36372
rect 7012 36320 7064 36372
rect 7380 36320 7432 36372
rect 8300 36320 8352 36372
rect 9588 36320 9640 36372
rect 9864 36320 9916 36372
rect 11060 36320 11112 36372
rect 11888 36320 11940 36372
rect 13452 36363 13504 36372
rect 13452 36329 13461 36363
rect 13461 36329 13495 36363
rect 13495 36329 13504 36363
rect 13452 36320 13504 36329
rect 14280 36320 14332 36372
rect 15476 36320 15528 36372
rect 16764 36320 16816 36372
rect 17592 36320 17644 36372
rect 17960 36320 18012 36372
rect 19984 36320 20036 36372
rect 20720 36363 20772 36372
rect 20720 36329 20729 36363
rect 20729 36329 20763 36363
rect 20763 36329 20772 36363
rect 20720 36320 20772 36329
rect 21548 36320 21600 36372
rect 22744 36320 22796 36372
rect 23388 36320 23440 36372
rect 23940 36320 23992 36372
rect 25136 36320 25188 36372
rect 25596 36320 25648 36372
rect 26424 36320 26476 36372
rect 27620 36320 27672 36372
rect 28540 36363 28592 36372
rect 28540 36329 28549 36363
rect 28549 36329 28583 36363
rect 28583 36329 28592 36363
rect 28540 36320 28592 36329
rect 30472 36363 30524 36372
rect 30472 36329 30481 36363
rect 30481 36329 30515 36363
rect 30515 36329 30524 36363
rect 30472 36320 30524 36329
rect 31208 36320 31260 36372
rect 33140 36363 33192 36372
rect 33140 36329 33149 36363
rect 33149 36329 33183 36363
rect 33183 36329 33192 36363
rect 33140 36320 33192 36329
rect 33692 36320 33744 36372
rect 34796 36320 34848 36372
rect 35716 36363 35768 36372
rect 35716 36329 35725 36363
rect 35725 36329 35759 36363
rect 35759 36329 35768 36363
rect 35716 36320 35768 36329
rect 35992 36320 36044 36372
rect 37096 36363 37148 36372
rect 37096 36329 37105 36363
rect 37105 36329 37139 36363
rect 37139 36329 37148 36363
rect 37096 36320 37148 36329
rect 37372 36320 37424 36372
rect 40040 36363 40092 36372
rect 40040 36329 40049 36363
rect 40049 36329 40083 36363
rect 40083 36329 40092 36363
rect 40040 36320 40092 36329
rect 40868 36320 40920 36372
rect 41512 36320 41564 36372
rect 42340 36363 42392 36372
rect 42340 36329 42349 36363
rect 42349 36329 42383 36363
rect 42383 36329 42392 36363
rect 42340 36320 42392 36329
rect 43076 36363 43128 36372
rect 43076 36329 43085 36363
rect 43085 36329 43119 36363
rect 43119 36329 43128 36363
rect 43076 36320 43128 36329
rect 44548 36320 44600 36372
rect 4620 36184 4672 36236
rect 3148 36159 3200 36168
rect 3148 36125 3157 36159
rect 3157 36125 3191 36159
rect 3191 36125 3200 36159
rect 3148 36116 3200 36125
rect 4988 36159 5040 36168
rect 3240 36048 3292 36100
rect 4988 36125 4997 36159
rect 4997 36125 5031 36159
rect 5031 36125 5040 36159
rect 4988 36116 5040 36125
rect 6920 36116 6972 36168
rect 7380 36159 7432 36168
rect 7380 36125 7389 36159
rect 7389 36125 7423 36159
rect 7423 36125 7432 36159
rect 7380 36116 7432 36125
rect 10140 36116 10192 36168
rect 13176 36116 13228 36168
rect 14372 36159 14424 36168
rect 14372 36125 14381 36159
rect 14381 36125 14415 36159
rect 14415 36125 14424 36159
rect 14372 36116 14424 36125
rect 15476 36116 15528 36168
rect 16948 36116 17000 36168
rect 17592 36159 17644 36168
rect 17592 36125 17601 36159
rect 17601 36125 17635 36159
rect 17635 36125 17644 36159
rect 17592 36116 17644 36125
rect 18328 36159 18380 36168
rect 18328 36125 18337 36159
rect 18337 36125 18371 36159
rect 18371 36125 18380 36159
rect 18328 36116 18380 36125
rect 5540 36048 5592 36100
rect 20536 36116 20588 36168
rect 22192 36116 22244 36168
rect 23296 36116 23348 36168
rect 23388 36116 23440 36168
rect 25044 36116 25096 36168
rect 26516 36159 26568 36168
rect 26516 36125 26525 36159
rect 26525 36125 26559 36159
rect 26559 36125 26568 36159
rect 26516 36116 26568 36125
rect 27620 36116 27672 36168
rect 30104 36116 30156 36168
rect 31116 36116 31168 36168
rect 33600 36116 33652 36168
rect 34704 36116 34756 36168
rect 38016 36159 38068 36168
rect 38016 36125 38025 36159
rect 38025 36125 38059 36159
rect 38059 36125 38068 36159
rect 38016 36116 38068 36125
rect 38660 36116 38712 36168
rect 39856 36159 39908 36168
rect 39856 36125 39865 36159
rect 39865 36125 39899 36159
rect 39899 36125 39908 36159
rect 39856 36116 39908 36125
rect 40776 36116 40828 36168
rect 43720 36116 43772 36168
rect 20444 36048 20496 36100
rect 2964 36023 3016 36032
rect 2964 35989 2973 36023
rect 2973 35989 3007 36023
rect 3007 35989 3016 36023
rect 2964 35980 3016 35989
rect 4068 35980 4120 36032
rect 8024 35980 8076 36032
rect 10876 36023 10928 36032
rect 10876 35989 10885 36023
rect 10885 35989 10919 36023
rect 10919 35989 10928 36023
rect 10876 35980 10928 35989
rect 19340 36023 19392 36032
rect 19340 35989 19349 36023
rect 19349 35989 19383 36023
rect 19383 35989 19392 36023
rect 19340 35980 19392 35989
rect 29644 36023 29696 36032
rect 29644 35989 29653 36023
rect 29653 35989 29687 36023
rect 29687 35989 29696 36023
rect 29644 35980 29696 35989
rect 30288 35980 30340 36032
rect 32128 35980 32180 36032
rect 38936 36023 38988 36032
rect 38936 35989 38945 36023
rect 38945 35989 38979 36023
rect 38979 35989 38988 36023
rect 38936 35980 38988 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 2412 35776 2464 35828
rect 3148 35776 3200 35828
rect 4896 35819 4948 35828
rect 4896 35785 4905 35819
rect 4905 35785 4939 35819
rect 4939 35785 4948 35819
rect 4896 35776 4948 35785
rect 17132 35819 17184 35828
rect 17132 35785 17141 35819
rect 17141 35785 17175 35819
rect 17175 35785 17184 35819
rect 17132 35776 17184 35785
rect 19064 35819 19116 35828
rect 19064 35785 19073 35819
rect 19073 35785 19107 35819
rect 19107 35785 19116 35819
rect 19064 35776 19116 35785
rect 19432 35776 19484 35828
rect 22100 35819 22152 35828
rect 22100 35785 22109 35819
rect 22109 35785 22143 35819
rect 22143 35785 22152 35819
rect 22100 35776 22152 35785
rect 24400 35776 24452 35828
rect 28816 35776 28868 35828
rect 29644 35776 29696 35828
rect 38108 35776 38160 35828
rect 38844 35776 38896 35828
rect 40132 35819 40184 35828
rect 40132 35785 40141 35819
rect 40141 35785 40175 35819
rect 40175 35785 40184 35819
rect 40132 35776 40184 35785
rect 41420 35776 41472 35828
rect 45744 35776 45796 35828
rect 2044 35572 2096 35624
rect 2688 35708 2740 35760
rect 22652 35751 22704 35760
rect 22652 35717 22661 35751
rect 22661 35717 22695 35751
rect 22695 35717 22704 35751
rect 22652 35708 22704 35717
rect 28724 35708 28776 35760
rect 38476 35708 38528 35760
rect 38936 35708 38988 35760
rect 2780 35640 2832 35692
rect 33508 35683 33560 35692
rect 2964 35572 3016 35624
rect 6460 35547 6512 35556
rect 6460 35513 6469 35547
rect 6469 35513 6503 35547
rect 6503 35513 6512 35547
rect 6460 35504 6512 35513
rect 9404 35504 9456 35556
rect 10140 35547 10192 35556
rect 10140 35513 10149 35547
rect 10149 35513 10183 35547
rect 10183 35513 10192 35547
rect 10140 35504 10192 35513
rect 12256 35504 12308 35556
rect 25596 35504 25648 35556
rect 33508 35649 33517 35683
rect 33517 35649 33551 35683
rect 33551 35649 33560 35683
rect 33508 35640 33560 35649
rect 43628 35640 43680 35692
rect 26332 35572 26384 35624
rect 30104 35615 30156 35624
rect 30104 35581 30113 35615
rect 30113 35581 30147 35615
rect 30147 35581 30156 35615
rect 30104 35572 30156 35581
rect 27620 35547 27672 35556
rect 27620 35513 27629 35547
rect 27629 35513 27663 35547
rect 27663 35513 27672 35547
rect 27620 35504 27672 35513
rect 1584 35479 1636 35488
rect 1584 35445 1593 35479
rect 1593 35445 1627 35479
rect 1627 35445 1636 35479
rect 1584 35436 1636 35445
rect 2412 35436 2464 35488
rect 8668 35436 8720 35488
rect 9496 35479 9548 35488
rect 9496 35445 9505 35479
rect 9505 35445 9539 35479
rect 9539 35445 9548 35479
rect 9496 35436 9548 35445
rect 10968 35479 11020 35488
rect 10968 35445 10977 35479
rect 10977 35445 11011 35479
rect 11011 35445 11020 35479
rect 10968 35436 11020 35445
rect 11980 35479 12032 35488
rect 11980 35445 11989 35479
rect 11989 35445 12023 35479
rect 12023 35445 12032 35479
rect 11980 35436 12032 35445
rect 12624 35479 12676 35488
rect 12624 35445 12633 35479
rect 12633 35445 12667 35479
rect 12667 35445 12676 35479
rect 12624 35436 12676 35445
rect 13176 35479 13228 35488
rect 13176 35445 13185 35479
rect 13185 35445 13219 35479
rect 13219 35445 13228 35479
rect 13176 35436 13228 35445
rect 14464 35479 14516 35488
rect 14464 35445 14473 35479
rect 14473 35445 14507 35479
rect 14507 35445 14516 35479
rect 14464 35436 14516 35445
rect 23204 35479 23256 35488
rect 23204 35445 23213 35479
rect 23213 35445 23247 35479
rect 23247 35445 23256 35479
rect 23204 35436 23256 35445
rect 23664 35479 23716 35488
rect 23664 35445 23673 35479
rect 23673 35445 23707 35479
rect 23707 35445 23716 35479
rect 23664 35436 23716 35445
rect 25228 35479 25280 35488
rect 25228 35445 25237 35479
rect 25237 35445 25271 35479
rect 25271 35445 25280 35479
rect 25228 35436 25280 35445
rect 26056 35436 26108 35488
rect 27068 35479 27120 35488
rect 27068 35445 27077 35479
rect 27077 35445 27111 35479
rect 27111 35445 27120 35479
rect 27068 35436 27120 35445
rect 29552 35479 29604 35488
rect 29552 35445 29561 35479
rect 29561 35445 29595 35479
rect 29595 35445 29604 35479
rect 29552 35436 29604 35445
rect 31024 35479 31076 35488
rect 31024 35445 31033 35479
rect 31033 35445 31067 35479
rect 31067 35445 31076 35479
rect 31024 35436 31076 35445
rect 32680 35479 32732 35488
rect 32680 35445 32689 35479
rect 32689 35445 32723 35479
rect 32723 35445 32732 35479
rect 32680 35436 32732 35445
rect 34244 35436 34296 35488
rect 34704 35436 34756 35488
rect 36268 35479 36320 35488
rect 36268 35445 36277 35479
rect 36277 35445 36311 35479
rect 36311 35445 36320 35479
rect 36268 35436 36320 35445
rect 37832 35479 37884 35488
rect 37832 35445 37841 35479
rect 37841 35445 37875 35479
rect 37875 35445 37884 35479
rect 37832 35436 37884 35445
rect 38568 35479 38620 35488
rect 38568 35445 38577 35479
rect 38577 35445 38611 35479
rect 38611 35445 38620 35479
rect 38568 35436 38620 35445
rect 39212 35479 39264 35488
rect 39212 35445 39221 35479
rect 39221 35445 39255 35479
rect 39255 35445 39264 35479
rect 39212 35436 39264 35445
rect 40592 35479 40644 35488
rect 40592 35445 40601 35479
rect 40601 35445 40635 35479
rect 40635 35445 40644 35479
rect 40592 35436 40644 35445
rect 42432 35479 42484 35488
rect 42432 35445 42441 35479
rect 42441 35445 42475 35479
rect 42475 35445 42484 35479
rect 42432 35436 42484 35445
rect 43352 35479 43404 35488
rect 43352 35445 43361 35479
rect 43361 35445 43395 35479
rect 43395 35445 43404 35479
rect 43352 35436 43404 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1584 35275 1636 35284
rect 1584 35241 1593 35275
rect 1593 35241 1627 35275
rect 1627 35241 1636 35275
rect 1584 35232 1636 35241
rect 2044 35275 2096 35284
rect 2044 35241 2053 35275
rect 2053 35241 2087 35275
rect 2087 35241 2096 35275
rect 2044 35232 2096 35241
rect 2228 35232 2280 35284
rect 22376 35232 22428 35284
rect 26332 35232 26384 35284
rect 26516 35232 26568 35284
rect 38016 35232 38068 35284
rect 22192 35164 22244 35216
rect 26240 35164 26292 35216
rect 24216 35096 24268 35148
rect 32680 35096 32732 35148
rect 1400 35071 1452 35080
rect 1400 35037 1409 35071
rect 1409 35037 1443 35071
rect 1443 35037 1452 35071
rect 1400 35028 1452 35037
rect 2872 35028 2924 35080
rect 18420 35028 18472 35080
rect 26516 35028 26568 35080
rect 4620 34960 4672 35012
rect 6368 34960 6420 35012
rect 20168 34960 20220 35012
rect 26056 34960 26108 35012
rect 3884 34935 3936 34944
rect 3884 34901 3893 34935
rect 3893 34901 3927 34935
rect 3927 34901 3936 34935
rect 3884 34892 3936 34901
rect 5540 34892 5592 34944
rect 6736 34892 6788 34944
rect 23296 34935 23348 34944
rect 23296 34901 23305 34935
rect 23305 34901 23339 34935
rect 23339 34901 23348 34935
rect 23296 34892 23348 34901
rect 23388 34892 23440 34944
rect 25044 34935 25096 34944
rect 25044 34901 25053 34935
rect 25053 34901 25087 34935
rect 25087 34901 25096 34935
rect 25044 34892 25096 34901
rect 30380 34935 30432 34944
rect 30380 34901 30389 34935
rect 30389 34901 30423 34935
rect 30423 34901 30432 34935
rect 30380 34892 30432 34901
rect 31116 34935 31168 34944
rect 31116 34901 31125 34935
rect 31125 34901 31159 34935
rect 31159 34901 31168 34935
rect 31116 34892 31168 34901
rect 33600 34935 33652 34944
rect 33600 34901 33609 34935
rect 33609 34901 33643 34935
rect 33643 34901 33652 34935
rect 33600 34892 33652 34901
rect 34520 34892 34572 34944
rect 38016 34892 38068 34944
rect 38660 34935 38712 34944
rect 38660 34901 38669 34935
rect 38669 34901 38703 34935
rect 38703 34901 38712 34935
rect 38660 34892 38712 34901
rect 39856 34935 39908 34944
rect 39856 34901 39865 34935
rect 39865 34901 39899 34935
rect 39899 34901 39908 34935
rect 39856 34892 39908 34901
rect 40776 34935 40828 34944
rect 40776 34901 40785 34935
rect 40785 34901 40819 34935
rect 40819 34901 40828 34935
rect 40776 34892 40828 34901
rect 41328 34892 41380 34944
rect 43168 34892 43220 34944
rect 43536 34892 43588 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2780 34688 2832 34740
rect 25780 34688 25832 34740
rect 33600 34688 33652 34740
rect 20996 34620 21048 34672
rect 23664 34620 23716 34672
rect 1400 34595 1452 34604
rect 1400 34561 1409 34595
rect 1409 34561 1443 34595
rect 1443 34561 1452 34595
rect 1400 34552 1452 34561
rect 3240 34595 3292 34604
rect 3240 34561 3249 34595
rect 3249 34561 3283 34595
rect 3283 34561 3292 34595
rect 3240 34552 3292 34561
rect 5172 34552 5224 34604
rect 10968 34552 11020 34604
rect 12992 34552 13044 34604
rect 22836 34552 22888 34604
rect 25228 34552 25280 34604
rect 3516 34484 3568 34536
rect 6828 34484 6880 34536
rect 11980 34484 12032 34536
rect 13268 34484 13320 34536
rect 14464 34484 14516 34536
rect 15016 34484 15068 34536
rect 22744 34484 22796 34536
rect 23388 34484 23440 34536
rect 26240 34484 26292 34536
rect 27252 34484 27304 34536
rect 43720 34527 43772 34536
rect 43720 34493 43729 34527
rect 43729 34493 43763 34527
rect 43763 34493 43772 34527
rect 43720 34484 43772 34493
rect 1584 34391 1636 34400
rect 1584 34357 1593 34391
rect 1593 34357 1627 34391
rect 1627 34357 1636 34391
rect 1584 34348 1636 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 1492 34187 1544 34196
rect 1492 34153 1501 34187
rect 1501 34153 1535 34187
rect 1535 34153 1544 34187
rect 1492 34144 1544 34153
rect 2872 34144 2924 34196
rect 2504 33847 2556 33856
rect 2504 33813 2513 33847
rect 2513 33813 2547 33847
rect 2547 33813 2556 33847
rect 2504 33804 2556 33813
rect 23204 33804 23256 33856
rect 29460 33804 29512 33856
rect 43628 33804 43680 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1492 33464 1544 33516
rect 1400 33303 1452 33312
rect 1400 33269 1409 33303
rect 1409 33269 1443 33303
rect 1443 33269 1452 33303
rect 1400 33260 1452 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 21548 33056 21600 33108
rect 28540 33056 28592 33108
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 2596 32444 2648 32496
rect 20076 32444 20128 32496
rect 35348 32444 35400 32496
rect 43720 32444 43772 32496
rect 1492 32376 1544 32428
rect 32772 32376 32824 32428
rect 43076 32376 43128 32428
rect 1676 32172 1728 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1768 31968 1820 32020
rect 1584 31875 1636 31884
rect 1584 31841 1593 31875
rect 1593 31841 1627 31875
rect 1627 31841 1636 31875
rect 1584 31832 1636 31841
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 1676 31807 1728 31816
rect 1676 31773 1685 31807
rect 1685 31773 1719 31807
rect 1719 31773 1728 31807
rect 1676 31764 1728 31773
rect 1860 31671 1912 31680
rect 1860 31637 1869 31671
rect 1869 31637 1903 31671
rect 1903 31637 1912 31671
rect 1860 31628 1912 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1768 31424 1820 31476
rect 1400 31331 1452 31340
rect 1400 31297 1409 31331
rect 1409 31297 1443 31331
rect 1443 31297 1452 31331
rect 1400 31288 1452 31297
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 1400 30243 1452 30252
rect 1400 30209 1409 30243
rect 1409 30209 1443 30243
rect 1443 30209 1452 30243
rect 1400 30200 1452 30209
rect 29000 30200 29052 30252
rect 1584 30039 1636 30048
rect 1584 30005 1593 30039
rect 1593 30005 1627 30039
rect 1627 30005 1636 30039
rect 1584 29996 1636 30005
rect 44088 30039 44140 30048
rect 44088 30005 44097 30039
rect 44097 30005 44131 30039
rect 44131 30005 44140 30039
rect 44088 29996 44140 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 33140 29656 33192 29708
rect 41328 29656 41380 29708
rect 28080 29588 28132 29640
rect 41604 29588 41656 29640
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 3516 28976 3568 29028
rect 4896 28976 4948 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1492 28500 1544 28552
rect 1400 28407 1452 28416
rect 1400 28373 1409 28407
rect 1409 28373 1443 28407
rect 1443 28373 1452 28407
rect 1400 28364 1452 28373
rect 29276 28364 29328 28416
rect 39856 28364 39908 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 1400 28135 1452 28144
rect 1400 28101 1409 28135
rect 1409 28101 1443 28135
rect 1443 28101 1452 28135
rect 1400 28092 1452 28101
rect 1676 28067 1728 28076
rect 1676 28033 1685 28067
rect 1685 28033 1719 28067
rect 1719 28033 1728 28067
rect 1676 28024 1728 28033
rect 1584 27999 1636 28008
rect 1584 27965 1593 27999
rect 1593 27965 1627 27999
rect 1627 27965 1636 27999
rect 1584 27956 1636 27965
rect 10876 27888 10928 27940
rect 1584 27863 1636 27872
rect 1584 27829 1593 27863
rect 1593 27829 1627 27863
rect 1627 27829 1636 27863
rect 1584 27820 1636 27829
rect 2780 27820 2832 27872
rect 11060 27820 11112 27872
rect 31116 27820 31168 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 1676 27616 1728 27668
rect 7472 27616 7524 27668
rect 29368 27616 29420 27668
rect 1860 27548 1912 27600
rect 2688 27591 2740 27600
rect 2688 27557 2697 27591
rect 2697 27557 2731 27591
rect 2731 27557 2740 27591
rect 2688 27548 2740 27557
rect 2780 27523 2832 27532
rect 2780 27489 2789 27523
rect 2789 27489 2823 27523
rect 2823 27489 2832 27523
rect 2780 27480 2832 27489
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 2412 27455 2464 27464
rect 2412 27421 2421 27455
rect 2421 27421 2455 27455
rect 2455 27421 2464 27455
rect 2412 27412 2464 27421
rect 3056 27319 3108 27328
rect 3056 27285 3065 27319
rect 3065 27285 3099 27319
rect 3099 27285 3108 27319
rect 3056 27276 3108 27285
rect 8484 27276 8536 27328
rect 9036 27319 9088 27328
rect 9036 27285 9045 27319
rect 9045 27285 9079 27319
rect 9079 27285 9088 27319
rect 9036 27276 9088 27285
rect 9588 27319 9640 27328
rect 9588 27285 9597 27319
rect 9597 27285 9631 27319
rect 9631 27285 9640 27319
rect 9588 27276 9640 27285
rect 10968 27276 11020 27328
rect 26608 27276 26660 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 1400 27115 1452 27124
rect 1400 27081 1409 27115
rect 1409 27081 1443 27115
rect 1443 27081 1452 27115
rect 1400 27072 1452 27081
rect 8024 27115 8076 27124
rect 8024 27081 8033 27115
rect 8033 27081 8067 27115
rect 8067 27081 8076 27115
rect 8024 27072 8076 27081
rect 9588 27072 9640 27124
rect 9036 27004 9088 27056
rect 17408 27004 17460 27056
rect 4068 26936 4120 26988
rect 11336 26936 11388 26988
rect 10508 26868 10560 26920
rect 25228 26868 25280 26920
rect 6644 26800 6696 26852
rect 11520 26843 11572 26852
rect 11520 26809 11529 26843
rect 11529 26809 11563 26843
rect 11563 26809 11572 26843
rect 11520 26800 11572 26809
rect 11704 26800 11756 26852
rect 1860 26732 1912 26784
rect 2228 26732 2280 26784
rect 8576 26775 8628 26784
rect 8576 26741 8585 26775
rect 8585 26741 8619 26775
rect 8619 26741 8628 26775
rect 8576 26732 8628 26741
rect 10048 26732 10100 26784
rect 10232 26732 10284 26784
rect 10876 26775 10928 26784
rect 10876 26741 10885 26775
rect 10885 26741 10919 26775
rect 10919 26741 10928 26775
rect 10876 26732 10928 26741
rect 16304 26732 16356 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 1584 26571 1636 26580
rect 1584 26537 1593 26571
rect 1593 26537 1627 26571
rect 1627 26537 1636 26571
rect 1584 26528 1636 26537
rect 2412 26528 2464 26580
rect 6644 26528 6696 26580
rect 6828 26528 6880 26580
rect 10416 26571 10468 26580
rect 6092 26460 6144 26512
rect 9496 26503 9548 26512
rect 9496 26469 9505 26503
rect 9505 26469 9539 26503
rect 9539 26469 9548 26503
rect 9496 26460 9548 26469
rect 10416 26537 10425 26571
rect 10425 26537 10459 26571
rect 10459 26537 10468 26571
rect 10416 26528 10468 26537
rect 11520 26460 11572 26512
rect 16488 26528 16540 26580
rect 12624 26503 12676 26512
rect 12624 26469 12633 26503
rect 12633 26469 12667 26503
rect 12667 26469 12676 26503
rect 12624 26460 12676 26469
rect 13360 26460 13412 26512
rect 31576 26460 31628 26512
rect 30196 26392 30248 26444
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 2136 26324 2188 26376
rect 9588 26324 9640 26376
rect 12072 26324 12124 26376
rect 3792 26299 3844 26308
rect 3792 26265 3801 26299
rect 3801 26265 3835 26299
rect 3835 26265 3844 26299
rect 3792 26256 3844 26265
rect 8760 26256 8812 26308
rect 10508 26256 10560 26308
rect 10600 26256 10652 26308
rect 2504 26188 2556 26240
rect 8300 26231 8352 26240
rect 8300 26197 8309 26231
rect 8309 26197 8343 26231
rect 8343 26197 8352 26231
rect 8300 26188 8352 26197
rect 9864 26188 9916 26240
rect 19340 26324 19392 26376
rect 13084 26299 13136 26308
rect 13084 26265 13093 26299
rect 13093 26265 13127 26299
rect 13127 26265 13136 26299
rect 13084 26256 13136 26265
rect 16488 26256 16540 26308
rect 33232 26324 33284 26376
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 6920 26027 6972 26036
rect 6920 25993 6929 26027
rect 6929 25993 6963 26027
rect 6963 25993 6972 26027
rect 6920 25984 6972 25993
rect 10324 25984 10376 26036
rect 12072 26027 12124 26036
rect 12072 25993 12081 26027
rect 12081 25993 12115 26027
rect 12115 25993 12124 26027
rect 12072 25984 12124 25993
rect 7656 25848 7708 25900
rect 10048 25848 10100 25900
rect 1400 25780 1452 25832
rect 8576 25780 8628 25832
rect 10140 25780 10192 25832
rect 12072 25712 12124 25764
rect 25136 25712 25188 25764
rect 1492 25687 1544 25696
rect 1492 25653 1501 25687
rect 1501 25653 1535 25687
rect 1535 25653 1544 25687
rect 1492 25644 1544 25653
rect 2320 25644 2372 25696
rect 2872 25687 2924 25696
rect 2872 25653 2881 25687
rect 2881 25653 2915 25687
rect 2915 25653 2924 25687
rect 2872 25644 2924 25653
rect 2964 25644 3016 25696
rect 3240 25644 3292 25696
rect 3516 25644 3568 25696
rect 5724 25644 5776 25696
rect 7656 25687 7708 25696
rect 7656 25653 7665 25687
rect 7665 25653 7699 25687
rect 7699 25653 7708 25687
rect 7656 25644 7708 25653
rect 8392 25644 8444 25696
rect 9220 25644 9272 25696
rect 9772 25644 9824 25696
rect 11520 25687 11572 25696
rect 11520 25653 11529 25687
rect 11529 25653 11563 25687
rect 11563 25653 11572 25687
rect 11520 25644 11572 25653
rect 13084 25644 13136 25696
rect 14096 25687 14148 25696
rect 14096 25653 14105 25687
rect 14105 25653 14139 25687
rect 14139 25653 14148 25687
rect 14096 25644 14148 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 4988 25440 5040 25492
rect 5080 25440 5132 25492
rect 5448 25440 5500 25492
rect 756 25372 808 25424
rect 3148 25372 3200 25424
rect 3608 25372 3660 25424
rect 7564 25440 7616 25492
rect 9036 25440 9088 25492
rect 9588 25440 9640 25492
rect 10508 25440 10560 25492
rect 11152 25483 11204 25492
rect 11152 25449 11161 25483
rect 11161 25449 11195 25483
rect 11195 25449 11204 25483
rect 11152 25440 11204 25449
rect 11428 25440 11480 25492
rect 12532 25440 12584 25492
rect 11244 25372 11296 25424
rect 12624 25372 12676 25424
rect 18880 25372 18932 25424
rect 1216 25304 1268 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 1952 25236 2004 25288
rect 5724 25236 5776 25288
rect 5908 25236 5960 25288
rect 8300 25236 8352 25288
rect 12440 25304 12492 25356
rect 31760 25304 31812 25356
rect 11336 25236 11388 25288
rect 11888 25236 11940 25288
rect 14464 25236 14516 25288
rect 23848 25236 23900 25288
rect 8484 25168 8536 25220
rect 18880 25168 18932 25220
rect 23020 25168 23072 25220
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 3148 25100 3200 25152
rect 3884 25100 3936 25152
rect 6644 25143 6696 25152
rect 6644 25109 6653 25143
rect 6653 25109 6687 25143
rect 6687 25109 6696 25143
rect 6644 25100 6696 25109
rect 7196 25143 7248 25152
rect 7196 25109 7205 25143
rect 7205 25109 7239 25143
rect 7239 25109 7248 25143
rect 7196 25100 7248 25109
rect 7288 25100 7340 25152
rect 12348 25100 12400 25152
rect 16764 25100 16816 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 3148 24896 3200 24948
rect 9864 24896 9916 24948
rect 11060 24896 11112 24948
rect 15752 24896 15804 24948
rect 18696 24896 18748 24948
rect 18788 24896 18840 24948
rect 26332 24896 26384 24948
rect 10048 24828 10100 24880
rect 12348 24828 12400 24880
rect 17684 24828 17736 24880
rect 18052 24828 18104 24880
rect 33508 24828 33560 24880
rect 3148 24760 3200 24812
rect 3424 24760 3476 24812
rect 5264 24760 5316 24812
rect 2780 24692 2832 24744
rect 3056 24692 3108 24744
rect 8300 24760 8352 24812
rect 8576 24803 8628 24812
rect 8576 24769 8585 24803
rect 8585 24769 8619 24803
rect 8619 24769 8628 24803
rect 8576 24760 8628 24769
rect 9772 24803 9824 24812
rect 9772 24769 9781 24803
rect 9781 24769 9815 24803
rect 9815 24769 9824 24803
rect 9772 24760 9824 24769
rect 10600 24803 10652 24812
rect 10600 24769 10609 24803
rect 10609 24769 10643 24803
rect 10643 24769 10652 24803
rect 10600 24760 10652 24769
rect 14096 24760 14148 24812
rect 15844 24760 15896 24812
rect 22928 24760 22980 24812
rect 2044 24624 2096 24676
rect 4160 24667 4212 24676
rect 4160 24633 4169 24667
rect 4169 24633 4203 24667
rect 4203 24633 4212 24667
rect 4160 24624 4212 24633
rect 2412 24599 2464 24608
rect 2412 24565 2421 24599
rect 2421 24565 2455 24599
rect 2455 24565 2464 24599
rect 2412 24556 2464 24565
rect 4712 24599 4764 24608
rect 4712 24565 4721 24599
rect 4721 24565 4755 24599
rect 4755 24565 4764 24599
rect 4712 24556 4764 24565
rect 5080 24556 5132 24608
rect 8392 24692 8444 24744
rect 7472 24624 7524 24676
rect 16396 24692 16448 24744
rect 26976 24692 27028 24744
rect 11612 24624 11664 24676
rect 17316 24624 17368 24676
rect 5816 24599 5868 24608
rect 5816 24565 5825 24599
rect 5825 24565 5859 24599
rect 5859 24565 5868 24599
rect 5816 24556 5868 24565
rect 6276 24556 6328 24608
rect 7104 24599 7156 24608
rect 7104 24565 7113 24599
rect 7113 24565 7147 24599
rect 7147 24565 7156 24599
rect 7104 24556 7156 24565
rect 8116 24556 8168 24608
rect 8300 24556 8352 24608
rect 8944 24556 8996 24608
rect 9956 24599 10008 24608
rect 9956 24565 9965 24599
rect 9965 24565 9999 24599
rect 9999 24565 10008 24599
rect 9956 24556 10008 24565
rect 12164 24599 12216 24608
rect 12164 24565 12173 24599
rect 12173 24565 12207 24599
rect 12207 24565 12216 24599
rect 12164 24556 12216 24565
rect 12808 24556 12860 24608
rect 14372 24599 14424 24608
rect 14372 24565 14381 24599
rect 14381 24565 14415 24599
rect 14415 24565 14424 24599
rect 14372 24556 14424 24565
rect 15936 24599 15988 24608
rect 15936 24565 15945 24599
rect 15945 24565 15979 24599
rect 15979 24565 15988 24599
rect 15936 24556 15988 24565
rect 17040 24556 17092 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1768 24352 1820 24404
rect 2688 24352 2740 24404
rect 11520 24395 11572 24404
rect 11520 24361 11529 24395
rect 11529 24361 11563 24395
rect 11563 24361 11572 24395
rect 11520 24352 11572 24361
rect 12072 24352 12124 24404
rect 13176 24352 13228 24404
rect 15200 24352 15252 24404
rect 16304 24395 16356 24404
rect 16304 24361 16313 24395
rect 16313 24361 16347 24395
rect 16347 24361 16356 24395
rect 16304 24352 16356 24361
rect 17224 24352 17276 24404
rect 17408 24395 17460 24404
rect 17408 24361 17417 24395
rect 17417 24361 17451 24395
rect 17451 24361 17460 24395
rect 17408 24352 17460 24361
rect 17776 24352 17828 24404
rect 18788 24352 18840 24404
rect 19156 24352 19208 24404
rect 19984 24352 20036 24404
rect 22100 24395 22152 24404
rect 22100 24361 22109 24395
rect 22109 24361 22143 24395
rect 22143 24361 22152 24395
rect 22100 24352 22152 24361
rect 7748 24327 7800 24336
rect 7748 24293 7757 24327
rect 7757 24293 7791 24327
rect 7791 24293 7800 24327
rect 7748 24284 7800 24293
rect 9588 24284 9640 24336
rect 9864 24284 9916 24336
rect 13636 24284 13688 24336
rect 1584 24259 1636 24268
rect 1584 24225 1593 24259
rect 1593 24225 1627 24259
rect 1627 24225 1636 24259
rect 1584 24216 1636 24225
rect 9036 24259 9088 24268
rect 9036 24225 9045 24259
rect 9045 24225 9079 24259
rect 9079 24225 9088 24259
rect 9036 24216 9088 24225
rect 14188 24259 14240 24268
rect 1676 24191 1728 24200
rect 1676 24157 1685 24191
rect 1685 24157 1719 24191
rect 1719 24157 1728 24191
rect 1676 24148 1728 24157
rect 5724 24148 5776 24200
rect 9680 24148 9732 24200
rect 11336 24191 11388 24200
rect 11336 24157 11345 24191
rect 11345 24157 11379 24191
rect 11379 24157 11388 24191
rect 11336 24148 11388 24157
rect 1400 24123 1452 24132
rect 1400 24089 1409 24123
rect 1409 24089 1443 24123
rect 1443 24089 1452 24123
rect 1400 24080 1452 24089
rect 2412 24055 2464 24064
rect 2412 24021 2421 24055
rect 2421 24021 2455 24055
rect 2455 24021 2464 24055
rect 2412 24012 2464 24021
rect 2872 24055 2924 24064
rect 2872 24021 2881 24055
rect 2881 24021 2915 24055
rect 2915 24021 2924 24055
rect 2872 24012 2924 24021
rect 3700 24012 3752 24064
rect 5080 24080 5132 24132
rect 6276 24080 6328 24132
rect 7932 24080 7984 24132
rect 8116 24123 8168 24132
rect 8116 24089 8125 24123
rect 8125 24089 8159 24123
rect 8159 24089 8168 24123
rect 8116 24080 8168 24089
rect 10048 24123 10100 24132
rect 10048 24089 10057 24123
rect 10057 24089 10091 24123
rect 10091 24089 10100 24123
rect 10048 24080 10100 24089
rect 10140 24080 10192 24132
rect 12072 24148 12124 24200
rect 3976 24012 4028 24064
rect 4804 24012 4856 24064
rect 6000 24012 6052 24064
rect 6460 24055 6512 24064
rect 6460 24021 6469 24055
rect 6469 24021 6503 24055
rect 6503 24021 6512 24055
rect 6460 24012 6512 24021
rect 7012 24055 7064 24064
rect 7012 24021 7021 24055
rect 7021 24021 7055 24055
rect 7055 24021 7064 24055
rect 7012 24012 7064 24021
rect 7656 24055 7708 24064
rect 7656 24021 7665 24055
rect 7665 24021 7699 24055
rect 7699 24021 7708 24055
rect 7656 24012 7708 24021
rect 8576 24012 8628 24064
rect 11796 24080 11848 24132
rect 14188 24225 14197 24259
rect 14197 24225 14231 24259
rect 14231 24225 14240 24259
rect 14188 24216 14240 24225
rect 13636 24148 13688 24200
rect 18788 24148 18840 24200
rect 19984 24216 20036 24268
rect 21732 24148 21784 24200
rect 29000 24148 29052 24200
rect 38660 24148 38712 24200
rect 11428 24012 11480 24064
rect 14096 24080 14148 24132
rect 19340 24080 19392 24132
rect 20260 24080 20312 24132
rect 27160 24080 27212 24132
rect 35992 24080 36044 24132
rect 14188 24012 14240 24064
rect 15752 24055 15804 24064
rect 15752 24021 15761 24055
rect 15761 24021 15795 24055
rect 15795 24021 15804 24055
rect 15752 24012 15804 24021
rect 16856 24055 16908 24064
rect 16856 24021 16865 24055
rect 16865 24021 16899 24055
rect 16899 24021 16908 24055
rect 16856 24012 16908 24021
rect 17224 24012 17276 24064
rect 29920 24012 29972 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1400 23851 1452 23860
rect 1400 23817 1409 23851
rect 1409 23817 1443 23851
rect 1443 23817 1452 23851
rect 1400 23808 1452 23817
rect 2872 23808 2924 23860
rect 1032 23740 1084 23792
rect 1492 23672 1544 23724
rect 2964 23536 3016 23588
rect 2872 23511 2924 23520
rect 2872 23477 2881 23511
rect 2881 23477 2915 23511
rect 2915 23477 2924 23511
rect 2872 23468 2924 23477
rect 4068 23808 4120 23860
rect 4988 23740 5040 23792
rect 5080 23740 5132 23792
rect 7932 23740 7984 23792
rect 8852 23740 8904 23792
rect 9036 23740 9088 23792
rect 3424 23672 3476 23724
rect 6460 23672 6512 23724
rect 8760 23672 8812 23724
rect 3240 23536 3292 23588
rect 3608 23536 3660 23588
rect 5632 23579 5684 23588
rect 5632 23545 5641 23579
rect 5641 23545 5675 23579
rect 5675 23545 5684 23579
rect 5632 23536 5684 23545
rect 6184 23536 6236 23588
rect 7196 23468 7248 23520
rect 9220 23604 9272 23656
rect 11336 23808 11388 23860
rect 11612 23808 11664 23860
rect 14280 23851 14332 23860
rect 10416 23740 10468 23792
rect 11704 23783 11756 23792
rect 11704 23749 11713 23783
rect 11713 23749 11747 23783
rect 11747 23749 11756 23783
rect 11704 23740 11756 23749
rect 9956 23672 10008 23724
rect 10876 23672 10928 23724
rect 12348 23740 12400 23792
rect 12072 23672 12124 23724
rect 13084 23715 13136 23724
rect 13084 23681 13093 23715
rect 13093 23681 13127 23715
rect 13127 23681 13136 23715
rect 13084 23672 13136 23681
rect 14280 23817 14289 23851
rect 14289 23817 14323 23851
rect 14323 23817 14332 23851
rect 14280 23808 14332 23817
rect 15292 23851 15344 23860
rect 15292 23817 15301 23851
rect 15301 23817 15335 23851
rect 15335 23817 15344 23851
rect 15292 23808 15344 23817
rect 15752 23808 15804 23860
rect 16764 23808 16816 23860
rect 17132 23808 17184 23860
rect 18696 23851 18748 23860
rect 18696 23817 18705 23851
rect 18705 23817 18739 23851
rect 18739 23817 18748 23851
rect 18696 23808 18748 23817
rect 18880 23808 18932 23860
rect 20076 23808 20128 23860
rect 16304 23740 16356 23792
rect 17408 23740 17460 23792
rect 11980 23604 12032 23656
rect 19064 23672 19116 23724
rect 19340 23672 19392 23724
rect 17684 23604 17736 23656
rect 28540 23808 28592 23860
rect 22100 23740 22152 23792
rect 30380 23740 30432 23792
rect 32312 23672 32364 23724
rect 8576 23536 8628 23588
rect 8852 23536 8904 23588
rect 8300 23511 8352 23520
rect 8300 23477 8309 23511
rect 8309 23477 8343 23511
rect 8343 23477 8352 23511
rect 8300 23468 8352 23477
rect 9496 23468 9548 23520
rect 10048 23536 10100 23588
rect 10416 23536 10468 23588
rect 10508 23579 10560 23588
rect 10508 23545 10517 23579
rect 10517 23545 10551 23579
rect 10551 23545 10560 23579
rect 11520 23579 11572 23588
rect 10508 23536 10560 23545
rect 11520 23545 11529 23579
rect 11529 23545 11563 23579
rect 11563 23545 11572 23579
rect 11520 23536 11572 23545
rect 12716 23536 12768 23588
rect 12900 23579 12952 23588
rect 12900 23545 12909 23579
rect 12909 23545 12943 23579
rect 12943 23545 12952 23579
rect 12900 23536 12952 23545
rect 13912 23536 13964 23588
rect 30472 23536 30524 23588
rect 12348 23468 12400 23520
rect 13360 23468 13412 23520
rect 14004 23468 14056 23520
rect 14372 23468 14424 23520
rect 17776 23468 17828 23520
rect 18328 23468 18380 23520
rect 20260 23468 20312 23520
rect 20720 23468 20772 23520
rect 42248 23468 42300 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1676 23264 1728 23316
rect 3240 23307 3292 23316
rect 3240 23273 3249 23307
rect 3249 23273 3283 23307
rect 3283 23273 3292 23307
rect 3240 23264 3292 23273
rect 4896 23264 4948 23316
rect 4988 23264 5040 23316
rect 6276 23264 6328 23316
rect 6644 23264 6696 23316
rect 4528 23196 4580 23248
rect 1584 23128 1636 23180
rect 2136 23128 2188 23180
rect 5540 23196 5592 23248
rect 6920 23196 6972 23248
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 3792 23060 3844 23112
rect 1124 22992 1176 23044
rect 7656 23128 7708 23180
rect 8300 23264 8352 23316
rect 13084 23264 13136 23316
rect 16120 23264 16172 23316
rect 16488 23264 16540 23316
rect 17592 23307 17644 23316
rect 17592 23273 17601 23307
rect 17601 23273 17635 23307
rect 17635 23273 17644 23307
rect 17592 23264 17644 23273
rect 17776 23264 17828 23316
rect 18604 23307 18656 23316
rect 18604 23273 18613 23307
rect 18613 23273 18647 23307
rect 18647 23273 18656 23307
rect 18604 23264 18656 23273
rect 27068 23264 27120 23316
rect 28448 23264 28500 23316
rect 29828 23264 29880 23316
rect 7840 23196 7892 23248
rect 9036 23196 9088 23248
rect 9220 23171 9272 23180
rect 9220 23137 9229 23171
rect 9229 23137 9263 23171
rect 9263 23137 9272 23171
rect 9220 23128 9272 23137
rect 9864 23171 9916 23180
rect 9864 23137 9873 23171
rect 9873 23137 9907 23171
rect 9907 23137 9916 23171
rect 9864 23128 9916 23137
rect 10324 23196 10376 23248
rect 10968 23196 11020 23248
rect 11336 23196 11388 23248
rect 12164 23196 12216 23248
rect 10784 23171 10836 23180
rect 10784 23137 10793 23171
rect 10793 23137 10827 23171
rect 10827 23137 10836 23171
rect 10784 23128 10836 23137
rect 11520 23128 11572 23180
rect 6000 23060 6052 23112
rect 8024 23060 8076 23112
rect 8760 23060 8812 23112
rect 9312 23060 9364 23112
rect 4068 22992 4120 23044
rect 5356 22992 5408 23044
rect 8116 22992 8168 23044
rect 8852 22992 8904 23044
rect 10048 22992 10100 23044
rect 10232 22992 10284 23044
rect 12348 23060 12400 23112
rect 12900 23196 12952 23248
rect 14372 23196 14424 23248
rect 18052 23239 18104 23248
rect 18052 23205 18061 23239
rect 18061 23205 18095 23239
rect 18095 23205 18104 23239
rect 18052 23196 18104 23205
rect 14832 23128 14884 23180
rect 21364 23196 21416 23248
rect 21548 23239 21600 23248
rect 21548 23205 21557 23239
rect 21557 23205 21591 23239
rect 21591 23205 21600 23239
rect 21548 23196 21600 23205
rect 21640 23196 21692 23248
rect 19248 23171 19300 23180
rect 19248 23137 19257 23171
rect 19257 23137 19291 23171
rect 19291 23137 19300 23171
rect 19248 23128 19300 23137
rect 20444 23128 20496 23180
rect 38476 23196 38528 23248
rect 30104 23128 30156 23180
rect 39212 23128 39264 23180
rect 14096 23103 14148 23112
rect 14096 23069 14105 23103
rect 14105 23069 14139 23103
rect 14139 23069 14148 23103
rect 14096 23060 14148 23069
rect 14372 23060 14424 23112
rect 15936 23060 15988 23112
rect 21272 23060 21324 23112
rect 14740 23035 14792 23044
rect 2136 22967 2188 22976
rect 2136 22933 2145 22967
rect 2145 22933 2179 22967
rect 2179 22933 2188 22967
rect 2136 22924 2188 22933
rect 3792 22924 3844 22976
rect 4988 22967 5040 22976
rect 4988 22933 4997 22967
rect 4997 22933 5031 22967
rect 5031 22933 5040 22967
rect 4988 22924 5040 22933
rect 5172 22924 5224 22976
rect 6276 22967 6328 22976
rect 6276 22933 6285 22967
rect 6285 22933 6319 22967
rect 6319 22933 6328 22967
rect 6276 22924 6328 22933
rect 7196 22967 7248 22976
rect 7196 22933 7205 22967
rect 7205 22933 7239 22967
rect 7239 22933 7248 22967
rect 7196 22924 7248 22933
rect 8392 22924 8444 22976
rect 10324 22967 10376 22976
rect 10324 22933 10333 22967
rect 10333 22933 10367 22967
rect 10367 22933 10376 22967
rect 10324 22924 10376 22933
rect 10600 22924 10652 22976
rect 10876 22924 10928 22976
rect 14740 23001 14749 23035
rect 14749 23001 14783 23035
rect 14783 23001 14792 23035
rect 14740 22992 14792 23001
rect 17316 22992 17368 23044
rect 17684 22992 17736 23044
rect 19340 22992 19392 23044
rect 11796 22924 11848 22976
rect 12808 22924 12860 22976
rect 13452 22924 13504 22976
rect 14188 22924 14240 22976
rect 16304 22967 16356 22976
rect 16304 22933 16313 22967
rect 16313 22933 16347 22967
rect 16347 22933 16356 22967
rect 16304 22924 16356 22933
rect 19248 22924 19300 22976
rect 22284 22992 22336 23044
rect 29552 23060 29604 23112
rect 40592 23060 40644 23112
rect 30012 23035 30064 23044
rect 30012 23001 30021 23035
rect 30021 23001 30055 23035
rect 30055 23001 30064 23035
rect 30012 22992 30064 23001
rect 30564 22992 30616 23044
rect 31300 22992 31352 23044
rect 42432 22992 42484 23044
rect 30932 22924 30984 22976
rect 32312 22967 32364 22976
rect 32312 22933 32321 22967
rect 32321 22933 32355 22967
rect 32355 22933 32364 22967
rect 32312 22924 32364 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 1768 22720 1820 22772
rect 2872 22720 2924 22772
rect 4712 22763 4764 22772
rect 4712 22729 4721 22763
rect 4721 22729 4755 22763
rect 4755 22729 4764 22763
rect 4712 22720 4764 22729
rect 5080 22720 5132 22772
rect 5908 22720 5960 22772
rect 7748 22720 7800 22772
rect 480 22652 532 22704
rect 3700 22652 3752 22704
rect 1584 22627 1636 22636
rect 1584 22593 1593 22627
rect 1593 22593 1627 22627
rect 1627 22593 1636 22627
rect 1584 22584 1636 22593
rect 2044 22627 2096 22636
rect 2044 22593 2053 22627
rect 2053 22593 2087 22627
rect 2087 22593 2096 22627
rect 2044 22584 2096 22593
rect 2688 22584 2740 22636
rect 2872 22627 2924 22636
rect 2872 22593 2881 22627
rect 2881 22593 2915 22627
rect 2915 22593 2924 22627
rect 2872 22584 2924 22593
rect 3884 22584 3936 22636
rect 2136 22516 2188 22568
rect 2320 22516 2372 22568
rect 6276 22652 6328 22704
rect 8760 22652 8812 22704
rect 5540 22584 5592 22636
rect 6460 22584 6512 22636
rect 5080 22516 5132 22568
rect 5356 22559 5408 22568
rect 5356 22525 5365 22559
rect 5365 22525 5399 22559
rect 5399 22525 5408 22559
rect 5356 22516 5408 22525
rect 6184 22516 6236 22568
rect 6644 22516 6696 22568
rect 7564 22584 7616 22636
rect 7932 22584 7984 22636
rect 9036 22584 9088 22636
rect 10232 22652 10284 22704
rect 10416 22652 10468 22704
rect 10876 22720 10928 22772
rect 11980 22763 12032 22772
rect 11980 22729 11989 22763
rect 11989 22729 12023 22763
rect 12023 22729 12032 22763
rect 11980 22720 12032 22729
rect 12164 22720 12216 22772
rect 12532 22763 12584 22772
rect 12532 22729 12541 22763
rect 12541 22729 12575 22763
rect 12575 22729 12584 22763
rect 12532 22720 12584 22729
rect 12808 22720 12860 22772
rect 14832 22763 14884 22772
rect 14832 22729 14841 22763
rect 14841 22729 14875 22763
rect 14875 22729 14884 22763
rect 14832 22720 14884 22729
rect 15844 22763 15896 22772
rect 15844 22729 15853 22763
rect 15853 22729 15887 22763
rect 15887 22729 15896 22763
rect 15844 22720 15896 22729
rect 16028 22720 16080 22772
rect 22376 22763 22428 22772
rect 10600 22627 10652 22636
rect 10600 22593 10609 22627
rect 10609 22593 10643 22627
rect 10643 22593 10652 22627
rect 10600 22584 10652 22593
rect 10784 22627 10836 22636
rect 10784 22593 10793 22627
rect 10793 22593 10827 22627
rect 10827 22593 10836 22627
rect 10784 22584 10836 22593
rect 13176 22652 13228 22704
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 12900 22584 12952 22636
rect 13728 22652 13780 22704
rect 13820 22652 13872 22704
rect 14372 22652 14424 22704
rect 17224 22652 17276 22704
rect 21180 22695 21232 22704
rect 21180 22661 21189 22695
rect 21189 22661 21223 22695
rect 21223 22661 21232 22695
rect 21180 22652 21232 22661
rect 13636 22584 13688 22636
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 17868 22627 17920 22636
rect 17868 22593 17877 22627
rect 17877 22593 17911 22627
rect 17911 22593 17920 22627
rect 17868 22584 17920 22593
rect 18236 22584 18288 22636
rect 20168 22627 20220 22636
rect 18144 22559 18196 22568
rect 18144 22525 18153 22559
rect 18153 22525 18187 22559
rect 18187 22525 18196 22559
rect 18144 22516 18196 22525
rect 19892 22559 19944 22568
rect 19892 22525 19901 22559
rect 19901 22525 19935 22559
rect 19935 22525 19944 22559
rect 19892 22516 19944 22525
rect 20168 22593 20177 22627
rect 20177 22593 20211 22627
rect 20211 22593 20220 22627
rect 20168 22584 20220 22593
rect 22376 22729 22385 22763
rect 22385 22729 22419 22763
rect 22419 22729 22428 22763
rect 22376 22720 22428 22729
rect 29828 22763 29880 22772
rect 29828 22729 29837 22763
rect 29837 22729 29871 22763
rect 29871 22729 29880 22763
rect 29828 22720 29880 22729
rect 30012 22720 30064 22772
rect 30104 22720 30156 22772
rect 34704 22720 34756 22772
rect 22192 22652 22244 22704
rect 22560 22584 22612 22636
rect 29184 22516 29236 22568
rect 1400 22423 1452 22432
rect 1400 22389 1409 22423
rect 1409 22389 1443 22423
rect 1443 22389 1452 22423
rect 1400 22380 1452 22389
rect 4068 22423 4120 22432
rect 4068 22389 4077 22423
rect 4077 22389 4111 22423
rect 4111 22389 4120 22423
rect 4068 22380 4120 22389
rect 7196 22448 7248 22500
rect 10416 22448 10468 22500
rect 10876 22448 10928 22500
rect 11060 22448 11112 22500
rect 11888 22491 11940 22500
rect 11888 22457 11897 22491
rect 11897 22457 11931 22491
rect 11931 22457 11940 22491
rect 11888 22448 11940 22457
rect 12624 22448 12676 22500
rect 21088 22448 21140 22500
rect 21272 22448 21324 22500
rect 26240 22448 26292 22500
rect 6000 22380 6052 22432
rect 6092 22380 6144 22432
rect 6460 22380 6512 22432
rect 8668 22380 8720 22432
rect 10784 22380 10836 22432
rect 12716 22423 12768 22432
rect 12716 22389 12725 22423
rect 12725 22389 12759 22423
rect 12759 22389 12768 22423
rect 12716 22380 12768 22389
rect 13912 22380 13964 22432
rect 15568 22380 15620 22432
rect 16028 22380 16080 22432
rect 30564 22423 30616 22432
rect 30564 22389 30573 22423
rect 30573 22389 30607 22423
rect 30607 22389 30616 22423
rect 30564 22380 30616 22389
rect 31300 22423 31352 22432
rect 31300 22389 31309 22423
rect 31309 22389 31343 22423
rect 31343 22389 31352 22423
rect 31300 22380 31352 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3424 22176 3476 22228
rect 5540 22176 5592 22228
rect 6000 22176 6052 22228
rect 6920 22219 6972 22228
rect 6920 22185 6929 22219
rect 6929 22185 6963 22219
rect 6963 22185 6972 22219
rect 6920 22176 6972 22185
rect 7564 22176 7616 22228
rect 10784 22176 10836 22228
rect 10968 22219 11020 22228
rect 10968 22185 10977 22219
rect 10977 22185 11011 22219
rect 11011 22185 11020 22219
rect 10968 22176 11020 22185
rect 1952 22108 2004 22160
rect 2596 22108 2648 22160
rect 3240 22108 3292 22160
rect 5632 22151 5684 22160
rect 2228 22015 2280 22024
rect 2228 21981 2237 22015
rect 2237 21981 2271 22015
rect 2271 21981 2280 22015
rect 2964 22040 3016 22092
rect 3148 22040 3200 22092
rect 3700 22040 3752 22092
rect 3792 22083 3844 22092
rect 3792 22049 3801 22083
rect 3801 22049 3835 22083
rect 3835 22049 3844 22083
rect 3792 22040 3844 22049
rect 5264 22040 5316 22092
rect 2228 21972 2280 21981
rect 2780 21972 2832 22024
rect 3516 21972 3568 22024
rect 4712 21972 4764 22024
rect 5632 22117 5641 22151
rect 5641 22117 5675 22151
rect 5675 22117 5684 22151
rect 5632 22108 5684 22117
rect 14648 22176 14700 22228
rect 11152 22108 11204 22160
rect 12900 22108 12952 22160
rect 13452 22108 13504 22160
rect 15200 22108 15252 22160
rect 22192 22176 22244 22228
rect 5724 22083 5776 22092
rect 5724 22049 5733 22083
rect 5733 22049 5767 22083
rect 5767 22049 5776 22083
rect 5724 22040 5776 22049
rect 6184 22040 6236 22092
rect 10324 22083 10376 22092
rect 10324 22049 10333 22083
rect 10333 22049 10367 22083
rect 10367 22049 10376 22083
rect 10324 22040 10376 22049
rect 10416 22040 10468 22092
rect 10692 22040 10744 22092
rect 15384 22083 15436 22092
rect 7564 21972 7616 22024
rect 7932 22015 7984 22024
rect 7932 21981 7941 22015
rect 7941 21981 7975 22015
rect 7975 21981 7984 22015
rect 7932 21972 7984 21981
rect 8116 21972 8168 22024
rect 8484 21972 8536 22024
rect 1860 21904 1912 21956
rect 1584 21879 1636 21888
rect 1584 21845 1593 21879
rect 1593 21845 1627 21879
rect 1627 21845 1636 21879
rect 1584 21836 1636 21845
rect 1676 21836 1728 21888
rect 2228 21836 2280 21888
rect 3148 21904 3200 21956
rect 5080 21904 5132 21956
rect 5172 21904 5224 21956
rect 5540 21904 5592 21956
rect 8944 21904 8996 21956
rect 12072 21972 12124 22024
rect 12348 22015 12400 22024
rect 12348 21981 12357 22015
rect 12357 21981 12391 22015
rect 12391 21981 12400 22015
rect 12348 21972 12400 21981
rect 12716 21972 12768 22024
rect 3516 21836 3568 21888
rect 6276 21836 6328 21888
rect 6920 21836 6972 21888
rect 8300 21836 8352 21888
rect 9128 21836 9180 21888
rect 10048 21836 10100 21888
rect 10508 21879 10560 21888
rect 10508 21845 10517 21879
rect 10517 21845 10551 21879
rect 10551 21845 10560 21879
rect 10508 21836 10560 21845
rect 10600 21879 10652 21888
rect 10600 21845 10609 21879
rect 10609 21845 10643 21879
rect 10643 21845 10652 21879
rect 10600 21836 10652 21845
rect 10968 21836 11020 21888
rect 11612 21904 11664 21956
rect 12624 21904 12676 21956
rect 14096 22015 14148 22024
rect 14096 21981 14105 22015
rect 14105 21981 14139 22015
rect 14139 21981 14148 22015
rect 14096 21972 14148 21981
rect 14832 21972 14884 22024
rect 15384 22049 15393 22083
rect 15393 22049 15427 22083
rect 15427 22049 15436 22083
rect 15384 22040 15436 22049
rect 16304 22040 16356 22092
rect 16764 22040 16816 22092
rect 17408 22040 17460 22092
rect 16856 22015 16908 22024
rect 15200 21904 15252 21956
rect 16856 21981 16865 22015
rect 16865 21981 16899 22015
rect 16899 21981 16908 22015
rect 16856 21972 16908 21981
rect 18144 21972 18196 22024
rect 26148 22108 26200 22160
rect 18420 22040 18472 22092
rect 19064 22040 19116 22092
rect 19340 22040 19392 22092
rect 19432 22040 19484 22092
rect 20536 22083 20588 22092
rect 20536 22049 20545 22083
rect 20545 22049 20579 22083
rect 20579 22049 20588 22083
rect 20536 22040 20588 22049
rect 20260 21972 20312 22024
rect 31300 21972 31352 22024
rect 17776 21904 17828 21956
rect 18328 21947 18380 21956
rect 18328 21913 18337 21947
rect 18337 21913 18371 21947
rect 18371 21913 18380 21947
rect 18328 21904 18380 21913
rect 19248 21904 19300 21956
rect 11888 21879 11940 21888
rect 11888 21845 11897 21879
rect 11897 21845 11931 21879
rect 11931 21845 11940 21879
rect 11888 21836 11940 21845
rect 12808 21879 12860 21888
rect 12808 21845 12817 21879
rect 12817 21845 12851 21879
rect 12851 21845 12860 21879
rect 12808 21836 12860 21845
rect 12900 21836 12952 21888
rect 13176 21836 13228 21888
rect 15752 21836 15804 21888
rect 17408 21836 17460 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2596 21632 2648 21684
rect 4068 21632 4120 21684
rect 1492 21539 1544 21548
rect 1492 21505 1501 21539
rect 1501 21505 1535 21539
rect 1535 21505 1544 21539
rect 1492 21496 1544 21505
rect 2504 21496 2556 21548
rect 3056 21496 3108 21548
rect 3792 21496 3844 21548
rect 5908 21632 5960 21684
rect 5356 21564 5408 21616
rect 6644 21607 6696 21616
rect 6644 21573 6653 21607
rect 6653 21573 6687 21607
rect 6687 21573 6696 21607
rect 6644 21564 6696 21573
rect 5448 21539 5500 21548
rect 5448 21505 5457 21539
rect 5457 21505 5491 21539
rect 5491 21505 5500 21539
rect 5448 21496 5500 21505
rect 1492 21360 1544 21412
rect 3884 21292 3936 21344
rect 5172 21428 5224 21480
rect 5264 21428 5316 21480
rect 10324 21632 10376 21684
rect 11336 21632 11388 21684
rect 11612 21632 11664 21684
rect 12624 21632 12676 21684
rect 13176 21675 13228 21684
rect 13176 21641 13185 21675
rect 13185 21641 13219 21675
rect 13219 21641 13228 21675
rect 13176 21632 13228 21641
rect 13360 21632 13412 21684
rect 23756 21632 23808 21684
rect 27712 21675 27764 21684
rect 27712 21641 27721 21675
rect 27721 21641 27755 21675
rect 27755 21641 27764 21675
rect 27712 21632 27764 21641
rect 11796 21564 11848 21616
rect 12256 21564 12308 21616
rect 14556 21564 14608 21616
rect 17316 21564 17368 21616
rect 19892 21564 19944 21616
rect 22284 21564 22336 21616
rect 22928 21607 22980 21616
rect 22928 21573 22937 21607
rect 22937 21573 22971 21607
rect 22971 21573 22980 21607
rect 22928 21564 22980 21573
rect 23112 21564 23164 21616
rect 9496 21539 9548 21548
rect 9496 21505 9505 21539
rect 9505 21505 9539 21539
rect 9539 21505 9548 21539
rect 9496 21496 9548 21505
rect 9680 21496 9732 21548
rect 8024 21471 8076 21480
rect 8024 21437 8033 21471
rect 8033 21437 8067 21471
rect 8067 21437 8076 21471
rect 8024 21428 8076 21437
rect 4620 21292 4672 21344
rect 4712 21292 4764 21344
rect 5264 21292 5316 21344
rect 8300 21360 8352 21412
rect 8392 21360 8444 21412
rect 9128 21360 9180 21412
rect 10416 21360 10468 21412
rect 10692 21496 10744 21548
rect 12164 21496 12216 21548
rect 12440 21496 12492 21548
rect 14280 21496 14332 21548
rect 15476 21539 15528 21548
rect 15476 21505 15485 21539
rect 15485 21505 15519 21539
rect 15519 21505 15528 21539
rect 15476 21496 15528 21505
rect 16948 21539 17000 21548
rect 16948 21505 16957 21539
rect 16957 21505 16991 21539
rect 16991 21505 17000 21539
rect 16948 21496 17000 21505
rect 17960 21496 18012 21548
rect 20628 21539 20680 21548
rect 20628 21505 20637 21539
rect 20637 21505 20671 21539
rect 20671 21505 20680 21539
rect 20628 21496 20680 21505
rect 12072 21471 12124 21480
rect 12072 21437 12081 21471
rect 12081 21437 12115 21471
rect 12115 21437 12124 21471
rect 12072 21428 12124 21437
rect 12624 21428 12676 21480
rect 14372 21428 14424 21480
rect 15384 21428 15436 21480
rect 16672 21471 16724 21480
rect 16672 21437 16681 21471
rect 16681 21437 16715 21471
rect 16715 21437 16724 21471
rect 16672 21428 16724 21437
rect 16764 21428 16816 21480
rect 31208 21496 31260 21548
rect 23480 21428 23532 21480
rect 12164 21360 12216 21412
rect 13176 21360 13228 21412
rect 8208 21292 8260 21344
rect 10232 21292 10284 21344
rect 11980 21292 12032 21344
rect 14372 21335 14424 21344
rect 14372 21301 14381 21335
rect 14381 21301 14415 21335
rect 14415 21301 14424 21335
rect 16212 21360 16264 21412
rect 27804 21360 27856 21412
rect 14372 21292 14424 21301
rect 16948 21292 17000 21344
rect 18236 21292 18288 21344
rect 18420 21292 18472 21344
rect 19248 21292 19300 21344
rect 20444 21292 20496 21344
rect 21732 21292 21784 21344
rect 22284 21292 22336 21344
rect 23480 21335 23532 21344
rect 23480 21301 23489 21335
rect 23489 21301 23523 21335
rect 23523 21301 23532 21335
rect 23480 21292 23532 21301
rect 23664 21292 23716 21344
rect 24124 21335 24176 21344
rect 24124 21301 24133 21335
rect 24133 21301 24167 21335
rect 24167 21301 24176 21335
rect 24124 21292 24176 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 388 21088 440 21140
rect 2044 21088 2096 21140
rect 3056 21088 3108 21140
rect 3332 21088 3384 21140
rect 4620 21088 4672 21140
rect 4436 21020 4488 21072
rect 5080 21088 5132 21140
rect 8392 21131 8444 21140
rect 8392 21097 8401 21131
rect 8401 21097 8435 21131
rect 8435 21097 8444 21131
rect 8392 21088 8444 21097
rect 8852 21088 8904 21140
rect 10692 21088 10744 21140
rect 11336 21088 11388 21140
rect 12716 21088 12768 21140
rect 13360 21088 13412 21140
rect 14372 21088 14424 21140
rect 1952 20884 2004 20936
rect 2136 20927 2188 20936
rect 2136 20893 2145 20927
rect 2145 20893 2179 20927
rect 2179 20893 2188 20927
rect 2136 20884 2188 20893
rect 4804 20952 4856 21004
rect 5724 21020 5776 21072
rect 8024 21020 8076 21072
rect 11612 21020 11664 21072
rect 15660 21063 15712 21072
rect 15660 21029 15669 21063
rect 15669 21029 15703 21063
rect 15703 21029 15712 21063
rect 15660 21020 15712 21029
rect 15844 21131 15896 21140
rect 15844 21097 15853 21131
rect 15853 21097 15887 21131
rect 15887 21097 15896 21131
rect 15844 21088 15896 21097
rect 16580 21063 16632 21072
rect 16580 21029 16589 21063
rect 16589 21029 16623 21063
rect 16623 21029 16632 21063
rect 16580 21020 16632 21029
rect 21364 21088 21416 21140
rect 25320 21088 25372 21140
rect 26608 21131 26660 21140
rect 26608 21097 26617 21131
rect 26617 21097 26651 21131
rect 26651 21097 26660 21131
rect 26608 21088 26660 21097
rect 28080 21131 28132 21140
rect 17500 21063 17552 21072
rect 17500 21029 17509 21063
rect 17509 21029 17543 21063
rect 17543 21029 17552 21063
rect 17500 21020 17552 21029
rect 18052 21020 18104 21072
rect 19800 21020 19852 21072
rect 3056 20816 3108 20868
rect 1308 20748 1360 20800
rect 4344 20816 4396 20868
rect 3884 20748 3936 20800
rect 4712 20748 4764 20800
rect 5448 20952 5500 21004
rect 6368 20952 6420 21004
rect 6460 20952 6512 21004
rect 6644 20952 6696 21004
rect 5540 20884 5592 20936
rect 9312 20952 9364 21004
rect 9404 20952 9456 21004
rect 12716 20995 12768 21004
rect 12716 20961 12725 20995
rect 12725 20961 12759 20995
rect 12759 20961 12768 20995
rect 12716 20952 12768 20961
rect 13360 20952 13412 21004
rect 14648 20995 14700 21004
rect 14648 20961 14657 20995
rect 14657 20961 14691 20995
rect 14691 20961 14700 20995
rect 14648 20952 14700 20961
rect 16212 20952 16264 21004
rect 16488 20952 16540 21004
rect 16764 20995 16816 21004
rect 16764 20961 16773 20995
rect 16773 20961 16807 20995
rect 16807 20961 16816 20995
rect 16764 20952 16816 20961
rect 18512 20952 18564 21004
rect 18880 20952 18932 21004
rect 8300 20884 8352 20936
rect 10784 20927 10836 20936
rect 10784 20893 10793 20927
rect 10793 20893 10827 20927
rect 10827 20893 10836 20927
rect 10784 20884 10836 20893
rect 12072 20927 12124 20936
rect 12072 20893 12081 20927
rect 12081 20893 12115 20927
rect 12115 20893 12124 20927
rect 12072 20884 12124 20893
rect 12808 20927 12860 20936
rect 12808 20893 12817 20927
rect 12817 20893 12851 20927
rect 12851 20893 12860 20927
rect 12808 20884 12860 20893
rect 13176 20884 13228 20936
rect 19156 20884 19208 20936
rect 6460 20816 6512 20868
rect 7288 20859 7340 20868
rect 7288 20825 7322 20859
rect 7322 20825 7340 20859
rect 7288 20816 7340 20825
rect 7932 20816 7984 20868
rect 8392 20816 8444 20868
rect 8852 20816 8904 20868
rect 9772 20816 9824 20868
rect 11612 20816 11664 20868
rect 13544 20816 13596 20868
rect 15292 20816 15344 20868
rect 15476 20816 15528 20868
rect 16580 20816 16632 20868
rect 17132 20816 17184 20868
rect 19064 20816 19116 20868
rect 13176 20748 13228 20800
rect 13360 20748 13412 20800
rect 19892 20884 19944 20936
rect 23204 21020 23256 21072
rect 24032 21020 24084 21072
rect 20444 20952 20496 21004
rect 22652 20952 22704 21004
rect 28080 21097 28089 21131
rect 28089 21097 28123 21131
rect 28123 21097 28132 21131
rect 28080 21088 28132 21097
rect 32220 20952 32272 21004
rect 25964 20884 26016 20936
rect 19340 20859 19392 20868
rect 19340 20825 19349 20859
rect 19349 20825 19383 20859
rect 19383 20825 19392 20859
rect 19340 20816 19392 20825
rect 19984 20816 20036 20868
rect 23204 20816 23256 20868
rect 24768 20816 24820 20868
rect 25688 20816 25740 20868
rect 26884 20816 26936 20868
rect 20536 20748 20588 20800
rect 20904 20791 20956 20800
rect 20904 20757 20913 20791
rect 20913 20757 20947 20791
rect 20947 20757 20956 20791
rect 20904 20748 20956 20757
rect 21456 20791 21508 20800
rect 21456 20757 21465 20791
rect 21465 20757 21499 20791
rect 21499 20757 21508 20791
rect 21456 20748 21508 20757
rect 22192 20748 22244 20800
rect 22468 20748 22520 20800
rect 22652 20791 22704 20800
rect 22652 20757 22661 20791
rect 22661 20757 22695 20791
rect 22695 20757 22704 20791
rect 22652 20748 22704 20757
rect 23296 20748 23348 20800
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 24492 20791 24544 20800
rect 24492 20757 24501 20791
rect 24501 20757 24535 20791
rect 24535 20757 24544 20791
rect 24492 20748 24544 20757
rect 29092 20748 29144 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1216 20544 1268 20596
rect 4344 20544 4396 20596
rect 6368 20544 6420 20596
rect 6552 20587 6604 20596
rect 6552 20553 6561 20587
rect 6561 20553 6595 20587
rect 6595 20553 6604 20587
rect 6552 20544 6604 20553
rect 6644 20544 6696 20596
rect 7012 20544 7064 20596
rect 7564 20544 7616 20596
rect 9128 20544 9180 20596
rect 9588 20544 9640 20596
rect 11704 20544 11756 20596
rect 11520 20476 11572 20528
rect 2320 20408 2372 20460
rect 2504 20408 2556 20460
rect 2596 20408 2648 20460
rect 3608 20408 3660 20460
rect 4252 20451 4304 20460
rect 4252 20417 4261 20451
rect 4261 20417 4295 20451
rect 4295 20417 4304 20451
rect 4252 20408 4304 20417
rect 2044 20340 2096 20392
rect 5172 20408 5224 20460
rect 5540 20451 5592 20460
rect 5540 20417 5549 20451
rect 5549 20417 5583 20451
rect 5583 20417 5592 20451
rect 5540 20408 5592 20417
rect 5816 20451 5868 20460
rect 5816 20417 5825 20451
rect 5825 20417 5859 20451
rect 5859 20417 5868 20451
rect 5816 20408 5868 20417
rect 6644 20451 6696 20460
rect 6644 20417 6653 20451
rect 6653 20417 6687 20451
rect 6687 20417 6696 20451
rect 6644 20408 6696 20417
rect 4528 20383 4580 20392
rect 4528 20349 4537 20383
rect 4537 20349 4571 20383
rect 4571 20349 4580 20383
rect 4528 20340 4580 20349
rect 6184 20340 6236 20392
rect 2320 20315 2372 20324
rect 2320 20281 2329 20315
rect 2329 20281 2363 20315
rect 2363 20281 2372 20315
rect 2320 20272 2372 20281
rect 3148 20315 3200 20324
rect 3148 20281 3157 20315
rect 3157 20281 3191 20315
rect 3191 20281 3200 20315
rect 3148 20272 3200 20281
rect 3424 20272 3476 20324
rect 9128 20408 9180 20460
rect 9312 20408 9364 20460
rect 9772 20451 9824 20460
rect 8852 20383 8904 20392
rect 8852 20349 8861 20383
rect 8861 20349 8895 20383
rect 8895 20349 8904 20383
rect 8852 20340 8904 20349
rect 2688 20204 2740 20256
rect 3056 20204 3108 20256
rect 4804 20204 4856 20256
rect 9772 20417 9781 20451
rect 9781 20417 9815 20451
rect 9815 20417 9824 20451
rect 9772 20408 9824 20417
rect 10692 20408 10744 20460
rect 16028 20476 16080 20528
rect 18052 20544 18104 20596
rect 18972 20587 19024 20596
rect 18328 20476 18380 20528
rect 18512 20519 18564 20528
rect 18512 20485 18521 20519
rect 18521 20485 18555 20519
rect 18555 20485 18564 20519
rect 18512 20476 18564 20485
rect 18972 20553 18981 20587
rect 18981 20553 19015 20587
rect 19015 20553 19024 20587
rect 18972 20544 19024 20553
rect 20444 20587 20496 20596
rect 20444 20553 20453 20587
rect 20453 20553 20487 20587
rect 20487 20553 20496 20587
rect 20444 20544 20496 20553
rect 20812 20544 20864 20596
rect 22652 20587 22704 20596
rect 22652 20553 22661 20587
rect 22661 20553 22695 20587
rect 22695 20553 22704 20587
rect 22652 20544 22704 20553
rect 24216 20587 24268 20596
rect 24216 20553 24225 20587
rect 24225 20553 24259 20587
rect 24259 20553 24268 20587
rect 24216 20544 24268 20553
rect 25780 20587 25832 20596
rect 25780 20553 25789 20587
rect 25789 20553 25823 20587
rect 25823 20553 25832 20587
rect 25780 20544 25832 20553
rect 28356 20587 28408 20596
rect 28356 20553 28365 20587
rect 28365 20553 28399 20587
rect 28399 20553 28408 20587
rect 28356 20544 28408 20553
rect 29736 20587 29788 20596
rect 29736 20553 29745 20587
rect 29745 20553 29779 20587
rect 29779 20553 29788 20587
rect 29736 20544 29788 20553
rect 24492 20476 24544 20528
rect 25320 20476 25372 20528
rect 27712 20476 27764 20528
rect 10416 20340 10468 20392
rect 12992 20408 13044 20460
rect 13820 20408 13872 20460
rect 14832 20408 14884 20460
rect 15016 20408 15068 20460
rect 11152 20340 11204 20392
rect 13544 20340 13596 20392
rect 13636 20340 13688 20392
rect 14648 20340 14700 20392
rect 18144 20408 18196 20460
rect 16120 20340 16172 20392
rect 17224 20340 17276 20392
rect 17500 20340 17552 20392
rect 17960 20272 18012 20324
rect 20904 20408 20956 20460
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 25780 20408 25832 20460
rect 27252 20408 27304 20460
rect 29092 20451 29144 20460
rect 29092 20417 29101 20451
rect 29101 20417 29135 20451
rect 29135 20417 29144 20451
rect 29092 20408 29144 20417
rect 19524 20340 19576 20392
rect 21640 20340 21692 20392
rect 33600 20340 33652 20392
rect 21916 20272 21968 20324
rect 16488 20204 16540 20256
rect 17132 20247 17184 20256
rect 17132 20213 17141 20247
rect 17141 20213 17175 20247
rect 17175 20213 17184 20247
rect 17132 20204 17184 20213
rect 17224 20204 17276 20256
rect 18696 20204 18748 20256
rect 20904 20204 20956 20256
rect 24860 20247 24912 20256
rect 24860 20213 24869 20247
rect 24869 20213 24903 20247
rect 24903 20213 24912 20247
rect 24860 20204 24912 20213
rect 27436 20247 27488 20256
rect 27436 20213 27445 20247
rect 27445 20213 27479 20247
rect 27479 20213 27488 20247
rect 27436 20204 27488 20213
rect 33784 20204 33836 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2136 20000 2188 20052
rect 3240 20043 3292 20052
rect 3240 20009 3249 20043
rect 3249 20009 3283 20043
rect 3283 20009 3292 20043
rect 3240 20000 3292 20009
rect 4712 20000 4764 20052
rect 5172 20000 5224 20052
rect 6644 20000 6696 20052
rect 9680 20000 9732 20052
rect 10692 20000 10744 20052
rect 18144 20000 18196 20052
rect 18420 20000 18472 20052
rect 18972 20000 19024 20052
rect 19156 20000 19208 20052
rect 20444 20000 20496 20052
rect 22192 20000 22244 20052
rect 25596 20000 25648 20052
rect 1952 19975 2004 19984
rect 1952 19941 1961 19975
rect 1961 19941 1995 19975
rect 1995 19941 2004 19975
rect 1952 19932 2004 19941
rect 2504 19932 2556 19984
rect 6184 19932 6236 19984
rect 6368 19932 6420 19984
rect 2044 19864 2096 19916
rect 2872 19864 2924 19916
rect 3792 19864 3844 19916
rect 4896 19864 4948 19916
rect 3332 19796 3384 19848
rect 4712 19796 4764 19848
rect 2044 19728 2096 19780
rect 5356 19796 5408 19848
rect 3332 19660 3384 19712
rect 4160 19660 4212 19712
rect 6736 19864 6788 19916
rect 7288 19907 7340 19916
rect 7288 19873 7297 19907
rect 7297 19873 7331 19907
rect 7331 19873 7340 19907
rect 7288 19864 7340 19873
rect 8852 19932 8904 19984
rect 16764 19932 16816 19984
rect 17408 19932 17460 19984
rect 17868 19932 17920 19984
rect 28172 20000 28224 20052
rect 32772 20043 32824 20052
rect 32772 20009 32781 20043
rect 32781 20009 32815 20043
rect 32815 20009 32824 20043
rect 32772 20000 32824 20009
rect 9404 19864 9456 19916
rect 11060 19864 11112 19916
rect 11796 19907 11848 19916
rect 11796 19873 11805 19907
rect 11805 19873 11839 19907
rect 11839 19873 11848 19907
rect 11796 19864 11848 19873
rect 13268 19907 13320 19916
rect 13268 19873 13277 19907
rect 13277 19873 13311 19907
rect 13311 19873 13320 19907
rect 13268 19864 13320 19873
rect 14372 19907 14424 19916
rect 14372 19873 14381 19907
rect 14381 19873 14415 19907
rect 14415 19873 14424 19907
rect 14372 19864 14424 19873
rect 15108 19864 15160 19916
rect 16212 19907 16264 19916
rect 16212 19873 16221 19907
rect 16221 19873 16255 19907
rect 16255 19873 16264 19907
rect 16212 19864 16264 19873
rect 16488 19864 16540 19916
rect 18236 19864 18288 19916
rect 20996 19864 21048 19916
rect 27160 19932 27212 19984
rect 28448 19932 28500 19984
rect 28816 19932 28868 19984
rect 30656 19975 30708 19984
rect 30656 19941 30665 19975
rect 30665 19941 30699 19975
rect 30699 19941 30708 19975
rect 30656 19932 30708 19941
rect 37832 20000 37884 20052
rect 22836 19864 22888 19916
rect 43628 19932 43680 19984
rect 43536 19864 43588 19916
rect 6092 19839 6144 19848
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 6368 19796 6420 19848
rect 8852 19796 8904 19848
rect 12348 19796 12400 19848
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 14096 19839 14148 19848
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 14832 19796 14884 19848
rect 5816 19728 5868 19780
rect 6736 19771 6788 19780
rect 6736 19737 6745 19771
rect 6745 19737 6779 19771
rect 6779 19737 6788 19771
rect 6736 19728 6788 19737
rect 9128 19771 9180 19780
rect 9128 19737 9137 19771
rect 9137 19737 9171 19771
rect 9171 19737 9180 19771
rect 9128 19728 9180 19737
rect 16212 19728 16264 19780
rect 16856 19728 16908 19780
rect 5540 19660 5592 19712
rect 7104 19660 7156 19712
rect 7196 19660 7248 19712
rect 8760 19660 8812 19712
rect 13544 19660 13596 19712
rect 16580 19660 16632 19712
rect 16672 19660 16724 19712
rect 17500 19728 17552 19780
rect 18604 19796 18656 19848
rect 20168 19796 20220 19848
rect 20628 19839 20680 19848
rect 20628 19805 20637 19839
rect 20637 19805 20671 19839
rect 20671 19805 20680 19839
rect 20628 19796 20680 19805
rect 21272 19796 21324 19848
rect 23388 19796 23440 19848
rect 24952 19796 25004 19848
rect 28356 19796 28408 19848
rect 29736 19796 29788 19848
rect 21548 19728 21600 19780
rect 23480 19771 23532 19780
rect 23480 19737 23489 19771
rect 23489 19737 23523 19771
rect 23523 19737 23532 19771
rect 23480 19728 23532 19737
rect 25044 19771 25096 19780
rect 25044 19737 25053 19771
rect 25053 19737 25087 19771
rect 25087 19737 25096 19771
rect 25044 19728 25096 19737
rect 26884 19771 26936 19780
rect 18144 19703 18196 19712
rect 18144 19669 18153 19703
rect 18153 19669 18187 19703
rect 18187 19669 18196 19703
rect 18144 19660 18196 19669
rect 18328 19660 18380 19712
rect 21180 19660 21232 19712
rect 21640 19660 21692 19712
rect 24768 19660 24820 19712
rect 26884 19737 26893 19771
rect 26893 19737 26927 19771
rect 26927 19737 26936 19771
rect 26884 19728 26936 19737
rect 27620 19771 27672 19780
rect 27620 19737 27629 19771
rect 27629 19737 27663 19771
rect 27663 19737 27672 19771
rect 27620 19728 27672 19737
rect 28448 19728 28500 19780
rect 30196 19771 30248 19780
rect 27160 19660 27212 19712
rect 28632 19703 28684 19712
rect 28632 19669 28641 19703
rect 28641 19669 28675 19703
rect 28675 19669 28684 19703
rect 28632 19660 28684 19669
rect 30196 19737 30205 19771
rect 30205 19737 30239 19771
rect 30239 19737 30248 19771
rect 30196 19728 30248 19737
rect 33416 19796 33468 19848
rect 43352 19796 43404 19848
rect 33784 19771 33836 19780
rect 31392 19703 31444 19712
rect 31392 19669 31401 19703
rect 31401 19669 31435 19703
rect 31435 19669 31444 19703
rect 31392 19660 31444 19669
rect 32036 19703 32088 19712
rect 32036 19669 32045 19703
rect 32045 19669 32079 19703
rect 32079 19669 32088 19703
rect 33784 19737 33793 19771
rect 33793 19737 33827 19771
rect 33827 19737 33836 19771
rect 33784 19728 33836 19737
rect 34612 19728 34664 19780
rect 35624 19728 35676 19780
rect 32036 19660 32088 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1952 19456 2004 19508
rect 2504 19499 2556 19508
rect 2504 19465 2513 19499
rect 2513 19465 2547 19499
rect 2547 19465 2556 19499
rect 2504 19456 2556 19465
rect 5632 19456 5684 19508
rect 5816 19499 5868 19508
rect 5816 19465 5825 19499
rect 5825 19465 5859 19499
rect 5859 19465 5868 19499
rect 5816 19456 5868 19465
rect 2320 19388 2372 19440
rect 1860 19320 1912 19372
rect 2136 19320 2188 19372
rect 2412 19363 2464 19372
rect 2412 19329 2421 19363
rect 2421 19329 2455 19363
rect 2455 19329 2464 19363
rect 2412 19320 2464 19329
rect 3424 19320 3476 19372
rect 3700 19320 3752 19372
rect 5540 19388 5592 19440
rect 5724 19388 5776 19440
rect 8484 19431 8536 19440
rect 8484 19397 8493 19431
rect 8493 19397 8527 19431
rect 8527 19397 8536 19431
rect 8484 19388 8536 19397
rect 2688 19295 2740 19304
rect 2688 19261 2697 19295
rect 2697 19261 2731 19295
rect 2731 19261 2740 19295
rect 2688 19252 2740 19261
rect 3792 19252 3844 19304
rect 4344 19252 4396 19304
rect 4160 19184 4212 19236
rect 4252 19184 4304 19236
rect 1952 19116 2004 19168
rect 3332 19116 3384 19168
rect 6460 19320 6512 19372
rect 8944 19456 8996 19508
rect 8760 19388 8812 19440
rect 13544 19388 13596 19440
rect 19432 19456 19484 19508
rect 5632 19252 5684 19304
rect 9404 19252 9456 19304
rect 11520 19295 11572 19304
rect 11520 19261 11529 19295
rect 11529 19261 11563 19295
rect 11563 19261 11572 19295
rect 11520 19252 11572 19261
rect 13544 19252 13596 19304
rect 14740 19388 14792 19440
rect 6092 19184 6144 19236
rect 6644 19184 6696 19236
rect 8116 19184 8168 19236
rect 9588 19184 9640 19236
rect 10876 19184 10928 19236
rect 13636 19184 13688 19236
rect 4620 19116 4672 19168
rect 5908 19116 5960 19168
rect 9772 19116 9824 19168
rect 13268 19116 13320 19168
rect 13544 19116 13596 19168
rect 15016 19320 15068 19372
rect 15200 19363 15252 19372
rect 15200 19329 15209 19363
rect 15209 19329 15243 19363
rect 15243 19329 15252 19363
rect 15200 19320 15252 19329
rect 16028 19320 16080 19372
rect 16120 19320 16172 19372
rect 19248 19388 19300 19440
rect 19616 19388 19668 19440
rect 19984 19388 20036 19440
rect 20444 19388 20496 19440
rect 21088 19431 21140 19440
rect 21088 19397 21097 19431
rect 21097 19397 21131 19431
rect 21131 19397 21140 19431
rect 21088 19388 21140 19397
rect 21364 19388 21416 19440
rect 23572 19388 23624 19440
rect 15108 19252 15160 19304
rect 15292 19252 15344 19304
rect 16488 19252 16540 19304
rect 18328 19320 18380 19372
rect 18512 19320 18564 19372
rect 19432 19320 19484 19372
rect 19892 19320 19944 19372
rect 22744 19320 22796 19372
rect 23664 19320 23716 19372
rect 28448 19456 28500 19508
rect 28724 19499 28776 19508
rect 28724 19465 28733 19499
rect 28733 19465 28767 19499
rect 28767 19465 28776 19499
rect 28724 19456 28776 19465
rect 29460 19499 29512 19508
rect 29460 19465 29469 19499
rect 29469 19465 29503 19499
rect 29503 19465 29512 19499
rect 29460 19456 29512 19465
rect 33140 19499 33192 19508
rect 33140 19465 33149 19499
rect 33149 19465 33183 19499
rect 33183 19465 33192 19499
rect 33140 19456 33192 19465
rect 33324 19388 33376 19440
rect 26700 19320 26752 19372
rect 27344 19320 27396 19372
rect 28908 19320 28960 19372
rect 30196 19320 30248 19372
rect 31760 19320 31812 19372
rect 32036 19320 32088 19372
rect 32404 19320 32456 19372
rect 33968 19320 34020 19372
rect 19156 19252 19208 19304
rect 19616 19252 19668 19304
rect 19984 19252 20036 19304
rect 21824 19295 21876 19304
rect 21824 19261 21833 19295
rect 21833 19261 21867 19295
rect 21867 19261 21876 19295
rect 21824 19252 21876 19261
rect 23204 19295 23256 19304
rect 23204 19261 23213 19295
rect 23213 19261 23247 19295
rect 23247 19261 23256 19295
rect 23204 19252 23256 19261
rect 25504 19295 25556 19304
rect 25504 19261 25513 19295
rect 25513 19261 25547 19295
rect 25547 19261 25556 19295
rect 25504 19252 25556 19261
rect 18236 19184 18288 19236
rect 18788 19184 18840 19236
rect 19524 19227 19576 19236
rect 19524 19193 19533 19227
rect 19533 19193 19567 19227
rect 19567 19193 19576 19227
rect 19524 19184 19576 19193
rect 19800 19184 19852 19236
rect 20260 19184 20312 19236
rect 18880 19116 18932 19168
rect 19156 19116 19208 19168
rect 19616 19116 19668 19168
rect 27620 19227 27672 19236
rect 27620 19193 27629 19227
rect 27629 19193 27663 19227
rect 27663 19193 27672 19227
rect 27620 19184 27672 19193
rect 20444 19116 20496 19168
rect 20904 19116 20956 19168
rect 21364 19116 21416 19168
rect 31024 19184 31076 19236
rect 35348 19252 35400 19304
rect 34244 19184 34296 19236
rect 28172 19116 28224 19168
rect 28724 19116 28776 19168
rect 30196 19159 30248 19168
rect 30196 19125 30205 19159
rect 30205 19125 30239 19159
rect 30239 19125 30248 19159
rect 30196 19116 30248 19125
rect 32404 19159 32456 19168
rect 32404 19125 32413 19159
rect 32413 19125 32447 19159
rect 32447 19125 32456 19159
rect 32404 19116 32456 19125
rect 34612 19116 34664 19168
rect 35624 19159 35676 19168
rect 35624 19125 35633 19159
rect 35633 19125 35667 19159
rect 35667 19125 35676 19159
rect 35624 19116 35676 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2044 18955 2096 18964
rect 2044 18921 2053 18955
rect 2053 18921 2087 18955
rect 2087 18921 2096 18955
rect 2044 18912 2096 18921
rect 3148 18912 3200 18964
rect 4712 18912 4764 18964
rect 3700 18844 3752 18896
rect 5908 18844 5960 18896
rect 1032 18776 1084 18828
rect 2688 18819 2740 18828
rect 2688 18785 2697 18819
rect 2697 18785 2731 18819
rect 2731 18785 2740 18819
rect 2688 18776 2740 18785
rect 5632 18776 5684 18828
rect 9588 18912 9640 18964
rect 13728 18912 13780 18964
rect 14096 18912 14148 18964
rect 16396 18912 16448 18964
rect 1124 18708 1176 18760
rect 2044 18751 2096 18760
rect 2044 18717 2053 18751
rect 2053 18717 2087 18751
rect 2087 18717 2096 18751
rect 2044 18708 2096 18717
rect 3240 18708 3292 18760
rect 4528 18708 4580 18760
rect 9680 18844 9732 18896
rect 8208 18819 8260 18828
rect 8208 18785 8217 18819
rect 8217 18785 8251 18819
rect 8251 18785 8260 18819
rect 8208 18776 8260 18785
rect 9036 18776 9088 18828
rect 10600 18819 10652 18828
rect 10600 18785 10609 18819
rect 10609 18785 10643 18819
rect 10643 18785 10652 18819
rect 10600 18776 10652 18785
rect 13544 18844 13596 18896
rect 11520 18776 11572 18828
rect 14280 18776 14332 18828
rect 15936 18819 15988 18828
rect 15936 18785 15945 18819
rect 15945 18785 15979 18819
rect 15979 18785 15988 18819
rect 15936 18776 15988 18785
rect 14372 18751 14424 18760
rect 4712 18640 4764 18692
rect 2688 18572 2740 18624
rect 3792 18572 3844 18624
rect 10416 18640 10468 18692
rect 10876 18640 10928 18692
rect 11060 18683 11112 18692
rect 11060 18649 11069 18683
rect 11069 18649 11103 18683
rect 11103 18649 11112 18683
rect 11060 18640 11112 18649
rect 9496 18572 9548 18624
rect 10508 18572 10560 18624
rect 13544 18640 13596 18692
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 17040 18844 17092 18896
rect 17868 18776 17920 18828
rect 12716 18572 12768 18624
rect 13176 18572 13228 18624
rect 14740 18572 14792 18624
rect 16672 18572 16724 18624
rect 17132 18640 17184 18692
rect 17500 18708 17552 18760
rect 17684 18708 17736 18760
rect 20260 18912 20312 18964
rect 21548 18955 21600 18964
rect 18144 18887 18196 18896
rect 18144 18853 18153 18887
rect 18153 18853 18187 18887
rect 18187 18853 18196 18887
rect 18144 18844 18196 18853
rect 18052 18776 18104 18828
rect 19524 18844 19576 18896
rect 19800 18844 19852 18896
rect 20076 18844 20128 18896
rect 20352 18844 20404 18896
rect 21548 18921 21557 18955
rect 21557 18921 21591 18955
rect 21591 18921 21600 18955
rect 21548 18912 21600 18921
rect 22560 18912 22612 18964
rect 23480 18912 23532 18964
rect 24308 18912 24360 18964
rect 24952 18955 25004 18964
rect 24952 18921 24961 18955
rect 24961 18921 24995 18955
rect 24995 18921 25004 18955
rect 24952 18912 25004 18921
rect 27252 18955 27304 18964
rect 27252 18921 27261 18955
rect 27261 18921 27295 18955
rect 27295 18921 27304 18955
rect 27252 18912 27304 18921
rect 27620 18912 27672 18964
rect 36268 18912 36320 18964
rect 21456 18844 21508 18896
rect 30104 18844 30156 18896
rect 35624 18844 35676 18896
rect 18052 18640 18104 18692
rect 19616 18708 19668 18760
rect 30564 18776 30616 18828
rect 20444 18708 20496 18760
rect 20812 18708 20864 18760
rect 21548 18708 21600 18760
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22376 18708 22428 18717
rect 22744 18708 22796 18760
rect 24768 18708 24820 18760
rect 30748 18708 30800 18760
rect 18788 18640 18840 18692
rect 19800 18640 19852 18692
rect 21640 18640 21692 18692
rect 22652 18640 22704 18692
rect 26976 18640 27028 18692
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 18512 18572 18564 18624
rect 20996 18572 21048 18624
rect 24492 18572 24544 18624
rect 26608 18615 26660 18624
rect 26608 18581 26617 18615
rect 26617 18581 26651 18615
rect 26651 18581 26660 18615
rect 30196 18640 30248 18692
rect 43996 18640 44048 18692
rect 33968 18615 34020 18624
rect 26608 18572 26660 18581
rect 33968 18581 33977 18615
rect 33977 18581 34011 18615
rect 34011 18581 34020 18615
rect 33968 18572 34020 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4160 18368 4212 18420
rect 9128 18368 9180 18420
rect 9220 18368 9272 18420
rect 11980 18368 12032 18420
rect 4988 18300 5040 18352
rect 5448 18300 5500 18352
rect 7840 18300 7892 18352
rect 14372 18368 14424 18420
rect 16028 18411 16080 18420
rect 16028 18377 16037 18411
rect 16037 18377 16071 18411
rect 16071 18377 16080 18411
rect 16028 18368 16080 18377
rect 17316 18368 17368 18420
rect 18236 18411 18288 18420
rect 18236 18377 18245 18411
rect 18245 18377 18279 18411
rect 18279 18377 18288 18411
rect 18236 18368 18288 18377
rect 18880 18368 18932 18420
rect 20812 18368 20864 18420
rect 21364 18368 21416 18420
rect 21456 18368 21508 18420
rect 22928 18411 22980 18420
rect 21732 18300 21784 18352
rect 22284 18343 22336 18352
rect 22284 18309 22293 18343
rect 22293 18309 22327 18343
rect 22327 18309 22336 18343
rect 22284 18300 22336 18309
rect 22928 18377 22937 18411
rect 22937 18377 22971 18411
rect 22971 18377 22980 18411
rect 22928 18368 22980 18377
rect 23572 18411 23624 18420
rect 23572 18377 23581 18411
rect 23581 18377 23615 18411
rect 23615 18377 23624 18411
rect 23572 18368 23624 18377
rect 24768 18411 24820 18420
rect 24768 18377 24777 18411
rect 24777 18377 24811 18411
rect 24811 18377 24820 18411
rect 24768 18368 24820 18377
rect 24952 18368 25004 18420
rect 27436 18368 27488 18420
rect 28080 18368 28132 18420
rect 29276 18411 29328 18420
rect 29276 18377 29285 18411
rect 29285 18377 29319 18411
rect 29319 18377 29328 18411
rect 29276 18368 29328 18377
rect 3976 18275 4028 18284
rect 3976 18241 3985 18275
rect 3985 18241 4019 18275
rect 4019 18241 4028 18275
rect 3976 18232 4028 18241
rect 4436 18275 4488 18284
rect 4436 18241 4445 18275
rect 4445 18241 4479 18275
rect 4479 18241 4488 18275
rect 4436 18232 4488 18241
rect 5632 18232 5684 18284
rect 6276 18232 6328 18284
rect 6920 18207 6972 18216
rect 2872 18096 2924 18148
rect 2596 18028 2648 18080
rect 3332 18028 3384 18080
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 11336 18232 11388 18284
rect 14096 18275 14148 18284
rect 14096 18241 14105 18275
rect 14105 18241 14139 18275
rect 14139 18241 14148 18275
rect 14096 18232 14148 18241
rect 16488 18232 16540 18284
rect 16672 18232 16724 18284
rect 17132 18275 17184 18284
rect 17132 18241 17141 18275
rect 17141 18241 17175 18275
rect 17175 18241 17184 18275
rect 17132 18232 17184 18241
rect 17408 18232 17460 18284
rect 9036 18207 9088 18216
rect 9036 18173 9045 18207
rect 9045 18173 9079 18207
rect 9079 18173 9088 18207
rect 9036 18164 9088 18173
rect 6368 18028 6420 18080
rect 8852 18028 8904 18080
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 15292 18164 15344 18216
rect 16856 18164 16908 18216
rect 17224 18207 17276 18216
rect 17224 18173 17233 18207
rect 17233 18173 17267 18207
rect 17267 18173 17276 18207
rect 17224 18164 17276 18173
rect 17316 18164 17368 18216
rect 18788 18232 18840 18284
rect 17868 18164 17920 18216
rect 19524 18207 19576 18216
rect 11152 18096 11204 18148
rect 11336 18096 11388 18148
rect 11428 18096 11480 18148
rect 12164 18096 12216 18148
rect 12992 18096 13044 18148
rect 11060 18028 11112 18080
rect 18512 18096 18564 18148
rect 19156 18139 19208 18148
rect 19156 18105 19165 18139
rect 19165 18105 19199 18139
rect 19199 18105 19208 18139
rect 19156 18096 19208 18105
rect 19524 18173 19533 18207
rect 19533 18173 19567 18207
rect 19567 18173 19576 18207
rect 19524 18164 19576 18173
rect 19708 18164 19760 18216
rect 20444 18207 20496 18216
rect 20444 18173 20453 18207
rect 20453 18173 20487 18207
rect 20487 18173 20496 18207
rect 20444 18164 20496 18173
rect 20996 18275 21048 18284
rect 20996 18241 21005 18275
rect 21005 18241 21039 18275
rect 21039 18241 21048 18275
rect 20996 18232 21048 18241
rect 23020 18232 23072 18284
rect 24032 18232 24084 18284
rect 24768 18232 24820 18284
rect 25320 18275 25372 18284
rect 25320 18241 25329 18275
rect 25329 18241 25363 18275
rect 25363 18241 25372 18275
rect 25320 18232 25372 18241
rect 27252 18232 27304 18284
rect 28172 18275 28224 18284
rect 28172 18241 28181 18275
rect 28181 18241 28215 18275
rect 28215 18241 28224 18275
rect 28172 18232 28224 18241
rect 21364 18164 21416 18216
rect 23296 18164 23348 18216
rect 26332 18207 26384 18216
rect 26332 18173 26341 18207
rect 26341 18173 26375 18207
rect 26375 18173 26384 18207
rect 26332 18164 26384 18173
rect 29000 18300 29052 18352
rect 30288 18300 30340 18352
rect 29920 18232 29972 18284
rect 28356 18164 28408 18216
rect 29184 18164 29236 18216
rect 19984 18096 20036 18148
rect 20536 18096 20588 18148
rect 16488 18028 16540 18080
rect 16948 18028 17000 18080
rect 18144 18028 18196 18080
rect 19524 18028 19576 18080
rect 21916 18028 21968 18080
rect 24032 18096 24084 18148
rect 31760 18096 31812 18148
rect 25320 18028 25372 18080
rect 27068 18071 27120 18080
rect 27068 18037 27077 18071
rect 27077 18037 27111 18071
rect 27111 18037 27120 18071
rect 27068 18028 27120 18037
rect 27252 18028 27304 18080
rect 30840 18028 30892 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 1768 17824 1820 17876
rect 6736 17824 6788 17876
rect 9864 17824 9916 17876
rect 11060 17824 11112 17876
rect 11244 17824 11296 17876
rect 12072 17824 12124 17876
rect 2228 17688 2280 17740
rect 6184 17756 6236 17808
rect 6644 17756 6696 17808
rect 13176 17824 13228 17876
rect 13360 17824 13412 17876
rect 14464 17824 14516 17876
rect 14740 17824 14792 17876
rect 16948 17824 17000 17876
rect 17132 17867 17184 17876
rect 17132 17833 17141 17867
rect 17141 17833 17175 17867
rect 17175 17833 17184 17867
rect 17132 17824 17184 17833
rect 17408 17824 17460 17876
rect 18420 17824 18472 17876
rect 19156 17824 19208 17876
rect 19248 17824 19300 17876
rect 19524 17824 19576 17876
rect 20444 17824 20496 17876
rect 20904 17867 20956 17876
rect 20904 17833 20913 17867
rect 20913 17833 20947 17867
rect 20947 17833 20956 17867
rect 20904 17824 20956 17833
rect 22192 17824 22244 17876
rect 19800 17756 19852 17808
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 1676 17663 1728 17672
rect 1676 17629 1685 17663
rect 1685 17629 1719 17663
rect 1719 17629 1728 17663
rect 1676 17620 1728 17629
rect 2872 17620 2924 17672
rect 3700 17688 3752 17740
rect 4068 17663 4120 17672
rect 4068 17629 4077 17663
rect 4077 17629 4111 17663
rect 4111 17629 4120 17663
rect 4620 17688 4672 17740
rect 5816 17688 5868 17740
rect 6736 17688 6788 17740
rect 7104 17688 7156 17740
rect 10508 17688 10560 17740
rect 12164 17688 12216 17740
rect 12440 17731 12492 17740
rect 12440 17697 12449 17731
rect 12449 17697 12483 17731
rect 12483 17697 12492 17731
rect 12440 17688 12492 17697
rect 13636 17688 13688 17740
rect 14096 17731 14148 17740
rect 14096 17697 14105 17731
rect 14105 17697 14139 17731
rect 14139 17697 14148 17731
rect 14096 17688 14148 17697
rect 16120 17731 16172 17740
rect 16120 17697 16129 17731
rect 16129 17697 16163 17731
rect 16163 17697 16172 17731
rect 16120 17688 16172 17697
rect 17224 17688 17276 17740
rect 17868 17688 17920 17740
rect 4068 17620 4120 17629
rect 5448 17620 5500 17672
rect 5540 17620 5592 17672
rect 6184 17620 6236 17672
rect 6460 17620 6512 17672
rect 10876 17620 10928 17672
rect 3056 17552 3108 17604
rect 3332 17552 3384 17604
rect 1860 17527 1912 17536
rect 1860 17493 1869 17527
rect 1869 17493 1903 17527
rect 1903 17493 1912 17527
rect 1860 17484 1912 17493
rect 3700 17484 3752 17536
rect 4804 17484 4856 17536
rect 5080 17552 5132 17604
rect 7104 17552 7156 17604
rect 7932 17552 7984 17604
rect 11428 17552 11480 17604
rect 12348 17552 12400 17604
rect 13360 17552 13412 17604
rect 13912 17620 13964 17672
rect 15660 17620 15712 17672
rect 15844 17620 15896 17672
rect 17316 17620 17368 17672
rect 17408 17620 17460 17672
rect 17500 17620 17552 17672
rect 18328 17620 18380 17672
rect 9772 17484 9824 17536
rect 17224 17552 17276 17604
rect 18696 17688 18748 17740
rect 18880 17688 18932 17740
rect 19524 17688 19576 17740
rect 22652 17756 22704 17808
rect 25688 17824 25740 17876
rect 26056 17867 26108 17876
rect 26056 17833 26065 17867
rect 26065 17833 26099 17867
rect 26099 17833 26108 17867
rect 26056 17824 26108 17833
rect 27896 17824 27948 17876
rect 28264 17867 28316 17876
rect 28264 17833 28273 17867
rect 28273 17833 28307 17867
rect 28307 17833 28316 17867
rect 28264 17824 28316 17833
rect 21088 17688 21140 17740
rect 19800 17620 19852 17672
rect 19984 17620 20036 17672
rect 18512 17595 18564 17604
rect 18512 17561 18539 17595
rect 18539 17561 18564 17595
rect 18512 17552 18564 17561
rect 16212 17527 16264 17536
rect 16212 17493 16221 17527
rect 16221 17493 16255 17527
rect 16255 17493 16264 17527
rect 16212 17484 16264 17493
rect 17316 17484 17368 17536
rect 17500 17527 17552 17536
rect 17500 17493 17509 17527
rect 17509 17493 17543 17527
rect 17543 17493 17552 17527
rect 17500 17484 17552 17493
rect 17868 17484 17920 17536
rect 17960 17484 18012 17536
rect 18052 17484 18104 17536
rect 18788 17552 18840 17604
rect 18972 17484 19024 17536
rect 19156 17484 19208 17536
rect 21364 17620 21416 17672
rect 22928 17688 22980 17740
rect 25136 17688 25188 17740
rect 21732 17552 21784 17604
rect 20260 17484 20312 17536
rect 20536 17484 20588 17536
rect 20996 17484 21048 17536
rect 21364 17484 21416 17536
rect 27068 17620 27120 17672
rect 27252 17620 27304 17672
rect 23020 17552 23072 17604
rect 23204 17484 23256 17536
rect 23572 17484 23624 17536
rect 24952 17527 25004 17536
rect 24952 17493 24961 17527
rect 24961 17493 24995 17527
rect 24995 17493 25004 17527
rect 24952 17484 25004 17493
rect 29184 17484 29236 17536
rect 29920 17484 29972 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 2780 17280 2832 17332
rect 3700 17280 3752 17332
rect 5632 17280 5684 17332
rect 5724 17280 5776 17332
rect 5908 17280 5960 17332
rect 10600 17280 10652 17332
rect 3884 17212 3936 17264
rect 4160 17212 4212 17264
rect 4804 17212 4856 17264
rect 10692 17212 10744 17264
rect 12256 17280 12308 17332
rect 17500 17280 17552 17332
rect 18604 17280 18656 17332
rect 22284 17280 22336 17332
rect 24032 17280 24084 17332
rect 28632 17280 28684 17332
rect 41604 17280 41656 17332
rect 11796 17212 11848 17264
rect 12348 17212 12400 17264
rect 13176 17255 13228 17264
rect 13176 17221 13185 17255
rect 13185 17221 13219 17255
rect 13219 17221 13228 17255
rect 13176 17212 13228 17221
rect 14188 17212 14240 17264
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 2320 17144 2372 17196
rect 2596 17187 2648 17196
rect 2596 17153 2605 17187
rect 2605 17153 2639 17187
rect 2639 17153 2648 17187
rect 2596 17144 2648 17153
rect 4436 17187 4488 17196
rect 4436 17153 4445 17187
rect 4445 17153 4479 17187
rect 4479 17153 4488 17187
rect 4436 17144 4488 17153
rect 756 17076 808 17128
rect 3976 17076 4028 17128
rect 6092 17144 6144 17196
rect 7104 17187 7156 17196
rect 7104 17153 7113 17187
rect 7113 17153 7147 17187
rect 7147 17153 7156 17187
rect 7104 17144 7156 17153
rect 7196 17144 7248 17196
rect 8484 17144 8536 17196
rect 8852 17144 8904 17196
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 9128 17076 9180 17128
rect 9864 17076 9916 17128
rect 13820 17076 13872 17128
rect 2136 17051 2188 17060
rect 2136 17017 2145 17051
rect 2145 17017 2179 17051
rect 2179 17017 2188 17051
rect 2136 17008 2188 17017
rect 12440 17008 12492 17060
rect 12532 17008 12584 17060
rect 15292 17076 15344 17128
rect 17960 17212 18012 17264
rect 18788 17212 18840 17264
rect 16672 17187 16724 17196
rect 16672 17153 16681 17187
rect 16681 17153 16715 17187
rect 16715 17153 16724 17187
rect 16672 17144 16724 17153
rect 16764 17144 16816 17196
rect 17224 17144 17276 17196
rect 18512 17144 18564 17196
rect 19984 17212 20036 17264
rect 20444 17212 20496 17264
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 21732 17144 21784 17196
rect 18788 17076 18840 17128
rect 19616 17076 19668 17128
rect 19800 17076 19852 17128
rect 20352 17076 20404 17128
rect 20536 17076 20588 17128
rect 22560 17144 22612 17196
rect 23480 17144 23532 17196
rect 29000 17212 29052 17264
rect 43904 17212 43956 17264
rect 27896 17144 27948 17196
rect 29644 17144 29696 17196
rect 23204 17076 23256 17128
rect 18328 17008 18380 17060
rect 480 16940 532 16992
rect 756 16940 808 16992
rect 3332 16940 3384 16992
rect 5724 16940 5776 16992
rect 5908 16940 5960 16992
rect 6000 16940 6052 16992
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 6736 16940 6788 16992
rect 10416 16940 10468 16992
rect 10600 16940 10652 16992
rect 15292 16940 15344 16992
rect 16396 16940 16448 16992
rect 16672 16940 16724 16992
rect 18512 16940 18564 16992
rect 18972 16940 19024 16992
rect 19340 16983 19392 16992
rect 19340 16949 19349 16983
rect 19349 16949 19383 16983
rect 19383 16949 19392 16983
rect 19340 16940 19392 16949
rect 21180 17008 21232 17060
rect 23388 17008 23440 17060
rect 24124 17076 24176 17128
rect 24768 17076 24820 17128
rect 29276 17076 29328 17128
rect 30380 17076 30432 17128
rect 20996 16940 21048 16992
rect 22192 16940 22244 16992
rect 22652 16940 22704 16992
rect 22928 16940 22980 16992
rect 23020 16940 23072 16992
rect 26056 17008 26108 17060
rect 24032 16983 24084 16992
rect 24032 16949 24041 16983
rect 24041 16949 24075 16983
rect 24075 16949 24084 16983
rect 24032 16940 24084 16949
rect 25412 16940 25464 16992
rect 26976 16983 27028 16992
rect 26976 16949 26985 16983
rect 26985 16949 27019 16983
rect 27019 16949 27028 16983
rect 26976 16940 27028 16949
rect 28908 16940 28960 16992
rect 29092 16940 29144 16992
rect 37924 16940 37976 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1768 16779 1820 16788
rect 1768 16745 1777 16779
rect 1777 16745 1811 16779
rect 1811 16745 1820 16779
rect 1768 16736 1820 16745
rect 1400 16600 1452 16652
rect 2872 16736 2924 16788
rect 4712 16600 4764 16652
rect 1584 16532 1636 16584
rect 3976 16532 4028 16584
rect 6736 16736 6788 16788
rect 7104 16736 7156 16788
rect 7196 16736 7248 16788
rect 8484 16736 8536 16788
rect 9128 16736 9180 16788
rect 8208 16668 8260 16720
rect 10140 16668 10192 16720
rect 10876 16668 10928 16720
rect 9312 16600 9364 16652
rect 9772 16643 9824 16652
rect 9772 16609 9781 16643
rect 9781 16609 9815 16643
rect 9815 16609 9824 16643
rect 9772 16600 9824 16609
rect 13636 16736 13688 16788
rect 14372 16736 14424 16788
rect 11520 16600 11572 16652
rect 6828 16532 6880 16584
rect 7472 16532 7524 16584
rect 12072 16575 12124 16584
rect 12072 16541 12081 16575
rect 12081 16541 12115 16575
rect 12115 16541 12124 16575
rect 12072 16532 12124 16541
rect 12440 16600 12492 16652
rect 16672 16736 16724 16788
rect 17684 16736 17736 16788
rect 18236 16736 18288 16788
rect 18788 16736 18840 16788
rect 19340 16736 19392 16788
rect 19708 16736 19760 16788
rect 20168 16736 20220 16788
rect 20904 16736 20956 16788
rect 23204 16736 23256 16788
rect 25872 16779 25924 16788
rect 13176 16600 13228 16652
rect 12992 16532 13044 16584
rect 16396 16600 16448 16652
rect 16672 16600 16724 16652
rect 17592 16600 17644 16652
rect 18144 16643 18196 16652
rect 18144 16609 18153 16643
rect 18153 16609 18187 16643
rect 18187 16609 18196 16643
rect 18144 16600 18196 16609
rect 19156 16668 19208 16720
rect 22468 16668 22520 16720
rect 24676 16668 24728 16720
rect 25504 16668 25556 16720
rect 25872 16745 25881 16779
rect 25881 16745 25915 16779
rect 25915 16745 25924 16779
rect 25872 16736 25924 16745
rect 27620 16736 27672 16788
rect 28356 16736 28408 16788
rect 27068 16711 27120 16720
rect 27068 16677 27077 16711
rect 27077 16677 27111 16711
rect 27111 16677 27120 16711
rect 27068 16668 27120 16677
rect 29552 16711 29604 16720
rect 29552 16677 29561 16711
rect 29561 16677 29595 16711
rect 29595 16677 29604 16711
rect 29552 16668 29604 16677
rect 19616 16643 19668 16652
rect 14740 16532 14792 16584
rect 14924 16575 14976 16584
rect 14924 16541 14958 16575
rect 14958 16541 14976 16575
rect 14924 16532 14976 16541
rect 16488 16532 16540 16584
rect 18328 16532 18380 16584
rect 19616 16609 19625 16643
rect 19625 16609 19659 16643
rect 19659 16609 19668 16643
rect 19616 16600 19668 16609
rect 20168 16600 20220 16652
rect 21272 16600 21324 16652
rect 21548 16643 21600 16652
rect 21548 16609 21557 16643
rect 21557 16609 21591 16643
rect 21591 16609 21600 16643
rect 21548 16600 21600 16609
rect 22100 16600 22152 16652
rect 22560 16600 22612 16652
rect 22928 16600 22980 16652
rect 25044 16600 25096 16652
rect 3332 16464 3384 16516
rect 5448 16464 5500 16516
rect 5632 16464 5684 16516
rect 10232 16464 10284 16516
rect 11612 16464 11664 16516
rect 15476 16464 15528 16516
rect 15844 16464 15896 16516
rect 3792 16396 3844 16448
rect 7380 16396 7432 16448
rect 8208 16396 8260 16448
rect 8852 16396 8904 16448
rect 13176 16439 13228 16448
rect 13176 16405 13185 16439
rect 13185 16405 13219 16439
rect 13219 16405 13228 16439
rect 13176 16396 13228 16405
rect 13820 16396 13872 16448
rect 17868 16464 17920 16516
rect 19340 16464 19392 16516
rect 19984 16532 20036 16584
rect 20260 16532 20312 16584
rect 21180 16532 21232 16584
rect 23296 16575 23348 16584
rect 23296 16541 23305 16575
rect 23305 16541 23339 16575
rect 23339 16541 23348 16575
rect 23296 16532 23348 16541
rect 20628 16507 20680 16516
rect 20628 16473 20637 16507
rect 20637 16473 20671 16507
rect 20671 16473 20680 16507
rect 20628 16464 20680 16473
rect 22008 16507 22060 16516
rect 22008 16473 22017 16507
rect 22017 16473 22051 16507
rect 22051 16473 22060 16507
rect 22008 16464 22060 16473
rect 25228 16507 25280 16516
rect 16120 16396 16172 16448
rect 18604 16396 18656 16448
rect 18696 16396 18748 16448
rect 20260 16396 20312 16448
rect 21272 16396 21324 16448
rect 23296 16396 23348 16448
rect 25228 16473 25237 16507
rect 25237 16473 25271 16507
rect 25271 16473 25280 16507
rect 25228 16464 25280 16473
rect 26424 16439 26476 16448
rect 26424 16405 26433 16439
rect 26433 16405 26467 16439
rect 26467 16405 26476 16439
rect 26424 16396 26476 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 1676 16235 1728 16244
rect 1676 16201 1685 16235
rect 1685 16201 1719 16235
rect 1719 16201 1728 16235
rect 1676 16192 1728 16201
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 848 16124 900 16176
rect 4068 16192 4120 16244
rect 5264 16124 5316 16176
rect 7932 16124 7984 16176
rect 1308 16056 1360 16108
rect 2596 16099 2648 16108
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 2596 16065 2605 16099
rect 2605 16065 2639 16099
rect 2639 16065 2648 16099
rect 2596 16056 2648 16065
rect 4528 16056 4580 16108
rect 5172 16056 5224 16108
rect 6460 16099 6512 16108
rect 6460 16065 6469 16099
rect 6469 16065 6503 16099
rect 6503 16065 6512 16099
rect 6460 16056 6512 16065
rect 6368 15920 6420 15972
rect 8576 16056 8628 16108
rect 9404 16192 9456 16244
rect 11336 16192 11388 16244
rect 11612 16235 11664 16244
rect 11612 16201 11621 16235
rect 11621 16201 11655 16235
rect 11655 16201 11664 16235
rect 11612 16192 11664 16201
rect 8944 16124 8996 16176
rect 9128 16099 9180 16108
rect 9128 16065 9137 16099
rect 9137 16065 9171 16099
rect 9171 16065 9180 16099
rect 9128 16056 9180 16065
rect 16672 16235 16724 16244
rect 16672 16201 16681 16235
rect 16681 16201 16715 16235
rect 16715 16201 16724 16235
rect 16672 16192 16724 16201
rect 16948 16192 17000 16244
rect 20904 16192 20956 16244
rect 21824 16235 21876 16244
rect 21824 16201 21833 16235
rect 21833 16201 21867 16235
rect 21867 16201 21876 16235
rect 21824 16192 21876 16201
rect 13084 16124 13136 16176
rect 14096 16124 14148 16176
rect 17776 16167 17828 16176
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 14832 16056 14884 16108
rect 17776 16133 17794 16167
rect 17794 16133 17828 16167
rect 17776 16124 17828 16133
rect 15844 16056 15896 16108
rect 16120 16056 16172 16108
rect 17960 16056 18012 16108
rect 19248 16124 19300 16176
rect 20076 16124 20128 16176
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 19892 16099 19944 16108
rect 19892 16065 19901 16099
rect 19901 16065 19935 16099
rect 19935 16065 19944 16099
rect 19892 16056 19944 16065
rect 19984 16099 20036 16108
rect 19984 16065 19993 16099
rect 19993 16065 20027 16099
rect 20027 16065 20036 16099
rect 19984 16056 20036 16065
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 15476 16031 15528 16040
rect 3884 15852 3936 15904
rect 6920 15852 6972 15904
rect 7380 15852 7432 15904
rect 10140 15852 10192 15904
rect 15476 15997 15485 16031
rect 15485 15997 15519 16031
rect 15519 15997 15528 16031
rect 15476 15988 15528 15997
rect 18604 16031 18656 16040
rect 18604 15997 18613 16031
rect 18613 15997 18647 16031
rect 18647 15997 18656 16031
rect 18604 15988 18656 15997
rect 19064 15988 19116 16040
rect 21456 16124 21508 16176
rect 23480 16192 23532 16244
rect 24400 16192 24452 16244
rect 25044 16235 25096 16244
rect 25044 16201 25053 16235
rect 25053 16201 25087 16235
rect 25087 16201 25096 16235
rect 25044 16192 25096 16201
rect 25320 16192 25372 16244
rect 26792 16192 26844 16244
rect 27620 16235 27672 16244
rect 27620 16201 27629 16235
rect 27629 16201 27663 16235
rect 27663 16201 27672 16235
rect 27620 16192 27672 16201
rect 22836 16124 22888 16176
rect 23204 16167 23256 16176
rect 23204 16133 23213 16167
rect 23213 16133 23247 16167
rect 23247 16133 23256 16167
rect 23204 16124 23256 16133
rect 23296 16124 23348 16176
rect 20536 16056 20588 16108
rect 20996 15988 21048 16040
rect 21548 16056 21600 16108
rect 26332 16124 26384 16176
rect 24952 16056 25004 16108
rect 26976 16099 27028 16108
rect 26976 16065 26985 16099
rect 26985 16065 27019 16099
rect 27019 16065 27028 16099
rect 26976 16056 27028 16065
rect 16488 15852 16540 15904
rect 19156 15920 19208 15972
rect 19432 15920 19484 15972
rect 17776 15852 17828 15904
rect 18420 15852 18472 15904
rect 20536 15852 20588 15904
rect 20720 15920 20772 15972
rect 22560 15920 22612 15972
rect 21180 15852 21232 15904
rect 22744 16031 22796 16040
rect 22744 15997 22753 16031
rect 22753 15997 22787 16031
rect 22787 15997 22796 16031
rect 22744 15988 22796 15997
rect 24032 15988 24084 16040
rect 23756 15920 23808 15972
rect 24308 15963 24360 15972
rect 24308 15929 24317 15963
rect 24317 15929 24351 15963
rect 24351 15929 24360 15963
rect 24308 15920 24360 15929
rect 24860 15920 24912 15972
rect 24676 15852 24728 15904
rect 26608 15852 26660 15904
rect 28632 15895 28684 15904
rect 28632 15861 28641 15895
rect 28641 15861 28675 15895
rect 28675 15861 28684 15895
rect 28632 15852 28684 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1768 15691 1820 15700
rect 1768 15657 1777 15691
rect 1777 15657 1811 15691
rect 1811 15657 1820 15691
rect 1768 15648 1820 15657
rect 2136 15648 2188 15700
rect 3884 15648 3936 15700
rect 756 15580 808 15632
rect 1400 15512 1452 15564
rect 4988 15580 5040 15632
rect 8760 15580 8812 15632
rect 4620 15555 4672 15564
rect 4620 15521 4629 15555
rect 4629 15521 4663 15555
rect 4663 15521 4672 15555
rect 4620 15512 4672 15521
rect 13636 15648 13688 15700
rect 14464 15648 14516 15700
rect 14832 15648 14884 15700
rect 10876 15555 10928 15564
rect 10876 15521 10885 15555
rect 10885 15521 10919 15555
rect 10919 15521 10928 15555
rect 10876 15512 10928 15521
rect 11612 15512 11664 15564
rect 13728 15512 13780 15564
rect 18144 15648 18196 15700
rect 17224 15580 17276 15632
rect 19248 15623 19300 15632
rect 19248 15589 19257 15623
rect 19257 15589 19291 15623
rect 19291 15589 19300 15623
rect 19248 15580 19300 15589
rect 20536 15648 20588 15700
rect 21548 15691 21600 15700
rect 20904 15580 20956 15632
rect 21548 15657 21557 15691
rect 21557 15657 21591 15691
rect 21591 15657 21600 15691
rect 21548 15648 21600 15657
rect 24952 15648 25004 15700
rect 26148 15648 26200 15700
rect 26332 15691 26384 15700
rect 26332 15657 26341 15691
rect 26341 15657 26375 15691
rect 26375 15657 26384 15691
rect 26332 15648 26384 15657
rect 26792 15691 26844 15700
rect 26792 15657 26801 15691
rect 26801 15657 26835 15691
rect 26835 15657 26844 15691
rect 26792 15648 26844 15657
rect 26976 15648 27028 15700
rect 29368 15648 29420 15700
rect 29644 15648 29696 15700
rect 21640 15580 21692 15632
rect 22284 15623 22336 15632
rect 22284 15589 22293 15623
rect 22293 15589 22327 15623
rect 22327 15589 22336 15623
rect 22284 15580 22336 15589
rect 22928 15623 22980 15632
rect 22928 15589 22937 15623
rect 22937 15589 22971 15623
rect 22971 15589 22980 15623
rect 22928 15580 22980 15589
rect 24216 15580 24268 15632
rect 24584 15580 24636 15632
rect 25872 15580 25924 15632
rect 26056 15580 26108 15632
rect 27436 15580 27488 15632
rect 19156 15512 19208 15564
rect 19616 15555 19668 15564
rect 19616 15521 19625 15555
rect 19625 15521 19659 15555
rect 19659 15521 19668 15555
rect 19616 15512 19668 15521
rect 20168 15512 20220 15564
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 3240 15444 3292 15496
rect 3332 15376 3384 15428
rect 4528 15444 4580 15496
rect 6644 15444 6696 15496
rect 6828 15444 6880 15496
rect 7196 15487 7248 15496
rect 7196 15453 7230 15487
rect 7230 15453 7248 15487
rect 7196 15444 7248 15453
rect 11152 15444 11204 15496
rect 12348 15444 12400 15496
rect 13820 15444 13872 15496
rect 14740 15444 14792 15496
rect 16672 15444 16724 15496
rect 17960 15444 18012 15496
rect 6552 15376 6604 15428
rect 11428 15376 11480 15428
rect 2136 15308 2188 15360
rect 5632 15308 5684 15360
rect 9956 15308 10008 15360
rect 15476 15376 15528 15428
rect 15752 15376 15804 15428
rect 19524 15444 19576 15496
rect 20076 15444 20128 15496
rect 20720 15512 20772 15564
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 22376 15512 22428 15564
rect 21548 15444 21600 15496
rect 22744 15444 22796 15496
rect 26332 15512 26384 15564
rect 26424 15512 26476 15564
rect 23848 15487 23900 15496
rect 16580 15308 16632 15360
rect 17224 15308 17276 15360
rect 17408 15351 17460 15360
rect 17408 15317 17417 15351
rect 17417 15317 17451 15351
rect 17451 15317 17460 15351
rect 17408 15308 17460 15317
rect 17868 15308 17920 15360
rect 19984 15376 20036 15428
rect 20628 15419 20680 15428
rect 18328 15308 18380 15360
rect 20168 15351 20220 15360
rect 20168 15317 20177 15351
rect 20177 15317 20211 15351
rect 20211 15317 20220 15351
rect 20628 15385 20637 15419
rect 20637 15385 20671 15419
rect 20671 15385 20680 15419
rect 20628 15376 20680 15385
rect 21272 15376 21324 15428
rect 22008 15419 22060 15428
rect 22008 15385 22017 15419
rect 22017 15385 22051 15419
rect 22051 15385 22060 15419
rect 22008 15376 22060 15385
rect 23296 15376 23348 15428
rect 23848 15453 23857 15487
rect 23857 15453 23891 15487
rect 23891 15453 23900 15487
rect 23848 15444 23900 15453
rect 24400 15444 24452 15496
rect 29368 15444 29420 15496
rect 25688 15376 25740 15428
rect 20168 15308 20220 15317
rect 27436 15308 27488 15360
rect 27528 15308 27580 15360
rect 28632 15308 28684 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2136 14968 2188 15020
rect 8484 15104 8536 15156
rect 8852 15104 8904 15156
rect 11244 15104 11296 15156
rect 13360 15104 13412 15156
rect 15292 15104 15344 15156
rect 18604 15104 18656 15156
rect 18696 15104 18748 15156
rect 4528 14968 4580 15020
rect 8208 15036 8260 15088
rect 2412 14943 2464 14952
rect 2412 14909 2421 14943
rect 2421 14909 2455 14943
rect 2455 14909 2464 14943
rect 2412 14900 2464 14909
rect 756 14832 808 14884
rect 5632 14900 5684 14952
rect 7104 14968 7156 15020
rect 7564 14968 7616 15020
rect 7748 14968 7800 15020
rect 12256 15036 12308 15088
rect 12900 15036 12952 15088
rect 15016 15036 15068 15088
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 14556 14968 14608 15020
rect 15844 15011 15896 15020
rect 15844 14977 15853 15011
rect 15853 14977 15887 15011
rect 15887 14977 15896 15011
rect 15844 14968 15896 14977
rect 16672 15011 16724 15020
rect 8944 14943 8996 14952
rect 8944 14909 8953 14943
rect 8953 14909 8987 14943
rect 8987 14909 8996 14943
rect 8944 14900 8996 14909
rect 8024 14832 8076 14884
rect 11612 14875 11664 14884
rect 11612 14841 11621 14875
rect 11621 14841 11655 14875
rect 11655 14841 11664 14875
rect 11612 14832 11664 14841
rect 5816 14807 5868 14816
rect 5816 14773 5825 14807
rect 5825 14773 5859 14807
rect 5859 14773 5868 14807
rect 5816 14764 5868 14773
rect 5908 14764 5960 14816
rect 6736 14764 6788 14816
rect 7656 14764 7708 14816
rect 9496 14764 9548 14816
rect 15568 14900 15620 14952
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 16580 14900 16632 14952
rect 18052 14968 18104 15020
rect 18880 14968 18932 15020
rect 19616 14900 19668 14952
rect 19892 15036 19944 15088
rect 20536 15104 20588 15156
rect 20812 15104 20864 15156
rect 21180 15147 21232 15156
rect 21180 15113 21189 15147
rect 21189 15113 21223 15147
rect 21223 15113 21232 15147
rect 21180 15104 21232 15113
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 20168 14968 20220 15020
rect 22376 15104 22428 15156
rect 24676 15104 24728 15156
rect 25596 15104 25648 15156
rect 26332 15147 26384 15156
rect 26332 15113 26341 15147
rect 26341 15113 26375 15147
rect 26375 15113 26384 15147
rect 26332 15104 26384 15113
rect 26424 15104 26476 15156
rect 28264 15104 28316 15156
rect 28448 15104 28500 15156
rect 23204 15036 23256 15088
rect 25504 15036 25556 15088
rect 27252 15036 27304 15088
rect 20996 15011 21048 15020
rect 20996 14977 21005 15011
rect 21005 14977 21039 15011
rect 21039 14977 21048 15011
rect 20996 14968 21048 14977
rect 21272 15011 21324 15020
rect 21272 14977 21281 15011
rect 21281 14977 21315 15011
rect 21315 14977 21324 15011
rect 21272 14968 21324 14977
rect 18972 14832 19024 14884
rect 19432 14832 19484 14884
rect 20812 14900 20864 14952
rect 21916 14968 21968 15020
rect 22192 14968 22244 15020
rect 22744 14968 22796 15020
rect 25044 14968 25096 15020
rect 26424 14968 26476 15020
rect 26700 14968 26752 15020
rect 27712 14968 27764 15020
rect 28448 14968 28500 15020
rect 28816 14968 28868 15020
rect 22836 14900 22888 14952
rect 20444 14832 20496 14884
rect 21364 14832 21416 14884
rect 23296 14900 23348 14952
rect 23572 14900 23624 14952
rect 24400 14900 24452 14952
rect 24032 14875 24084 14884
rect 24032 14841 24041 14875
rect 24041 14841 24075 14875
rect 24075 14841 24084 14875
rect 24032 14832 24084 14841
rect 24676 14832 24728 14884
rect 14096 14764 14148 14816
rect 15108 14764 15160 14816
rect 16580 14764 16632 14816
rect 18420 14764 18472 14816
rect 19708 14764 19760 14816
rect 20996 14764 21048 14816
rect 22836 14764 22888 14816
rect 23296 14764 23348 14816
rect 23848 14807 23900 14816
rect 23848 14773 23857 14807
rect 23857 14773 23891 14807
rect 23891 14773 23900 14807
rect 23848 14764 23900 14773
rect 24584 14764 24636 14816
rect 24952 14832 25004 14884
rect 27436 14764 27488 14816
rect 27804 14764 27856 14816
rect 28264 14764 28316 14816
rect 28632 14807 28684 14816
rect 28632 14773 28641 14807
rect 28641 14773 28675 14807
rect 28675 14773 28684 14807
rect 28632 14764 28684 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 940 14560 992 14612
rect 3976 14560 4028 14612
rect 4068 14560 4120 14612
rect 8944 14560 8996 14612
rect 9864 14560 9916 14612
rect 12992 14560 13044 14612
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 13268 14560 13320 14612
rect 4344 14492 4396 14544
rect 3792 14424 3844 14476
rect 4804 14492 4856 14544
rect 6276 14492 6328 14544
rect 8300 14492 8352 14544
rect 11152 14492 11204 14544
rect 12624 14535 12676 14544
rect 12624 14501 12633 14535
rect 12633 14501 12667 14535
rect 12667 14501 12676 14535
rect 12624 14492 12676 14501
rect 12716 14492 12768 14544
rect 4712 14467 4764 14476
rect 4712 14433 4721 14467
rect 4721 14433 4755 14467
rect 4755 14433 4764 14467
rect 4712 14424 4764 14433
rect 6828 14424 6880 14476
rect 15660 14492 15712 14544
rect 17408 14535 17460 14544
rect 17408 14501 17417 14535
rect 17417 14501 17451 14535
rect 17451 14501 17460 14535
rect 17408 14492 17460 14501
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 3608 14356 3660 14408
rect 3700 14288 3752 14340
rect 4620 14356 4672 14408
rect 5439 14399 5491 14408
rect 5439 14365 5448 14399
rect 5448 14365 5482 14399
rect 5482 14365 5491 14399
rect 5439 14356 5491 14365
rect 6276 14356 6328 14408
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 11244 14399 11296 14408
rect 10784 14356 10836 14365
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 11520 14399 11572 14408
rect 11520 14365 11554 14399
rect 11554 14365 11572 14399
rect 11520 14356 11572 14365
rect 6184 14288 6236 14340
rect 6368 14288 6420 14340
rect 3240 14220 3292 14272
rect 3884 14220 3936 14272
rect 6460 14220 6512 14272
rect 7840 14288 7892 14340
rect 7932 14288 7984 14340
rect 8576 14288 8628 14340
rect 10048 14288 10100 14340
rect 11152 14288 11204 14340
rect 11980 14288 12032 14340
rect 8024 14220 8076 14272
rect 13912 14356 13964 14408
rect 14096 14399 14148 14408
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 19616 14560 19668 14612
rect 19984 14560 20036 14612
rect 20444 14560 20496 14612
rect 21732 14560 21784 14612
rect 22008 14560 22060 14612
rect 26056 14560 26108 14612
rect 26976 14560 27028 14612
rect 27436 14603 27488 14612
rect 27436 14569 27445 14603
rect 27445 14569 27479 14603
rect 27479 14569 27488 14603
rect 27436 14560 27488 14569
rect 27620 14560 27672 14612
rect 20076 14492 20128 14544
rect 20352 14535 20404 14544
rect 20352 14501 20361 14535
rect 20361 14501 20395 14535
rect 20395 14501 20404 14535
rect 20352 14492 20404 14501
rect 22192 14535 22244 14544
rect 22192 14501 22201 14535
rect 22201 14501 22235 14535
rect 22235 14501 22244 14535
rect 22192 14492 22244 14501
rect 22836 14492 22888 14544
rect 15568 14356 15620 14408
rect 16672 14356 16724 14408
rect 16764 14356 16816 14408
rect 18696 14399 18748 14408
rect 18696 14365 18705 14399
rect 18705 14365 18739 14399
rect 18739 14365 18748 14399
rect 18696 14356 18748 14365
rect 19248 14399 19300 14408
rect 19248 14365 19257 14399
rect 19257 14365 19291 14399
rect 19291 14365 19300 14399
rect 19248 14356 19300 14365
rect 19432 14356 19484 14408
rect 19708 14399 19760 14408
rect 19708 14365 19717 14399
rect 19717 14365 19751 14399
rect 19751 14365 19760 14399
rect 19708 14356 19760 14365
rect 20812 14399 20864 14408
rect 13360 14331 13412 14340
rect 13360 14297 13369 14331
rect 13369 14297 13403 14331
rect 13403 14297 13412 14331
rect 13360 14288 13412 14297
rect 13544 14331 13596 14340
rect 13544 14297 13553 14331
rect 13553 14297 13587 14331
rect 13587 14297 13596 14331
rect 13544 14288 13596 14297
rect 14004 14288 14056 14340
rect 16304 14331 16356 14340
rect 16304 14297 16338 14331
rect 16338 14297 16356 14331
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 21456 14399 21508 14408
rect 21456 14365 21465 14399
rect 21465 14365 21499 14399
rect 21499 14365 21508 14399
rect 21456 14356 21508 14365
rect 16304 14288 16356 14297
rect 13636 14220 13688 14272
rect 16580 14220 16632 14272
rect 18420 14220 18472 14272
rect 19248 14220 19300 14272
rect 20168 14220 20220 14272
rect 21088 14288 21140 14340
rect 21272 14331 21324 14340
rect 21272 14297 21281 14331
rect 21281 14297 21315 14331
rect 21315 14297 21324 14331
rect 21272 14288 21324 14297
rect 22376 14424 22428 14476
rect 23388 14492 23440 14544
rect 27068 14492 27120 14544
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 22468 14288 22520 14340
rect 23572 14424 23624 14476
rect 22100 14220 22152 14272
rect 24032 14356 24084 14408
rect 24676 14356 24728 14408
rect 24860 14356 24912 14408
rect 30012 14560 30064 14612
rect 24952 14288 25004 14340
rect 26792 14288 26844 14340
rect 26332 14263 26384 14272
rect 26332 14229 26341 14263
rect 26341 14229 26375 14263
rect 26375 14229 26384 14263
rect 26332 14220 26384 14229
rect 27896 14263 27948 14272
rect 27896 14229 27905 14263
rect 27905 14229 27939 14263
rect 27939 14229 27948 14263
rect 27896 14220 27948 14229
rect 30656 14263 30708 14272
rect 30656 14229 30665 14263
rect 30665 14229 30699 14263
rect 30699 14229 30708 14263
rect 30656 14220 30708 14229
rect 33508 14220 33560 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 388 14016 440 14068
rect 2688 14016 2740 14068
rect 7472 14016 7524 14068
rect 7932 14016 7984 14068
rect 8208 14016 8260 14068
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 3516 13880 3568 13932
rect 5632 13948 5684 14000
rect 4528 13880 4580 13932
rect 4988 13880 5040 13932
rect 5264 13880 5316 13932
rect 6276 13880 6328 13932
rect 6460 13948 6512 14000
rect 6828 13948 6880 14000
rect 8024 13948 8076 14000
rect 9312 13948 9364 14000
rect 6644 13923 6696 13932
rect 6644 13889 6678 13923
rect 6678 13889 6696 13923
rect 6644 13880 6696 13889
rect 2596 13812 2648 13864
rect 1584 13787 1636 13796
rect 1584 13753 1593 13787
rect 1593 13753 1627 13787
rect 1627 13753 1636 13787
rect 3608 13812 3660 13864
rect 3976 13855 4028 13864
rect 1584 13744 1636 13753
rect 2228 13719 2280 13728
rect 2228 13685 2237 13719
rect 2237 13685 2271 13719
rect 2271 13685 2280 13719
rect 2228 13676 2280 13685
rect 3240 13676 3292 13728
rect 3976 13821 3985 13855
rect 3985 13821 4019 13855
rect 4019 13821 4028 13855
rect 3976 13812 4028 13821
rect 7932 13744 7984 13796
rect 10508 13948 10560 14000
rect 11060 13948 11112 14000
rect 12256 14016 12308 14068
rect 18052 14016 18104 14068
rect 11980 13948 12032 14000
rect 14096 13948 14148 14000
rect 8576 13812 8628 13864
rect 9864 13812 9916 13864
rect 9128 13676 9180 13728
rect 9680 13744 9732 13796
rect 10416 13812 10468 13864
rect 10600 13812 10652 13864
rect 11244 13812 11296 13864
rect 11152 13744 11204 13796
rect 13820 13812 13872 13864
rect 14464 13880 14516 13932
rect 17040 13948 17092 14000
rect 19248 14016 19300 14068
rect 20352 14016 20404 14068
rect 14924 13923 14976 13932
rect 14924 13889 14958 13923
rect 14958 13889 14976 13923
rect 14924 13880 14976 13889
rect 15660 13880 15712 13932
rect 16672 13923 16724 13932
rect 14004 13855 14056 13864
rect 14004 13821 14013 13855
rect 14013 13821 14047 13855
rect 14047 13821 14056 13855
rect 14004 13812 14056 13821
rect 15752 13812 15804 13864
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 16672 13880 16724 13889
rect 18512 13948 18564 14000
rect 18052 13880 18104 13932
rect 18604 13923 18656 13932
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 14464 13744 14516 13796
rect 14648 13744 14700 13796
rect 18328 13812 18380 13864
rect 20076 13880 20128 13932
rect 20168 13880 20220 13932
rect 20536 13923 20588 13932
rect 20536 13889 20545 13923
rect 20545 13889 20579 13923
rect 20579 13889 20588 13923
rect 20536 13880 20588 13889
rect 20904 13880 20956 13932
rect 21088 13948 21140 14000
rect 23388 14016 23440 14068
rect 23756 14016 23808 14068
rect 22652 13923 22704 13932
rect 22652 13889 22683 13923
rect 22683 13889 22704 13923
rect 22652 13880 22704 13889
rect 18604 13744 18656 13796
rect 19432 13812 19484 13864
rect 18880 13744 18932 13796
rect 19524 13787 19576 13796
rect 19524 13753 19533 13787
rect 19533 13753 19567 13787
rect 19567 13753 19576 13787
rect 19524 13744 19576 13753
rect 19708 13744 19760 13796
rect 20260 13812 20312 13864
rect 21824 13812 21876 13864
rect 20168 13744 20220 13796
rect 22100 13744 22152 13796
rect 10876 13719 10928 13728
rect 10876 13685 10885 13719
rect 10885 13685 10919 13719
rect 10919 13685 10928 13719
rect 10876 13676 10928 13685
rect 12716 13676 12768 13728
rect 13544 13676 13596 13728
rect 18144 13676 18196 13728
rect 19064 13719 19116 13728
rect 19064 13685 19073 13719
rect 19073 13685 19107 13719
rect 19107 13685 19116 13719
rect 19064 13676 19116 13685
rect 19156 13676 19208 13728
rect 21916 13676 21968 13728
rect 22376 13676 22428 13728
rect 23940 13948 23992 14000
rect 24308 13923 24360 13932
rect 23388 13744 23440 13796
rect 23572 13744 23624 13796
rect 24308 13889 24317 13923
rect 24317 13889 24351 13923
rect 24351 13889 24360 13923
rect 24308 13880 24360 13889
rect 24676 14016 24728 14068
rect 28540 14016 28592 14068
rect 29276 14059 29328 14068
rect 29276 14025 29285 14059
rect 29285 14025 29319 14059
rect 29319 14025 29328 14059
rect 29276 14016 29328 14025
rect 30840 14059 30892 14068
rect 30840 14025 30849 14059
rect 30849 14025 30883 14059
rect 30883 14025 30892 14059
rect 30840 14016 30892 14025
rect 25320 13991 25372 14000
rect 25320 13957 25329 13991
rect 25329 13957 25363 13991
rect 25363 13957 25372 13991
rect 25320 13948 25372 13957
rect 25688 13948 25740 14000
rect 27528 13991 27580 14000
rect 27528 13957 27537 13991
rect 27537 13957 27571 13991
rect 27571 13957 27580 13991
rect 27528 13948 27580 13957
rect 28356 13948 28408 14000
rect 26148 13880 26200 13932
rect 26976 13855 27028 13864
rect 26976 13821 26985 13855
rect 26985 13821 27019 13855
rect 27019 13821 27028 13855
rect 26976 13812 27028 13821
rect 29000 13812 29052 13864
rect 28540 13744 28592 13796
rect 23664 13676 23716 13728
rect 25228 13676 25280 13728
rect 25964 13676 26016 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1768 13472 1820 13524
rect 848 13404 900 13456
rect 2044 13404 2096 13456
rect 2228 13404 2280 13456
rect 2320 13404 2372 13456
rect 2504 13404 2556 13456
rect 1492 13379 1544 13388
rect 1492 13345 1501 13379
rect 1501 13345 1535 13379
rect 1535 13345 1544 13379
rect 1492 13336 1544 13345
rect 3332 13404 3384 13456
rect 3884 13472 3936 13524
rect 5356 13472 5408 13524
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 6184 13472 6236 13524
rect 9680 13472 9732 13524
rect 1216 13268 1268 13320
rect 2044 13268 2096 13320
rect 1400 13243 1452 13252
rect 1400 13209 1409 13243
rect 1409 13209 1443 13243
rect 1443 13209 1452 13243
rect 1400 13200 1452 13209
rect 1492 13200 1544 13252
rect 2320 13200 2372 13252
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 3884 13379 3936 13388
rect 2780 13336 2832 13345
rect 3884 13345 3893 13379
rect 3893 13345 3927 13379
rect 3927 13345 3936 13379
rect 3884 13336 3936 13345
rect 2872 13311 2924 13320
rect 2872 13277 2881 13311
rect 2881 13277 2915 13311
rect 2915 13277 2924 13311
rect 2872 13268 2924 13277
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 3792 13268 3844 13277
rect 4160 13404 4212 13456
rect 6920 13404 6972 13456
rect 9496 13404 9548 13456
rect 8208 13336 8260 13388
rect 8852 13336 8904 13388
rect 14004 13472 14056 13524
rect 16304 13472 16356 13524
rect 19432 13472 19484 13524
rect 21272 13472 21324 13524
rect 22100 13515 22152 13524
rect 22100 13481 22109 13515
rect 22109 13481 22143 13515
rect 22143 13481 22152 13515
rect 22100 13472 22152 13481
rect 22376 13472 22428 13524
rect 22560 13472 22612 13524
rect 23848 13472 23900 13524
rect 25320 13472 25372 13524
rect 25504 13472 25556 13524
rect 27620 13472 27672 13524
rect 28264 13515 28316 13524
rect 28264 13481 28273 13515
rect 28273 13481 28307 13515
rect 28307 13481 28316 13515
rect 28264 13472 28316 13481
rect 28356 13472 28408 13524
rect 12256 13404 12308 13456
rect 17408 13404 17460 13456
rect 19524 13404 19576 13456
rect 12348 13336 12400 13388
rect 12716 13336 12768 13388
rect 17868 13336 17920 13388
rect 4068 13311 4120 13320
rect 4068 13277 4077 13311
rect 4077 13277 4111 13311
rect 4111 13277 4120 13311
rect 4068 13268 4120 13277
rect 4620 13268 4672 13320
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 11244 13311 11296 13320
rect 10784 13268 10836 13277
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 2504 13132 2556 13184
rect 6552 13200 6604 13252
rect 3792 13132 3844 13184
rect 8300 13132 8352 13184
rect 8576 13200 8628 13252
rect 10416 13200 10468 13252
rect 10876 13200 10928 13252
rect 8760 13132 8812 13184
rect 11704 13132 11756 13184
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 14096 13268 14148 13277
rect 14832 13268 14884 13320
rect 16672 13268 16724 13320
rect 18328 13268 18380 13320
rect 12716 13200 12768 13252
rect 15108 13200 15160 13252
rect 15200 13200 15252 13252
rect 18880 13336 18932 13388
rect 20628 13404 20680 13456
rect 19708 13379 19760 13388
rect 19708 13345 19717 13379
rect 19717 13345 19751 13379
rect 19751 13345 19760 13379
rect 21088 13379 21140 13388
rect 19708 13336 19760 13345
rect 21088 13345 21097 13379
rect 21097 13345 21131 13379
rect 21131 13345 21140 13379
rect 21088 13336 21140 13345
rect 18512 13268 18564 13320
rect 12992 13132 13044 13184
rect 13452 13132 13504 13184
rect 14280 13132 14332 13184
rect 16304 13132 16356 13184
rect 17224 13132 17276 13184
rect 17408 13132 17460 13184
rect 18144 13175 18196 13184
rect 18144 13141 18153 13175
rect 18153 13141 18187 13175
rect 18187 13141 18196 13175
rect 18880 13200 18932 13252
rect 20260 13268 20312 13320
rect 20628 13311 20680 13320
rect 20628 13277 20637 13311
rect 20637 13277 20671 13311
rect 20671 13277 20680 13311
rect 20628 13268 20680 13277
rect 21916 13404 21968 13456
rect 29000 13404 29052 13456
rect 21364 13336 21416 13388
rect 21456 13243 21508 13252
rect 21456 13209 21465 13243
rect 21465 13209 21499 13243
rect 21499 13209 21508 13243
rect 21456 13200 21508 13209
rect 21732 13200 21784 13252
rect 21916 13200 21968 13252
rect 18144 13132 18196 13141
rect 20076 13132 20128 13184
rect 20720 13132 20772 13184
rect 22560 13200 22612 13252
rect 23204 13268 23256 13320
rect 24768 13336 24820 13388
rect 26056 13336 26108 13388
rect 27896 13336 27948 13388
rect 28264 13336 28316 13388
rect 24492 13311 24544 13320
rect 24492 13277 24501 13311
rect 24501 13277 24535 13311
rect 24535 13277 24544 13311
rect 24492 13268 24544 13277
rect 26332 13268 26384 13320
rect 26148 13200 26200 13252
rect 26700 13200 26752 13252
rect 24308 13132 24360 13184
rect 27528 13132 27580 13184
rect 29644 13132 29696 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 2136 12928 2188 12980
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 6092 12928 6144 12980
rect 1492 12792 1544 12844
rect 2228 12860 2280 12912
rect 2872 12860 2924 12912
rect 3608 12903 3660 12912
rect 3608 12869 3617 12903
rect 3617 12869 3651 12903
rect 3651 12869 3660 12903
rect 3608 12860 3660 12869
rect 6184 12860 6236 12912
rect 6828 12860 6880 12912
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 2596 12792 2648 12844
rect 4068 12792 4120 12844
rect 4528 12792 4580 12844
rect 4712 12835 4764 12844
rect 4712 12801 4746 12835
rect 4746 12801 4764 12835
rect 6460 12835 6512 12844
rect 4712 12792 4764 12801
rect 6460 12801 6469 12835
rect 6469 12801 6503 12835
rect 6503 12801 6512 12835
rect 6460 12792 6512 12801
rect 6736 12835 6788 12844
rect 6736 12801 6770 12835
rect 6770 12801 6788 12835
rect 6736 12792 6788 12801
rect 9680 12928 9732 12980
rect 10324 12928 10376 12980
rect 15936 12928 15988 12980
rect 16212 12928 16264 12980
rect 16580 12928 16632 12980
rect 18328 12928 18380 12980
rect 18696 12928 18748 12980
rect 19156 12928 19208 12980
rect 19340 12928 19392 12980
rect 8484 12903 8536 12912
rect 8484 12869 8493 12903
rect 8493 12869 8527 12903
rect 8527 12869 8536 12903
rect 8484 12860 8536 12869
rect 7932 12792 7984 12844
rect 9956 12792 10008 12844
rect 11060 12792 11112 12844
rect 14096 12792 14148 12844
rect 14832 12835 14884 12844
rect 14832 12801 14841 12835
rect 14841 12801 14875 12835
rect 14875 12801 14884 12835
rect 15292 12835 15344 12844
rect 14832 12792 14884 12801
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 15476 12792 15528 12844
rect 17408 12792 17460 12844
rect 17500 12792 17552 12844
rect 17960 12792 18012 12844
rect 19248 12860 19300 12912
rect 19708 12860 19760 12912
rect 20720 12928 20772 12980
rect 23480 12928 23532 12980
rect 23664 12928 23716 12980
rect 24768 12928 24820 12980
rect 25964 12971 26016 12980
rect 19984 12860 20036 12912
rect 20628 12860 20680 12912
rect 21180 12903 21232 12912
rect 21180 12869 21189 12903
rect 21189 12869 21223 12903
rect 21223 12869 21232 12903
rect 21180 12860 21232 12869
rect 22560 12860 22612 12912
rect 24492 12860 24544 12912
rect 25964 12937 25973 12971
rect 25973 12937 26007 12971
rect 26007 12937 26016 12971
rect 25964 12928 26016 12937
rect 26148 12928 26200 12980
rect 28172 12971 28224 12980
rect 26516 12860 26568 12912
rect 27620 12860 27672 12912
rect 27804 12860 27856 12912
rect 28172 12937 28181 12971
rect 28181 12937 28215 12971
rect 28215 12937 28224 12971
rect 28172 12928 28224 12937
rect 29000 12928 29052 12980
rect 28908 12860 28960 12912
rect 29644 12928 29696 12980
rect 19064 12792 19116 12844
rect 22192 12835 22244 12844
rect 2964 12724 3016 12776
rect 3332 12767 3384 12776
rect 3332 12733 3341 12767
rect 3341 12733 3375 12767
rect 3375 12733 3384 12767
rect 3332 12724 3384 12733
rect 10600 12767 10652 12776
rect 1124 12656 1176 12708
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 2596 12588 2648 12640
rect 3700 12588 3752 12640
rect 3884 12588 3936 12640
rect 7748 12656 7800 12708
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 11152 12656 11204 12708
rect 11980 12656 12032 12708
rect 15016 12656 15068 12708
rect 16948 12656 17000 12708
rect 4712 12588 4764 12640
rect 5908 12588 5960 12640
rect 6368 12588 6420 12640
rect 6736 12588 6788 12640
rect 9220 12588 9272 12640
rect 11336 12588 11388 12640
rect 14648 12588 14700 12640
rect 16396 12588 16448 12640
rect 16580 12588 16632 12640
rect 16672 12588 16724 12640
rect 18328 12656 18380 12708
rect 19340 12724 19392 12776
rect 20444 12724 20496 12776
rect 21088 12656 21140 12708
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 23020 12792 23072 12844
rect 23664 12835 23716 12844
rect 23664 12801 23673 12835
rect 23673 12801 23707 12835
rect 23707 12801 23716 12835
rect 23664 12792 23716 12801
rect 23848 12835 23900 12844
rect 23848 12801 23857 12835
rect 23857 12801 23891 12835
rect 23891 12801 23900 12835
rect 23848 12792 23900 12801
rect 29828 12792 29880 12844
rect 22928 12724 22980 12776
rect 25228 12724 25280 12776
rect 23480 12699 23532 12708
rect 23480 12665 23489 12699
rect 23489 12665 23523 12699
rect 23523 12665 23532 12699
rect 23480 12656 23532 12665
rect 24308 12656 24360 12708
rect 28448 12656 28500 12708
rect 18604 12588 18656 12640
rect 18972 12588 19024 12640
rect 19432 12631 19484 12640
rect 19432 12597 19441 12631
rect 19441 12597 19475 12631
rect 19475 12597 19484 12631
rect 19432 12588 19484 12597
rect 19616 12631 19668 12640
rect 19616 12597 19625 12631
rect 19625 12597 19659 12631
rect 19659 12597 19668 12631
rect 19616 12588 19668 12597
rect 20260 12588 20312 12640
rect 20444 12631 20496 12640
rect 20444 12597 20453 12631
rect 20453 12597 20487 12631
rect 20487 12597 20496 12631
rect 20444 12588 20496 12597
rect 20720 12588 20772 12640
rect 24860 12588 24912 12640
rect 27068 12631 27120 12640
rect 27068 12597 27077 12631
rect 27077 12597 27111 12631
rect 27111 12597 27120 12631
rect 27068 12588 27120 12597
rect 27252 12588 27304 12640
rect 34612 12588 34664 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2596 12427 2648 12436
rect 2596 12393 2605 12427
rect 2605 12393 2639 12427
rect 2639 12393 2648 12427
rect 2596 12384 2648 12393
rect 5908 12384 5960 12436
rect 6276 12384 6328 12436
rect 6368 12384 6420 12436
rect 1860 12359 1912 12368
rect 1860 12325 1869 12359
rect 1869 12325 1903 12359
rect 1903 12325 1912 12359
rect 1860 12316 1912 12325
rect 2504 12291 2556 12300
rect 2504 12257 2513 12291
rect 2513 12257 2547 12291
rect 2547 12257 2556 12291
rect 2504 12248 2556 12257
rect 3700 12248 3752 12300
rect 4252 12248 4304 12300
rect 4528 12291 4580 12300
rect 4528 12257 4537 12291
rect 4537 12257 4571 12291
rect 4571 12257 4580 12291
rect 5264 12316 5316 12368
rect 5448 12316 5500 12368
rect 7196 12316 7248 12368
rect 7472 12316 7524 12368
rect 8116 12316 8168 12368
rect 8300 12316 8352 12368
rect 4528 12248 4580 12257
rect 1952 12180 2004 12232
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 2872 12180 2924 12232
rect 3424 12180 3476 12232
rect 3792 12180 3844 12232
rect 5540 12248 5592 12300
rect 8944 12291 8996 12300
rect 8944 12257 8953 12291
rect 8953 12257 8987 12291
rect 8987 12257 8996 12291
rect 8944 12248 8996 12257
rect 9128 12291 9180 12300
rect 9128 12257 9137 12291
rect 9137 12257 9171 12291
rect 9171 12257 9180 12291
rect 9128 12248 9180 12257
rect 12532 12384 12584 12436
rect 12716 12384 12768 12436
rect 10968 12316 11020 12368
rect 11888 12316 11940 12368
rect 15108 12384 15160 12436
rect 15292 12384 15344 12436
rect 15660 12384 15712 12436
rect 16396 12384 16448 12436
rect 16488 12359 16540 12368
rect 5816 12223 5868 12232
rect 5816 12189 5825 12223
rect 5825 12189 5859 12223
rect 5859 12189 5868 12223
rect 5816 12180 5868 12189
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 2504 12112 2556 12164
rect 3884 12112 3936 12164
rect 5080 12112 5132 12164
rect 5448 12112 5500 12164
rect 7472 12112 7524 12164
rect 7748 12112 7800 12164
rect 8208 12155 8260 12164
rect 8208 12121 8217 12155
rect 8217 12121 8251 12155
rect 8251 12121 8260 12155
rect 8208 12112 8260 12121
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 2320 12044 2372 12096
rect 2780 12044 2832 12096
rect 3056 12044 3108 12096
rect 4068 12087 4120 12096
rect 4068 12053 4077 12087
rect 4077 12053 4111 12087
rect 4111 12053 4120 12087
rect 4068 12044 4120 12053
rect 4896 12044 4948 12096
rect 9312 12112 9364 12164
rect 16488 12325 16497 12359
rect 16497 12325 16531 12359
rect 16531 12325 16540 12359
rect 16488 12316 16540 12325
rect 12716 12291 12768 12300
rect 12716 12257 12725 12291
rect 12725 12257 12759 12291
rect 12759 12257 12768 12291
rect 12716 12248 12768 12257
rect 15108 12248 15160 12300
rect 17316 12359 17368 12368
rect 17316 12325 17325 12359
rect 17325 12325 17359 12359
rect 17359 12325 17368 12359
rect 17316 12316 17368 12325
rect 16672 12248 16724 12300
rect 18696 12384 18748 12436
rect 19064 12384 19116 12436
rect 19432 12384 19484 12436
rect 19524 12384 19576 12436
rect 18052 12316 18104 12368
rect 19340 12248 19392 12300
rect 19708 12248 19760 12300
rect 14832 12180 14884 12232
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 16304 12223 16356 12232
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 17316 12180 17368 12232
rect 17500 12180 17552 12232
rect 17592 12180 17644 12232
rect 18328 12223 18380 12232
rect 18328 12189 18337 12223
rect 18337 12189 18371 12223
rect 18371 12189 18380 12223
rect 18328 12180 18380 12189
rect 19156 12180 19208 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 20352 12316 20404 12368
rect 20904 12316 20956 12368
rect 24124 12384 24176 12436
rect 25688 12384 25740 12436
rect 26148 12427 26200 12436
rect 26148 12393 26157 12427
rect 26157 12393 26191 12427
rect 26191 12393 26200 12427
rect 26148 12384 26200 12393
rect 26976 12384 27028 12436
rect 21732 12316 21784 12368
rect 20444 12180 20496 12232
rect 11152 12112 11204 12164
rect 16672 12112 16724 12164
rect 16948 12155 17000 12164
rect 16948 12121 16957 12155
rect 16957 12121 16991 12155
rect 16991 12121 17000 12155
rect 16948 12112 17000 12121
rect 19248 12155 19300 12164
rect 9036 12044 9088 12096
rect 15108 12044 15160 12096
rect 15292 12044 15344 12096
rect 15660 12044 15712 12096
rect 16120 12044 16172 12096
rect 16396 12044 16448 12096
rect 16488 12044 16540 12096
rect 17316 12044 17368 12096
rect 17592 12044 17644 12096
rect 19248 12121 19257 12155
rect 19257 12121 19291 12155
rect 19291 12121 19300 12155
rect 19248 12112 19300 12121
rect 19340 12112 19392 12164
rect 21732 12223 21784 12232
rect 21732 12189 21741 12223
rect 21741 12189 21775 12223
rect 21775 12189 21784 12223
rect 21732 12180 21784 12189
rect 22468 12180 22520 12232
rect 23204 12223 23256 12232
rect 23204 12189 23213 12223
rect 23213 12189 23247 12223
rect 23247 12189 23256 12223
rect 23204 12180 23256 12189
rect 20444 12044 20496 12096
rect 21180 12112 21232 12164
rect 28540 12316 28592 12368
rect 25228 12248 25280 12300
rect 27988 12248 28040 12300
rect 29552 12291 29604 12300
rect 29552 12257 29561 12291
rect 29561 12257 29595 12291
rect 29595 12257 29604 12291
rect 29552 12248 29604 12257
rect 27804 12180 27856 12232
rect 24400 12155 24452 12164
rect 24400 12121 24409 12155
rect 24409 12121 24443 12155
rect 24443 12121 24452 12155
rect 24400 12112 24452 12121
rect 24492 12112 24544 12164
rect 23296 12087 23348 12096
rect 23296 12053 23305 12087
rect 23305 12053 23339 12087
rect 23339 12053 23348 12087
rect 23296 12044 23348 12053
rect 23388 12044 23440 12096
rect 26700 12044 26752 12096
rect 27436 12044 27488 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 1860 11840 1912 11892
rect 3608 11840 3660 11892
rect 3976 11840 4028 11892
rect 1308 11772 1360 11824
rect 2964 11704 3016 11756
rect 3424 11747 3476 11756
rect 3424 11713 3433 11747
rect 3433 11713 3467 11747
rect 3467 11713 3476 11747
rect 3424 11704 3476 11713
rect 3516 11747 3568 11756
rect 3516 11713 3525 11747
rect 3525 11713 3559 11747
rect 3559 11713 3568 11747
rect 3516 11704 3568 11713
rect 3884 11704 3936 11756
rect 3976 11704 4028 11756
rect 4160 11840 4212 11892
rect 5724 11840 5776 11892
rect 8116 11840 8168 11892
rect 8392 11840 8444 11892
rect 12900 11840 12952 11892
rect 13360 11883 13412 11892
rect 13360 11849 13369 11883
rect 13369 11849 13403 11883
rect 13403 11849 13412 11883
rect 13360 11840 13412 11849
rect 4252 11704 4304 11756
rect 4712 11704 4764 11756
rect 6184 11772 6236 11824
rect 2504 11636 2556 11688
rect 2872 11636 2924 11688
rect 2228 11568 2280 11620
rect 4068 11568 4120 11620
rect 1584 11500 1636 11552
rect 3056 11500 3108 11552
rect 3976 11500 4028 11552
rect 6368 11704 6420 11756
rect 5264 11679 5316 11688
rect 5264 11645 5273 11679
rect 5273 11645 5307 11679
rect 5307 11645 5316 11679
rect 7748 11772 7800 11824
rect 10324 11815 10376 11824
rect 6828 11679 6880 11688
rect 5264 11636 5316 11645
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 8852 11636 8904 11688
rect 9036 11679 9088 11688
rect 9036 11645 9045 11679
rect 9045 11645 9079 11679
rect 9079 11645 9088 11679
rect 9036 11636 9088 11645
rect 10324 11781 10333 11815
rect 10333 11781 10367 11815
rect 10367 11781 10376 11815
rect 10324 11772 10376 11781
rect 11796 11815 11848 11824
rect 11796 11781 11830 11815
rect 11830 11781 11848 11815
rect 11796 11772 11848 11781
rect 15292 11840 15344 11892
rect 15752 11883 15804 11892
rect 15752 11849 15761 11883
rect 15761 11849 15795 11883
rect 15795 11849 15804 11883
rect 15752 11840 15804 11849
rect 16304 11840 16356 11892
rect 17500 11840 17552 11892
rect 18604 11840 18656 11892
rect 20260 11883 20312 11892
rect 20260 11849 20269 11883
rect 20269 11849 20303 11883
rect 20303 11849 20312 11883
rect 20260 11840 20312 11849
rect 20720 11840 20772 11892
rect 21824 11883 21876 11892
rect 21824 11849 21833 11883
rect 21833 11849 21867 11883
rect 21867 11849 21876 11883
rect 21824 11840 21876 11849
rect 22652 11883 22704 11892
rect 22652 11849 22661 11883
rect 22661 11849 22695 11883
rect 22695 11849 22704 11883
rect 22652 11840 22704 11849
rect 23480 11840 23532 11892
rect 24124 11840 24176 11892
rect 25320 11840 25372 11892
rect 27528 11883 27580 11892
rect 27528 11849 27537 11883
rect 27537 11849 27571 11883
rect 27571 11849 27580 11883
rect 27528 11840 27580 11849
rect 27804 11840 27856 11892
rect 28632 11883 28684 11892
rect 28632 11849 28641 11883
rect 28641 11849 28675 11883
rect 28675 11849 28684 11883
rect 28632 11840 28684 11849
rect 15016 11772 15068 11824
rect 15476 11815 15528 11824
rect 15476 11781 15485 11815
rect 15485 11781 15519 11815
rect 15519 11781 15528 11815
rect 15476 11772 15528 11781
rect 15936 11772 15988 11824
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 4988 11568 5040 11620
rect 6460 11568 6512 11620
rect 8392 11568 8444 11620
rect 12164 11704 12216 11756
rect 15568 11747 15620 11756
rect 11244 11636 11296 11688
rect 13268 11636 13320 11688
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 15292 11636 15344 11688
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 15752 11704 15804 11756
rect 16028 11636 16080 11688
rect 5632 11500 5684 11552
rect 7104 11500 7156 11552
rect 7564 11500 7616 11552
rect 9772 11500 9824 11552
rect 13452 11568 13504 11620
rect 10508 11500 10560 11552
rect 11520 11500 11572 11552
rect 14004 11500 14056 11552
rect 17040 11704 17092 11756
rect 19340 11772 19392 11824
rect 19708 11815 19760 11824
rect 19708 11781 19717 11815
rect 19717 11781 19751 11815
rect 19751 11781 19760 11815
rect 19708 11772 19760 11781
rect 18972 11704 19024 11756
rect 21548 11772 21600 11824
rect 22008 11815 22060 11824
rect 22008 11781 22017 11815
rect 22017 11781 22051 11815
rect 22051 11781 22060 11815
rect 22008 11772 22060 11781
rect 22100 11772 22152 11824
rect 27620 11772 27672 11824
rect 17500 11636 17552 11688
rect 19892 11704 19944 11756
rect 20168 11747 20220 11756
rect 20168 11713 20177 11747
rect 20177 11713 20211 11747
rect 20211 11713 20220 11747
rect 20168 11704 20220 11713
rect 20720 11704 20772 11756
rect 20996 11747 21048 11756
rect 20996 11713 21005 11747
rect 21005 11713 21039 11747
rect 21039 11713 21048 11747
rect 20996 11704 21048 11713
rect 21824 11704 21876 11756
rect 19156 11636 19208 11688
rect 19708 11636 19760 11688
rect 17776 11568 17828 11620
rect 20536 11636 20588 11688
rect 21916 11636 21968 11688
rect 24492 11704 24544 11756
rect 27988 11704 28040 11756
rect 20812 11611 20864 11620
rect 20812 11577 20821 11611
rect 20821 11577 20855 11611
rect 20855 11577 20864 11611
rect 20812 11568 20864 11577
rect 20996 11568 21048 11620
rect 21732 11568 21784 11620
rect 22836 11568 22888 11620
rect 28632 11636 28684 11688
rect 23664 11568 23716 11620
rect 31300 11568 31352 11620
rect 17500 11500 17552 11552
rect 18788 11500 18840 11552
rect 19616 11500 19668 11552
rect 19708 11500 19760 11552
rect 20076 11500 20128 11552
rect 23572 11543 23624 11552
rect 23572 11509 23581 11543
rect 23581 11509 23615 11543
rect 23615 11509 23624 11543
rect 23572 11500 23624 11509
rect 24492 11500 24544 11552
rect 25228 11543 25280 11552
rect 25228 11509 25237 11543
rect 25237 11509 25271 11543
rect 25271 11509 25280 11543
rect 25228 11500 25280 11509
rect 26976 11543 27028 11552
rect 26976 11509 26985 11543
rect 26985 11509 27019 11543
rect 27019 11509 27028 11543
rect 26976 11500 27028 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1492 11296 1544 11348
rect 2964 11296 3016 11348
rect 2872 11228 2924 11280
rect 3424 11296 3476 11348
rect 5172 11296 5224 11348
rect 6644 11296 6696 11348
rect 12624 11339 12676 11348
rect 5816 11228 5868 11280
rect 4252 11160 4304 11212
rect 5540 11203 5592 11212
rect 2320 11092 2372 11144
rect 3148 11092 3200 11144
rect 3424 11092 3476 11144
rect 3884 11024 3936 11076
rect 4528 11024 4580 11076
rect 5540 11169 5549 11203
rect 5549 11169 5583 11203
rect 5583 11169 5592 11203
rect 5540 11160 5592 11169
rect 6552 11203 6604 11212
rect 5448 11135 5500 11144
rect 5448 11101 5457 11135
rect 5457 11101 5491 11135
rect 5491 11101 5500 11135
rect 5448 11092 5500 11101
rect 4160 10999 4212 11008
rect 4160 10965 4169 10999
rect 4169 10965 4203 10999
rect 4203 10965 4212 10999
rect 4160 10956 4212 10965
rect 5540 11024 5592 11076
rect 5356 10956 5408 11008
rect 5724 10956 5776 11008
rect 6552 11169 6561 11203
rect 6561 11169 6595 11203
rect 6595 11169 6604 11203
rect 6552 11160 6604 11169
rect 8024 11160 8076 11212
rect 9312 11160 9364 11212
rect 9680 11160 9732 11212
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 7564 11135 7616 11144
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 11244 11135 11296 11144
rect 6000 11024 6052 11076
rect 6368 11024 6420 11076
rect 6644 11024 6696 11076
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 12624 11305 12633 11339
rect 12633 11305 12667 11339
rect 12667 11305 12676 11339
rect 12624 11296 12676 11305
rect 12992 11296 13044 11348
rect 14648 11296 14700 11348
rect 15292 11296 15344 11348
rect 15568 11296 15620 11348
rect 16120 11296 16172 11348
rect 16488 11296 16540 11348
rect 17868 11296 17920 11348
rect 19340 11296 19392 11348
rect 19708 11296 19760 11348
rect 20076 11339 20128 11348
rect 20076 11305 20085 11339
rect 20085 11305 20119 11339
rect 20119 11305 20128 11339
rect 20076 11296 20128 11305
rect 21088 11296 21140 11348
rect 22560 11339 22612 11348
rect 22560 11305 22569 11339
rect 22569 11305 22603 11339
rect 22603 11305 22612 11339
rect 22560 11296 22612 11305
rect 23204 11296 23256 11348
rect 12900 11160 12952 11212
rect 13636 11228 13688 11280
rect 13912 11228 13964 11280
rect 14740 11228 14792 11280
rect 15200 11160 15252 11212
rect 9128 11024 9180 11076
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 13544 11092 13596 11144
rect 14740 11092 14792 11144
rect 13176 11024 13228 11076
rect 14004 11024 14056 11076
rect 14648 11067 14700 11076
rect 14648 11033 14657 11067
rect 14657 11033 14691 11067
rect 14691 11033 14700 11067
rect 15844 11160 15896 11212
rect 16028 11203 16080 11212
rect 16028 11169 16037 11203
rect 16037 11169 16071 11203
rect 16071 11169 16080 11203
rect 16028 11160 16080 11169
rect 15660 11092 15712 11144
rect 16120 11135 16172 11144
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 17132 11160 17184 11212
rect 20720 11160 20772 11212
rect 23296 11228 23348 11280
rect 23664 11296 23716 11348
rect 24400 11339 24452 11348
rect 24400 11305 24409 11339
rect 24409 11305 24443 11339
rect 24443 11305 24452 11339
rect 24400 11296 24452 11305
rect 27252 11339 27304 11348
rect 27252 11305 27261 11339
rect 27261 11305 27295 11339
rect 27295 11305 27304 11339
rect 27252 11296 27304 11305
rect 32036 11228 32088 11280
rect 23756 11160 23808 11212
rect 24768 11160 24820 11212
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 18880 11092 18932 11144
rect 20628 11092 20680 11144
rect 14648 11024 14700 11033
rect 17040 11024 17092 11076
rect 8944 10956 8996 11008
rect 10784 10956 10836 11008
rect 12992 10956 13044 11008
rect 15016 10956 15068 11008
rect 15200 10956 15252 11008
rect 16672 10956 16724 11008
rect 18052 11024 18104 11076
rect 18696 11024 18748 11076
rect 19156 11024 19208 11076
rect 20168 11024 20220 11076
rect 20260 11067 20312 11076
rect 20260 11033 20269 11067
rect 20269 11033 20303 11067
rect 20303 11033 20312 11067
rect 20444 11067 20496 11076
rect 20260 11024 20312 11033
rect 20444 11033 20453 11067
rect 20453 11033 20487 11067
rect 20487 11033 20496 11067
rect 20444 11024 20496 11033
rect 21364 11092 21416 11144
rect 22836 11092 22888 11144
rect 23664 11135 23716 11144
rect 23664 11101 23673 11135
rect 23673 11101 23707 11135
rect 23707 11101 23716 11135
rect 23664 11092 23716 11101
rect 24216 11092 24268 11144
rect 21088 11067 21140 11076
rect 18328 10956 18380 11008
rect 18788 10956 18840 11008
rect 21088 11033 21097 11067
rect 21097 11033 21131 11067
rect 21131 11033 21140 11067
rect 21088 11024 21140 11033
rect 21548 11024 21600 11076
rect 20628 10956 20680 11008
rect 22468 10956 22520 11008
rect 22744 11067 22796 11076
rect 22744 11033 22753 11067
rect 22753 11033 22787 11067
rect 22787 11033 22796 11067
rect 22928 11067 22980 11076
rect 22744 11024 22796 11033
rect 22928 11033 22937 11067
rect 22937 11033 22971 11067
rect 22971 11033 22980 11067
rect 22928 11024 22980 11033
rect 24124 11024 24176 11076
rect 25688 11067 25740 11076
rect 25688 11033 25697 11067
rect 25697 11033 25731 11067
rect 25731 11033 25740 11067
rect 25688 11024 25740 11033
rect 26240 11067 26292 11076
rect 26240 11033 26249 11067
rect 26249 11033 26283 11067
rect 26283 11033 26292 11067
rect 26240 11024 26292 11033
rect 24308 10956 24360 11008
rect 24676 10956 24728 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 2136 10752 2188 10804
rect 2412 10752 2464 10804
rect 3332 10752 3384 10804
rect 5724 10752 5776 10804
rect 7564 10752 7616 10804
rect 7748 10752 7800 10804
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 2412 10616 2464 10668
rect 572 10548 624 10600
rect 1584 10523 1636 10532
rect 1584 10489 1593 10523
rect 1593 10489 1627 10523
rect 1627 10489 1636 10523
rect 1584 10480 1636 10489
rect 2504 10548 2556 10600
rect 5264 10684 5316 10736
rect 5540 10684 5592 10736
rect 6460 10727 6512 10736
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 3792 10616 3844 10668
rect 4252 10616 4304 10668
rect 4988 10616 5040 10668
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 6460 10693 6469 10727
rect 6469 10693 6503 10727
rect 6503 10693 6512 10727
rect 6460 10684 6512 10693
rect 6644 10684 6696 10736
rect 8300 10684 8352 10736
rect 8484 10752 8536 10804
rect 10508 10752 10560 10804
rect 10600 10752 10652 10804
rect 10876 10752 10928 10804
rect 11980 10752 12032 10804
rect 12256 10752 12308 10804
rect 12440 10752 12492 10804
rect 13452 10752 13504 10804
rect 14556 10795 14608 10804
rect 14556 10761 14565 10795
rect 14565 10761 14599 10795
rect 14599 10761 14608 10795
rect 14556 10752 14608 10761
rect 14924 10795 14976 10804
rect 14924 10761 14933 10795
rect 14933 10761 14967 10795
rect 14967 10761 14976 10795
rect 14924 10752 14976 10761
rect 15292 10752 15344 10804
rect 15660 10752 15712 10804
rect 9496 10684 9548 10736
rect 10140 10684 10192 10736
rect 5816 10616 5868 10668
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 4528 10548 4580 10600
rect 5448 10548 5500 10600
rect 6276 10548 6328 10600
rect 7288 10548 7340 10600
rect 7380 10548 7432 10600
rect 3792 10480 3844 10532
rect 2780 10412 2832 10464
rect 3976 10412 4028 10464
rect 4896 10455 4948 10464
rect 4896 10421 4905 10455
rect 4905 10421 4939 10455
rect 4939 10421 4948 10455
rect 4896 10412 4948 10421
rect 5172 10412 5224 10464
rect 5540 10412 5592 10464
rect 6276 10412 6328 10464
rect 7012 10412 7064 10464
rect 8300 10412 8352 10464
rect 10416 10616 10468 10668
rect 11612 10616 11664 10668
rect 13544 10727 13596 10736
rect 13544 10693 13553 10727
rect 13553 10693 13587 10727
rect 13587 10693 13596 10727
rect 13544 10684 13596 10693
rect 11244 10548 11296 10600
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 8668 10480 8720 10532
rect 9772 10480 9824 10532
rect 13268 10480 13320 10532
rect 12716 10412 12768 10464
rect 13452 10591 13504 10600
rect 13452 10557 13461 10591
rect 13461 10557 13495 10591
rect 13495 10557 13504 10591
rect 14280 10616 14332 10668
rect 14832 10616 14884 10668
rect 13452 10548 13504 10557
rect 15568 10548 15620 10600
rect 19432 10752 19484 10804
rect 19984 10752 20036 10804
rect 21640 10752 21692 10804
rect 22008 10752 22060 10804
rect 23664 10752 23716 10804
rect 24768 10752 24820 10804
rect 26700 10752 26752 10804
rect 28264 10752 28316 10804
rect 19248 10727 19300 10736
rect 19248 10693 19257 10727
rect 19257 10693 19291 10727
rect 19291 10693 19300 10727
rect 19248 10684 19300 10693
rect 22192 10684 22244 10736
rect 22744 10684 22796 10736
rect 23296 10684 23348 10736
rect 25504 10684 25556 10736
rect 32128 10684 32180 10736
rect 16580 10616 16632 10668
rect 18144 10616 18196 10668
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 17684 10591 17736 10600
rect 17684 10557 17693 10591
rect 17693 10557 17727 10591
rect 17727 10557 17736 10591
rect 17684 10548 17736 10557
rect 18696 10616 18748 10668
rect 20352 10616 20404 10668
rect 26976 10659 27028 10668
rect 18972 10548 19024 10600
rect 14004 10523 14056 10532
rect 14004 10489 14013 10523
rect 14013 10489 14047 10523
rect 14047 10489 14056 10523
rect 14004 10480 14056 10489
rect 14280 10480 14332 10532
rect 14832 10480 14884 10532
rect 16488 10480 16540 10532
rect 18512 10480 18564 10532
rect 18880 10523 18932 10532
rect 18880 10489 18889 10523
rect 18889 10489 18923 10523
rect 18923 10489 18932 10523
rect 19892 10523 19944 10532
rect 18880 10480 18932 10489
rect 19892 10489 19901 10523
rect 19901 10489 19935 10523
rect 19935 10489 19944 10523
rect 19892 10480 19944 10489
rect 20260 10548 20312 10600
rect 26976 10625 26985 10659
rect 26985 10625 27019 10659
rect 27019 10625 27028 10659
rect 26976 10616 27028 10625
rect 21364 10548 21416 10600
rect 22008 10548 22060 10600
rect 24676 10548 24728 10600
rect 25596 10548 25648 10600
rect 32220 10548 32272 10600
rect 20536 10480 20588 10532
rect 23204 10480 23256 10532
rect 30564 10480 30616 10532
rect 15200 10412 15252 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 15936 10455 15988 10464
rect 15936 10421 15945 10455
rect 15945 10421 15979 10455
rect 15979 10421 15988 10455
rect 15936 10412 15988 10421
rect 16672 10455 16724 10464
rect 16672 10421 16681 10455
rect 16681 10421 16715 10455
rect 16715 10421 16724 10455
rect 16672 10412 16724 10421
rect 18788 10455 18840 10464
rect 18788 10421 18797 10455
rect 18797 10421 18831 10455
rect 18831 10421 18840 10455
rect 18788 10412 18840 10421
rect 20996 10412 21048 10464
rect 21916 10455 21968 10464
rect 21916 10421 21925 10455
rect 21925 10421 21959 10455
rect 21959 10421 21968 10455
rect 21916 10412 21968 10421
rect 24124 10412 24176 10464
rect 26332 10412 26384 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 2688 10208 2740 10260
rect 5540 10251 5592 10260
rect 2596 10183 2648 10192
rect 2596 10149 2605 10183
rect 2605 10149 2639 10183
rect 2639 10149 2648 10183
rect 2596 10140 2648 10149
rect 2320 10072 2372 10124
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 4620 10140 4672 10192
rect 5080 10140 5132 10192
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 6092 10208 6144 10260
rect 6184 10208 6236 10260
rect 7472 10208 7524 10260
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 10600 10208 10652 10260
rect 11612 10208 11664 10260
rect 14556 10208 14608 10260
rect 15108 10208 15160 10260
rect 17592 10208 17644 10260
rect 17960 10208 18012 10260
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 18512 10208 18564 10260
rect 3608 10072 3660 10124
rect 3884 10072 3936 10124
rect 4528 10072 4580 10124
rect 5448 10072 5500 10124
rect 5724 10072 5776 10124
rect 6644 10072 6696 10124
rect 4068 10004 4120 10056
rect 4160 10004 4212 10056
rect 5816 10047 5868 10056
rect 2136 9936 2188 9988
rect 2228 9936 2280 9988
rect 3976 9979 4028 9988
rect 3976 9945 3985 9979
rect 3985 9945 4019 9979
rect 4019 9945 4028 9979
rect 3976 9936 4028 9945
rect 4528 9936 4580 9988
rect 3884 9868 3936 9920
rect 5080 9911 5132 9920
rect 5080 9877 5089 9911
rect 5089 9877 5123 9911
rect 5123 9877 5132 9911
rect 5080 9868 5132 9877
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 6460 10004 6512 10056
rect 9220 10140 9272 10192
rect 10140 10140 10192 10192
rect 12716 10140 12768 10192
rect 12992 10140 13044 10192
rect 15292 10183 15344 10192
rect 15292 10149 15301 10183
rect 15301 10149 15335 10183
rect 15335 10149 15344 10183
rect 15292 10140 15344 10149
rect 16764 10140 16816 10192
rect 7748 10115 7800 10124
rect 7748 10081 7757 10115
rect 7757 10081 7791 10115
rect 7791 10081 7800 10115
rect 7748 10072 7800 10081
rect 7932 10115 7984 10124
rect 7932 10081 7941 10115
rect 7941 10081 7975 10115
rect 7975 10081 7984 10115
rect 7932 10072 7984 10081
rect 8024 10072 8076 10124
rect 5356 9936 5408 9988
rect 6368 9936 6420 9988
rect 6644 9936 6696 9988
rect 7288 9936 7340 9988
rect 8944 10047 8996 10056
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 13544 10072 13596 10124
rect 15568 10072 15620 10124
rect 15660 10072 15712 10124
rect 17868 10140 17920 10192
rect 18972 10140 19024 10192
rect 19340 10140 19392 10192
rect 20536 10140 20588 10192
rect 21548 10208 21600 10260
rect 23296 10251 23348 10260
rect 23296 10217 23305 10251
rect 23305 10217 23339 10251
rect 23339 10217 23348 10251
rect 23296 10208 23348 10217
rect 24860 10208 24912 10260
rect 30656 10208 30708 10260
rect 43352 10251 43404 10260
rect 43352 10217 43361 10251
rect 43361 10217 43395 10251
rect 43395 10217 43404 10251
rect 43352 10208 43404 10217
rect 25504 10140 25556 10192
rect 25780 10140 25832 10192
rect 22652 10072 22704 10124
rect 7656 9868 7708 9920
rect 7748 9868 7800 9920
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 9036 9936 9088 9988
rect 10416 10004 10468 10056
rect 11520 10004 11572 10056
rect 12348 10004 12400 10056
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 14556 10047 14608 10056
rect 14556 10013 14565 10047
rect 14565 10013 14599 10047
rect 14599 10013 14608 10047
rect 15016 10047 15068 10056
rect 14556 10004 14608 10013
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17727 10047
rect 17727 10013 17736 10047
rect 17684 10004 17736 10013
rect 17868 10004 17920 10056
rect 18696 10004 18748 10056
rect 19248 10047 19300 10056
rect 19248 10013 19257 10047
rect 19257 10013 19291 10047
rect 19291 10013 19300 10047
rect 19248 10004 19300 10013
rect 20352 10004 20404 10056
rect 10600 9936 10652 9988
rect 11796 9936 11848 9988
rect 16672 9936 16724 9988
rect 16764 9979 16816 9988
rect 16764 9945 16773 9979
rect 16773 9945 16807 9979
rect 16807 9945 16816 9979
rect 16764 9936 16816 9945
rect 17224 9936 17276 9988
rect 18512 9979 18564 9988
rect 18512 9945 18521 9979
rect 18521 9945 18555 9979
rect 18555 9945 18564 9979
rect 18512 9936 18564 9945
rect 12992 9868 13044 9920
rect 14280 9868 14332 9920
rect 14924 9868 14976 9920
rect 15200 9868 15252 9920
rect 19432 9868 19484 9920
rect 20628 9936 20680 9988
rect 22468 10004 22520 10056
rect 25596 10004 25648 10056
rect 27252 10072 27304 10124
rect 28356 10072 28408 10124
rect 27896 10004 27948 10056
rect 29000 10047 29052 10056
rect 29000 10013 29009 10047
rect 29009 10013 29043 10047
rect 29043 10013 29052 10047
rect 29000 10004 29052 10013
rect 43352 10004 43404 10056
rect 21180 9936 21232 9988
rect 24860 9936 24912 9988
rect 25504 9936 25556 9988
rect 26792 9936 26844 9988
rect 21732 9868 21784 9920
rect 22008 9868 22060 9920
rect 22192 9868 22244 9920
rect 24032 9868 24084 9920
rect 24308 9868 24360 9920
rect 27620 9868 27672 9920
rect 27988 9868 28040 9920
rect 44088 9911 44140 9920
rect 44088 9877 44097 9911
rect 44097 9877 44131 9911
rect 44131 9877 44140 9911
rect 44088 9868 44140 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2228 9664 2280 9716
rect 2412 9664 2464 9716
rect 3608 9664 3660 9716
rect 4344 9664 4396 9716
rect 6552 9664 6604 9716
rect 1952 9596 2004 9648
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 2412 9571 2464 9580
rect 2412 9537 2421 9571
rect 2421 9537 2455 9571
rect 2455 9537 2464 9571
rect 2412 9528 2464 9537
rect 3792 9596 3844 9648
rect 4344 9528 4396 9580
rect 4620 9528 4672 9580
rect 3424 9460 3476 9512
rect 5172 9528 5224 9580
rect 5816 9596 5868 9648
rect 7380 9664 7432 9716
rect 9128 9664 9180 9716
rect 9312 9664 9364 9716
rect 9772 9664 9824 9716
rect 9956 9664 10008 9716
rect 10508 9664 10560 9716
rect 10692 9664 10744 9716
rect 14556 9664 14608 9716
rect 6000 9528 6052 9580
rect 6368 9528 6420 9580
rect 7288 9596 7340 9648
rect 7380 9528 7432 9580
rect 5448 9460 5500 9512
rect 7932 9528 7984 9580
rect 8208 9528 8260 9580
rect 9312 9528 9364 9580
rect 7656 9503 7708 9512
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 8484 9460 8536 9512
rect 9496 9460 9548 9512
rect 9772 9528 9824 9580
rect 10232 9460 10284 9512
rect 11612 9460 11664 9512
rect 16948 9664 17000 9716
rect 17776 9664 17828 9716
rect 15844 9596 15896 9648
rect 17684 9596 17736 9648
rect 13912 9528 13964 9580
rect 12992 9460 13044 9512
rect 15016 9528 15068 9580
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 16396 9528 16448 9580
rect 1032 9392 1084 9444
rect 3516 9435 3568 9444
rect 3516 9401 3525 9435
rect 3525 9401 3559 9435
rect 3559 9401 3568 9435
rect 3516 9392 3568 9401
rect 3608 9392 3660 9444
rect 1952 9367 2004 9376
rect 1952 9333 1961 9367
rect 1961 9333 1995 9367
rect 1995 9333 2004 9367
rect 1952 9324 2004 9333
rect 5356 9324 5408 9376
rect 7840 9392 7892 9444
rect 13360 9392 13412 9444
rect 14464 9392 14516 9444
rect 14648 9392 14700 9444
rect 6184 9324 6236 9376
rect 6276 9324 6328 9376
rect 7472 9367 7524 9376
rect 7472 9333 7481 9367
rect 7481 9333 7515 9367
rect 7515 9333 7524 9367
rect 7472 9324 7524 9333
rect 7656 9324 7708 9376
rect 8024 9324 8076 9376
rect 8300 9324 8352 9376
rect 10876 9367 10928 9376
rect 10876 9333 10885 9367
rect 10885 9333 10919 9367
rect 10919 9333 10928 9367
rect 10876 9324 10928 9333
rect 11888 9324 11940 9376
rect 15200 9460 15252 9512
rect 17868 9528 17920 9580
rect 18328 9596 18380 9648
rect 18512 9596 18564 9648
rect 19064 9664 19116 9716
rect 21916 9664 21968 9716
rect 16580 9460 16632 9512
rect 16672 9460 16724 9512
rect 17224 9460 17276 9512
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 18328 9460 18380 9512
rect 14924 9435 14976 9444
rect 14924 9401 14933 9435
rect 14933 9401 14967 9435
rect 14967 9401 14976 9435
rect 14924 9392 14976 9401
rect 15752 9392 15804 9444
rect 16488 9392 16540 9444
rect 17040 9435 17092 9444
rect 17040 9401 17049 9435
rect 17049 9401 17083 9435
rect 17083 9401 17092 9435
rect 17592 9435 17644 9444
rect 17040 9392 17092 9401
rect 17592 9401 17601 9435
rect 17601 9401 17635 9435
rect 17635 9401 17644 9435
rect 17592 9392 17644 9401
rect 20352 9596 20404 9648
rect 20720 9596 20772 9648
rect 22100 9664 22152 9716
rect 25228 9664 25280 9716
rect 27252 9707 27304 9716
rect 27252 9673 27261 9707
rect 27261 9673 27295 9707
rect 27295 9673 27304 9707
rect 27252 9664 27304 9673
rect 27896 9664 27948 9716
rect 24216 9639 24268 9648
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 18788 9460 18840 9512
rect 19064 9503 19116 9512
rect 19064 9469 19073 9503
rect 19073 9469 19107 9503
rect 19107 9469 19116 9503
rect 19064 9460 19116 9469
rect 19248 9460 19300 9512
rect 21732 9528 21784 9580
rect 24216 9605 24225 9639
rect 24225 9605 24259 9639
rect 24259 9605 24268 9639
rect 24216 9596 24268 9605
rect 25964 9639 26016 9648
rect 25964 9605 25973 9639
rect 25973 9605 26007 9639
rect 26007 9605 26016 9639
rect 25964 9596 26016 9605
rect 19892 9392 19944 9444
rect 22744 9528 22796 9580
rect 26700 9528 26752 9580
rect 23388 9460 23440 9512
rect 15108 9324 15160 9376
rect 16672 9324 16724 9376
rect 16948 9324 17000 9376
rect 17960 9324 18012 9376
rect 22100 9392 22152 9444
rect 22376 9392 22428 9444
rect 22468 9392 22520 9444
rect 27344 9460 27396 9512
rect 20628 9324 20680 9376
rect 21456 9324 21508 9376
rect 22560 9324 22612 9376
rect 22652 9367 22704 9376
rect 22652 9333 22661 9367
rect 22661 9333 22695 9367
rect 22695 9333 22704 9367
rect 22652 9324 22704 9333
rect 27068 9324 27120 9376
rect 42156 9324 42208 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1400 9163 1452 9172
rect 1400 9129 1409 9163
rect 1409 9129 1443 9163
rect 1443 9129 1452 9163
rect 1400 9120 1452 9129
rect 1676 9120 1728 9172
rect 2136 9120 2188 9172
rect 5448 9120 5500 9172
rect 6736 9120 6788 9172
rect 5724 9052 5776 9104
rect 6184 9052 6236 9104
rect 7104 9095 7156 9104
rect 7104 9061 7113 9095
rect 7113 9061 7147 9095
rect 7147 9061 7156 9095
rect 7104 9052 7156 9061
rect 7472 9120 7524 9172
rect 9036 9120 9088 9172
rect 7656 9052 7708 9104
rect 7840 9052 7892 9104
rect 1768 8984 1820 9036
rect 1492 8916 1544 8968
rect 1768 8848 1820 8900
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3240 8916 3292 8968
rect 3792 8916 3844 8968
rect 4620 8916 4672 8968
rect 5448 8916 5500 8968
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 6092 8916 6144 8968
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 3332 8848 3384 8900
rect 6184 8848 6236 8900
rect 6736 8916 6788 8968
rect 7288 8916 7340 8968
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 8668 9052 8720 9104
rect 8576 8984 8628 9036
rect 11060 9120 11112 9172
rect 11980 9163 12032 9172
rect 11980 9129 11989 9163
rect 11989 9129 12023 9163
rect 12023 9129 12032 9163
rect 11980 9120 12032 9129
rect 13084 9120 13136 9172
rect 14188 9120 14240 9172
rect 14372 9120 14424 9172
rect 16488 9163 16540 9172
rect 16488 9129 16497 9163
rect 16497 9129 16531 9163
rect 16531 9129 16540 9163
rect 16488 9120 16540 9129
rect 16580 9120 16632 9172
rect 16856 9120 16908 9172
rect 17224 9120 17276 9172
rect 17592 9120 17644 9172
rect 18512 9120 18564 9172
rect 20076 9120 20128 9172
rect 9956 9052 10008 9104
rect 10232 9052 10284 9104
rect 10784 9052 10836 9104
rect 13544 9052 13596 9104
rect 14004 9052 14056 9104
rect 14924 9052 14976 9104
rect 15936 9095 15988 9104
rect 15936 9061 15945 9095
rect 15945 9061 15979 9095
rect 15979 9061 15988 9095
rect 15936 9052 15988 9061
rect 16764 9052 16816 9104
rect 9312 8984 9364 9036
rect 10968 8984 11020 9036
rect 11612 8984 11664 9036
rect 11980 8984 12032 9036
rect 12624 9027 12676 9036
rect 12624 8993 12633 9027
rect 12633 8993 12667 9027
rect 12667 8993 12676 9027
rect 12624 8984 12676 8993
rect 13452 8984 13504 9036
rect 18696 9052 18748 9104
rect 19984 9095 20036 9104
rect 19984 9061 19993 9095
rect 19993 9061 20027 9095
rect 20027 9061 20036 9095
rect 19984 9052 20036 9061
rect 7288 8780 7340 8832
rect 7472 8891 7524 8900
rect 7472 8857 7481 8891
rect 7481 8857 7515 8891
rect 7515 8857 7524 8891
rect 7472 8848 7524 8857
rect 8300 8916 8352 8968
rect 8484 8916 8536 8968
rect 9036 8848 9088 8900
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 10140 8916 10192 8968
rect 10508 8916 10560 8968
rect 8116 8780 8168 8832
rect 9680 8848 9732 8900
rect 11244 8848 11296 8900
rect 11612 8848 11664 8900
rect 11796 8848 11848 8900
rect 13360 8916 13412 8968
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 14924 8916 14976 8925
rect 16764 8916 16816 8968
rect 17224 8916 17276 8968
rect 17500 8916 17552 8968
rect 20536 9120 20588 9172
rect 22100 9120 22152 9172
rect 24492 9120 24544 9172
rect 25964 9120 26016 9172
rect 26424 9120 26476 9172
rect 26976 9163 27028 9172
rect 26976 9129 26985 9163
rect 26985 9129 27019 9163
rect 27019 9129 27028 9163
rect 26976 9120 27028 9129
rect 27068 9120 27120 9172
rect 41420 9120 41472 9172
rect 20812 9052 20864 9104
rect 22468 9052 22520 9104
rect 23664 9052 23716 9104
rect 31208 9052 31260 9104
rect 20996 8984 21048 9036
rect 22560 9027 22612 9036
rect 22560 8993 22569 9027
rect 22569 8993 22603 9027
rect 22603 8993 22612 9027
rect 22560 8984 22612 8993
rect 24124 8984 24176 9036
rect 27436 8984 27488 9036
rect 21640 8959 21692 8968
rect 21640 8925 21649 8959
rect 21649 8925 21683 8959
rect 21683 8925 21692 8959
rect 21640 8916 21692 8925
rect 33324 9052 33376 9104
rect 15200 8848 15252 8900
rect 15752 8848 15804 8900
rect 17040 8848 17092 8900
rect 18052 8891 18104 8900
rect 18052 8857 18061 8891
rect 18061 8857 18095 8891
rect 18095 8857 18104 8891
rect 18052 8848 18104 8857
rect 18512 8848 18564 8900
rect 11336 8780 11388 8832
rect 12992 8780 13044 8832
rect 13360 8780 13412 8832
rect 14556 8780 14608 8832
rect 14924 8780 14976 8832
rect 16212 8780 16264 8832
rect 17500 8780 17552 8832
rect 20076 8848 20128 8900
rect 20260 8891 20312 8900
rect 20260 8857 20269 8891
rect 20269 8857 20303 8891
rect 20303 8857 20312 8891
rect 20260 8848 20312 8857
rect 20352 8848 20404 8900
rect 23664 8891 23716 8900
rect 23664 8857 23673 8891
rect 23673 8857 23707 8891
rect 23707 8857 23716 8891
rect 23664 8848 23716 8857
rect 26976 8848 27028 8900
rect 23756 8823 23808 8832
rect 23756 8789 23765 8823
rect 23765 8789 23799 8823
rect 23799 8789 23808 8823
rect 23756 8780 23808 8789
rect 23848 8780 23900 8832
rect 24216 8780 24268 8832
rect 25044 8823 25096 8832
rect 25044 8789 25053 8823
rect 25053 8789 25087 8823
rect 25087 8789 25096 8823
rect 25044 8780 25096 8789
rect 27712 8823 27764 8832
rect 27712 8789 27721 8823
rect 27721 8789 27755 8823
rect 27755 8789 27764 8823
rect 27712 8780 27764 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1860 8576 1912 8628
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 2320 8576 2372 8628
rect 3424 8619 3476 8628
rect 3424 8585 3433 8619
rect 3433 8585 3467 8619
rect 3467 8585 3476 8619
rect 3424 8576 3476 8585
rect 4804 8576 4856 8628
rect 7196 8576 7248 8628
rect 3976 8508 4028 8560
rect 6828 8551 6880 8560
rect 6828 8517 6837 8551
rect 6837 8517 6871 8551
rect 6871 8517 6880 8551
rect 6828 8508 6880 8517
rect 6920 8508 6972 8560
rect 7840 8508 7892 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 2228 8483 2280 8492
rect 2228 8449 2237 8483
rect 2237 8449 2271 8483
rect 2271 8449 2280 8483
rect 2228 8440 2280 8449
rect 3148 8440 3200 8492
rect 4712 8440 4764 8492
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 5632 8440 5684 8492
rect 7012 8440 7064 8492
rect 7196 8440 7248 8492
rect 8208 8508 8260 8560
rect 8760 8576 8812 8628
rect 9956 8576 10008 8628
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 11428 8576 11480 8628
rect 12164 8576 12216 8628
rect 5264 8372 5316 8424
rect 9312 8440 9364 8492
rect 9496 8440 9548 8492
rect 10140 8483 10192 8492
rect 3240 8304 3292 8356
rect 5908 8304 5960 8356
rect 7380 8372 7432 8424
rect 3884 8236 3936 8288
rect 4068 8236 4120 8288
rect 5264 8236 5316 8288
rect 5448 8236 5500 8288
rect 6920 8304 6972 8356
rect 7748 8304 7800 8356
rect 8300 8372 8352 8424
rect 9128 8372 9180 8424
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 10784 8508 10836 8560
rect 8116 8304 8168 8356
rect 8392 8347 8444 8356
rect 8392 8313 8401 8347
rect 8401 8313 8435 8347
rect 8435 8313 8444 8347
rect 8392 8304 8444 8313
rect 8668 8304 8720 8356
rect 9956 8372 10008 8424
rect 12164 8440 12216 8492
rect 12716 8576 12768 8628
rect 12808 8551 12860 8560
rect 12808 8517 12817 8551
rect 12817 8517 12851 8551
rect 12851 8517 12860 8551
rect 12808 8508 12860 8517
rect 13452 8508 13504 8560
rect 14096 8508 14148 8560
rect 17868 8576 17920 8628
rect 19156 8576 19208 8628
rect 20168 8576 20220 8628
rect 21640 8576 21692 8628
rect 21732 8576 21784 8628
rect 22744 8576 22796 8628
rect 25504 8619 25556 8628
rect 25504 8585 25513 8619
rect 25513 8585 25547 8619
rect 25547 8585 25556 8619
rect 25504 8576 25556 8585
rect 27712 8576 27764 8628
rect 42984 8576 43036 8628
rect 14924 8508 14976 8560
rect 16212 8508 16264 8560
rect 19248 8508 19300 8560
rect 20076 8508 20128 8560
rect 22560 8551 22612 8560
rect 22560 8517 22569 8551
rect 22569 8517 22603 8551
rect 22603 8517 22612 8551
rect 22560 8508 22612 8517
rect 23756 8508 23808 8560
rect 40776 8508 40828 8560
rect 11060 8372 11112 8424
rect 12348 8372 12400 8424
rect 12716 8304 12768 8356
rect 15108 8372 15160 8424
rect 15568 8440 15620 8492
rect 15752 8440 15804 8492
rect 17776 8440 17828 8492
rect 18512 8483 18564 8492
rect 18512 8449 18521 8483
rect 18521 8449 18555 8483
rect 18555 8449 18564 8483
rect 18512 8440 18564 8449
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 15384 8347 15436 8356
rect 15384 8313 15393 8347
rect 15393 8313 15427 8347
rect 15427 8313 15436 8347
rect 15384 8304 15436 8313
rect 8024 8236 8076 8288
rect 8208 8236 8260 8288
rect 9128 8236 9180 8288
rect 12992 8279 13044 8288
rect 12992 8245 13001 8279
rect 13001 8245 13035 8279
rect 13035 8245 13044 8279
rect 12992 8236 13044 8245
rect 13544 8236 13596 8288
rect 15568 8236 15620 8288
rect 16028 8415 16080 8424
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 16028 8372 16080 8381
rect 16580 8372 16632 8424
rect 21272 8440 21324 8492
rect 22376 8440 22428 8492
rect 26332 8440 26384 8492
rect 20260 8415 20312 8424
rect 20260 8381 20269 8415
rect 20269 8381 20303 8415
rect 20303 8381 20312 8415
rect 20260 8372 20312 8381
rect 25964 8415 26016 8424
rect 16948 8347 17000 8356
rect 16948 8313 16957 8347
rect 16957 8313 16991 8347
rect 16991 8313 17000 8347
rect 16948 8304 17000 8313
rect 17592 8304 17644 8356
rect 19524 8347 19576 8356
rect 16672 8236 16724 8288
rect 16856 8236 16908 8288
rect 17960 8236 18012 8288
rect 18604 8236 18656 8288
rect 19524 8313 19533 8347
rect 19533 8313 19567 8347
rect 19567 8313 19576 8347
rect 19524 8304 19576 8313
rect 19892 8304 19944 8356
rect 20352 8304 20404 8356
rect 20536 8347 20588 8356
rect 20536 8313 20545 8347
rect 20545 8313 20579 8347
rect 20579 8313 20588 8347
rect 20536 8304 20588 8313
rect 20812 8304 20864 8356
rect 20996 8304 21048 8356
rect 21272 8347 21324 8356
rect 21272 8313 21281 8347
rect 21281 8313 21315 8347
rect 21315 8313 21324 8347
rect 21272 8304 21324 8313
rect 22744 8347 22796 8356
rect 21916 8279 21968 8288
rect 21916 8245 21925 8279
rect 21925 8245 21959 8279
rect 21959 8245 21968 8279
rect 21916 8236 21968 8245
rect 22744 8313 22753 8347
rect 22753 8313 22787 8347
rect 22787 8313 22796 8347
rect 22744 8304 22796 8313
rect 23480 8304 23532 8356
rect 23848 8347 23900 8356
rect 23848 8313 23857 8347
rect 23857 8313 23891 8347
rect 23891 8313 23900 8347
rect 23848 8304 23900 8313
rect 25964 8381 25973 8415
rect 25973 8381 26007 8415
rect 26007 8381 26016 8415
rect 25964 8372 26016 8381
rect 26884 8304 26936 8356
rect 23388 8236 23440 8288
rect 28632 8236 28684 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2044 8075 2096 8084
rect 2044 8041 2053 8075
rect 2053 8041 2087 8075
rect 2087 8041 2096 8075
rect 2044 8032 2096 8041
rect 2596 8075 2648 8084
rect 2596 8041 2605 8075
rect 2605 8041 2639 8075
rect 2639 8041 2648 8075
rect 2596 8032 2648 8041
rect 3240 8075 3292 8084
rect 3240 8041 3249 8075
rect 3249 8041 3283 8075
rect 3283 8041 3292 8075
rect 3240 8032 3292 8041
rect 3792 8075 3844 8084
rect 3792 8041 3801 8075
rect 3801 8041 3835 8075
rect 3835 8041 3844 8075
rect 3792 8032 3844 8041
rect 6184 8075 6236 8084
rect 6184 8041 6193 8075
rect 6193 8041 6227 8075
rect 6227 8041 6236 8075
rect 6184 8032 6236 8041
rect 6736 8032 6788 8084
rect 6920 8032 6972 8084
rect 7472 8032 7524 8084
rect 7564 8032 7616 8084
rect 9956 8032 10008 8084
rect 12072 8032 12124 8084
rect 12992 8032 13044 8084
rect 1216 7964 1268 8016
rect 8300 7964 8352 8016
rect 9404 7964 9456 8016
rect 13268 7964 13320 8016
rect 15384 7964 15436 8016
rect 15752 7964 15804 8016
rect 17408 8032 17460 8084
rect 18604 8075 18656 8084
rect 18604 8041 18613 8075
rect 18613 8041 18647 8075
rect 18647 8041 18656 8075
rect 18604 8032 18656 8041
rect 19156 8032 19208 8084
rect 22008 8032 22060 8084
rect 25044 8075 25096 8084
rect 25044 8041 25053 8075
rect 25053 8041 25087 8075
rect 25087 8041 25096 8075
rect 25044 8032 25096 8041
rect 25596 8075 25648 8084
rect 25596 8041 25605 8075
rect 25605 8041 25639 8075
rect 25639 8041 25648 8075
rect 25596 8032 25648 8041
rect 18420 7964 18472 8016
rect 5172 7896 5224 7948
rect 7932 7896 7984 7948
rect 9956 7896 10008 7948
rect 5080 7828 5132 7880
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 7196 7828 7248 7880
rect 7656 7828 7708 7880
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 10692 7896 10744 7948
rect 11520 7896 11572 7948
rect 13176 7939 13228 7948
rect 13176 7905 13185 7939
rect 13185 7905 13219 7939
rect 13219 7905 13228 7939
rect 13176 7896 13228 7905
rect 13360 7896 13412 7948
rect 10784 7828 10836 7880
rect 11152 7828 11204 7880
rect 13820 7828 13872 7880
rect 15016 7871 15068 7880
rect 15016 7837 15025 7871
rect 15025 7837 15059 7871
rect 15059 7837 15068 7871
rect 15016 7828 15068 7837
rect 15108 7828 15160 7880
rect 15476 7828 15528 7880
rect 15660 7871 15712 7880
rect 15660 7837 15669 7871
rect 15669 7837 15703 7871
rect 15703 7837 15712 7871
rect 15660 7828 15712 7837
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 16948 7871 17000 7880
rect 16948 7837 16957 7871
rect 16957 7837 16991 7871
rect 16991 7837 17000 7871
rect 16948 7828 17000 7837
rect 18144 7896 18196 7948
rect 19800 7871 19852 7880
rect 19800 7837 19809 7871
rect 19809 7837 19843 7871
rect 19843 7837 19852 7871
rect 19800 7828 19852 7837
rect 25412 7964 25464 8016
rect 22376 7939 22428 7948
rect 22376 7905 22385 7939
rect 22385 7905 22419 7939
rect 22419 7905 22428 7939
rect 22376 7896 22428 7905
rect 4988 7760 5040 7812
rect 6736 7760 6788 7812
rect 7932 7803 7984 7812
rect 3608 7692 3660 7744
rect 4344 7735 4396 7744
rect 4344 7701 4353 7735
rect 4353 7701 4387 7735
rect 4387 7701 4396 7735
rect 4344 7692 4396 7701
rect 5540 7735 5592 7744
rect 5540 7701 5549 7735
rect 5549 7701 5583 7735
rect 5583 7701 5592 7735
rect 5540 7692 5592 7701
rect 7564 7692 7616 7744
rect 7932 7769 7941 7803
rect 7941 7769 7975 7803
rect 7975 7769 7984 7803
rect 7932 7760 7984 7769
rect 14096 7803 14148 7812
rect 14096 7769 14105 7803
rect 14105 7769 14139 7803
rect 14139 7769 14148 7803
rect 14096 7760 14148 7769
rect 16028 7760 16080 7812
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 9588 7735 9640 7744
rect 8392 7692 8444 7701
rect 9588 7701 9597 7735
rect 9597 7701 9631 7735
rect 9631 7701 9640 7735
rect 9588 7692 9640 7701
rect 10784 7692 10836 7744
rect 11428 7735 11480 7744
rect 11428 7701 11437 7735
rect 11437 7701 11471 7735
rect 11471 7701 11480 7735
rect 11428 7692 11480 7701
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 13084 7692 13136 7744
rect 14004 7692 14056 7744
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 15568 7692 15620 7744
rect 17408 7760 17460 7812
rect 18144 7803 18196 7812
rect 18144 7769 18153 7803
rect 18153 7769 18187 7803
rect 18187 7769 18196 7803
rect 18144 7760 18196 7769
rect 21916 7828 21968 7880
rect 22008 7828 22060 7880
rect 25136 7896 25188 7948
rect 23388 7828 23440 7880
rect 21272 7760 21324 7812
rect 21364 7760 21416 7812
rect 29184 7760 29236 7812
rect 20076 7692 20128 7744
rect 20812 7735 20864 7744
rect 20812 7701 20821 7735
rect 20821 7701 20855 7735
rect 20855 7701 20864 7735
rect 20812 7692 20864 7701
rect 21640 7735 21692 7744
rect 21640 7701 21649 7735
rect 21649 7701 21683 7735
rect 21683 7701 21692 7735
rect 21640 7692 21692 7701
rect 22100 7692 22152 7744
rect 23204 7692 23256 7744
rect 23756 7735 23808 7744
rect 23756 7701 23765 7735
rect 23765 7701 23799 7735
rect 23799 7701 23808 7735
rect 23756 7692 23808 7701
rect 24400 7735 24452 7744
rect 24400 7701 24409 7735
rect 24409 7701 24443 7735
rect 24443 7701 24452 7735
rect 24400 7692 24452 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 3608 7488 3660 7540
rect 3792 7488 3844 7540
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 2872 7352 2924 7404
rect 5080 7488 5132 7540
rect 8300 7488 8352 7540
rect 8852 7531 8904 7540
rect 8852 7497 8861 7531
rect 8861 7497 8895 7531
rect 8895 7497 8904 7531
rect 8852 7488 8904 7497
rect 9496 7488 9548 7540
rect 14464 7531 14516 7540
rect 10416 7463 10468 7472
rect 10416 7429 10425 7463
rect 10425 7429 10459 7463
rect 10459 7429 10468 7463
rect 10416 7420 10468 7429
rect 12716 7420 12768 7472
rect 13176 7420 13228 7472
rect 13360 7420 13412 7472
rect 14464 7497 14473 7531
rect 14473 7497 14507 7531
rect 14507 7497 14516 7531
rect 14464 7488 14516 7497
rect 14648 7420 14700 7472
rect 15936 7420 15988 7472
rect 16948 7420 17000 7472
rect 21180 7488 21232 7540
rect 21640 7488 21692 7540
rect 29552 7488 29604 7540
rect 17592 7420 17644 7472
rect 18420 7420 18472 7472
rect 18604 7420 18656 7472
rect 5540 7352 5592 7404
rect 6828 7352 6880 7404
rect 5264 7284 5316 7336
rect 8208 7352 8260 7404
rect 8300 7284 8352 7336
rect 8944 7352 8996 7404
rect 11520 7352 11572 7404
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 11888 7352 11940 7361
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 16488 7352 16540 7404
rect 19248 7420 19300 7472
rect 21548 7420 21600 7472
rect 7472 7216 7524 7268
rect 10784 7284 10836 7336
rect 11980 7327 12032 7336
rect 11980 7293 11989 7327
rect 11989 7293 12023 7327
rect 12023 7293 12032 7327
rect 11980 7284 12032 7293
rect 12256 7284 12308 7336
rect 12716 7284 12768 7336
rect 13820 7284 13872 7336
rect 16028 7284 16080 7336
rect 19432 7352 19484 7404
rect 20260 7352 20312 7404
rect 22008 7352 22060 7404
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 23756 7352 23808 7404
rect 32588 7352 32640 7404
rect 9496 7259 9548 7268
rect 9496 7225 9505 7259
rect 9505 7225 9539 7259
rect 9539 7225 9548 7259
rect 9496 7216 9548 7225
rect 11612 7216 11664 7268
rect 17960 7216 18012 7268
rect 20720 7284 20772 7336
rect 22376 7327 22428 7336
rect 22376 7293 22385 7327
rect 22385 7293 22419 7327
rect 22419 7293 22428 7327
rect 22376 7284 22428 7293
rect 24124 7284 24176 7336
rect 28356 7216 28408 7268
rect 6368 7148 6420 7200
rect 10140 7148 10192 7200
rect 11428 7148 11480 7200
rect 12256 7148 12308 7200
rect 12992 7148 13044 7200
rect 14464 7148 14516 7200
rect 15292 7148 15344 7200
rect 15752 7148 15804 7200
rect 19984 7148 20036 7200
rect 20628 7191 20680 7200
rect 20628 7157 20637 7191
rect 20637 7157 20671 7191
rect 20671 7157 20680 7191
rect 20628 7148 20680 7157
rect 24768 7191 24820 7200
rect 24768 7157 24777 7191
rect 24777 7157 24811 7191
rect 24811 7157 24820 7191
rect 24768 7148 24820 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3332 6944 3384 6996
rect 4804 6944 4856 6996
rect 6276 6944 6328 6996
rect 9128 6944 9180 6996
rect 9220 6944 9272 6996
rect 9772 6944 9824 6996
rect 10600 6944 10652 6996
rect 12440 6944 12492 6996
rect 13268 6944 13320 6996
rect 15200 6944 15252 6996
rect 17316 6944 17368 6996
rect 20444 6944 20496 6996
rect 22652 6944 22704 6996
rect 2872 6876 2924 6928
rect 7564 6876 7616 6928
rect 8576 6876 8628 6928
rect 8760 6876 8812 6928
rect 4436 6851 4488 6860
rect 4436 6817 4445 6851
rect 4445 6817 4479 6851
rect 4479 6817 4488 6851
rect 4436 6808 4488 6817
rect 5172 6851 5224 6860
rect 5172 6817 5181 6851
rect 5181 6817 5215 6851
rect 5215 6817 5224 6851
rect 5172 6808 5224 6817
rect 6092 6808 6144 6860
rect 7196 6808 7248 6860
rect 10968 6876 11020 6928
rect 1492 6740 1544 6792
rect 7104 6740 7156 6792
rect 7288 6783 7340 6792
rect 7288 6749 7297 6783
rect 7297 6749 7331 6783
rect 7331 6749 7340 6783
rect 7288 6740 7340 6749
rect 9404 6808 9456 6860
rect 9588 6851 9640 6860
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 10692 6808 10744 6860
rect 12072 6808 12124 6860
rect 12900 6808 12952 6860
rect 14648 6876 14700 6928
rect 17960 6876 18012 6928
rect 2780 6672 2832 6724
rect 2872 6672 2924 6724
rect 3700 6672 3752 6724
rect 6920 6672 6972 6724
rect 9956 6672 10008 6724
rect 10692 6715 10744 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 7472 6647 7524 6656
rect 7472 6613 7481 6647
rect 7481 6613 7515 6647
rect 7515 6613 7524 6647
rect 7472 6604 7524 6613
rect 7932 6604 7984 6656
rect 8300 6604 8352 6656
rect 8576 6604 8628 6656
rect 10232 6604 10284 6656
rect 10692 6681 10719 6715
rect 10719 6681 10744 6715
rect 10692 6672 10744 6681
rect 13084 6740 13136 6792
rect 12072 6672 12124 6724
rect 12440 6672 12492 6724
rect 11152 6604 11204 6656
rect 13268 6740 13320 6792
rect 13728 6808 13780 6860
rect 16304 6808 16356 6860
rect 15108 6740 15160 6792
rect 19708 6808 19760 6860
rect 20720 6876 20772 6928
rect 31024 6876 31076 6928
rect 21364 6808 21416 6860
rect 23020 6808 23072 6860
rect 24492 6808 24544 6860
rect 31116 6808 31168 6860
rect 42064 6808 42116 6860
rect 42708 6808 42760 6860
rect 18604 6740 18656 6792
rect 18236 6672 18288 6724
rect 19064 6740 19116 6792
rect 20628 6783 20680 6792
rect 19248 6672 19300 6724
rect 19524 6672 19576 6724
rect 13636 6604 13688 6656
rect 14096 6604 14148 6656
rect 14372 6604 14424 6656
rect 16672 6647 16724 6656
rect 16672 6613 16681 6647
rect 16681 6613 16715 6647
rect 16715 6613 16724 6647
rect 16672 6604 16724 6613
rect 17224 6647 17276 6656
rect 17224 6613 17233 6647
rect 17233 6613 17267 6647
rect 17267 6613 17276 6647
rect 17224 6604 17276 6613
rect 20260 6604 20312 6656
rect 20628 6749 20637 6783
rect 20637 6749 20671 6783
rect 20671 6749 20680 6783
rect 20628 6740 20680 6749
rect 21732 6647 21784 6656
rect 21732 6613 21741 6647
rect 21741 6613 21775 6647
rect 21775 6613 21784 6647
rect 21732 6604 21784 6613
rect 23940 6740 23992 6792
rect 24584 6783 24636 6792
rect 24584 6749 24593 6783
rect 24593 6749 24627 6783
rect 24627 6749 24636 6783
rect 24584 6740 24636 6749
rect 27896 6672 27948 6724
rect 23204 6604 23256 6656
rect 23480 6647 23532 6656
rect 23480 6613 23489 6647
rect 23489 6613 23523 6647
rect 23523 6613 23532 6647
rect 23480 6604 23532 6613
rect 23756 6604 23808 6656
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 25228 6604 25280 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2504 6400 2556 6452
rect 2964 6400 3016 6452
rect 3884 6443 3936 6452
rect 3884 6409 3893 6443
rect 3893 6409 3927 6443
rect 3927 6409 3936 6443
rect 3884 6400 3936 6409
rect 4068 6400 4120 6452
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 7196 6443 7248 6452
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 7932 6400 7984 6452
rect 8668 6400 8720 6452
rect 10048 6400 10100 6452
rect 2412 6332 2464 6384
rect 8576 6332 8628 6384
rect 11060 6400 11112 6452
rect 10508 6375 10560 6384
rect 10508 6341 10517 6375
rect 10517 6341 10551 6375
rect 10551 6341 10560 6375
rect 11888 6400 11940 6452
rect 14464 6400 14516 6452
rect 15292 6400 15344 6452
rect 15660 6400 15712 6452
rect 16120 6400 16172 6452
rect 17868 6400 17920 6452
rect 10508 6332 10560 6341
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 2780 6264 2832 6316
rect 7748 6264 7800 6316
rect 8116 6264 8168 6316
rect 9036 6264 9088 6316
rect 9772 6307 9824 6316
rect 4896 6196 4948 6248
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 10048 6264 10100 6316
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 10692 6264 10744 6316
rect 12348 6332 12400 6384
rect 11060 6264 11112 6316
rect 11612 6307 11664 6316
rect 11612 6273 11621 6307
rect 11621 6273 11655 6307
rect 11655 6273 11664 6307
rect 11612 6264 11664 6273
rect 14188 6332 14240 6384
rect 15108 6332 15160 6384
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 12900 6264 12952 6273
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 14648 6264 14700 6316
rect 20352 6400 20404 6452
rect 20628 6400 20680 6452
rect 31760 6400 31812 6452
rect 19708 6375 19760 6384
rect 19708 6341 19717 6375
rect 19717 6341 19751 6375
rect 19751 6341 19760 6375
rect 19708 6332 19760 6341
rect 19800 6332 19852 6384
rect 21916 6375 21968 6384
rect 21916 6341 21925 6375
rect 21925 6341 21959 6375
rect 21959 6341 21968 6375
rect 21916 6332 21968 6341
rect 23572 6375 23624 6384
rect 23572 6341 23581 6375
rect 23581 6341 23615 6375
rect 23615 6341 23624 6375
rect 23572 6332 23624 6341
rect 24032 6332 24084 6384
rect 2136 6128 2188 6180
rect 8024 6128 8076 6180
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 8116 6060 8168 6112
rect 10232 6060 10284 6112
rect 11060 6060 11112 6112
rect 15384 6239 15436 6248
rect 14188 6171 14240 6180
rect 14188 6137 14197 6171
rect 14197 6137 14231 6171
rect 14231 6137 14240 6171
rect 14188 6128 14240 6137
rect 13820 6060 13872 6112
rect 15384 6205 15393 6239
rect 15393 6205 15427 6239
rect 15427 6205 15436 6239
rect 15384 6196 15436 6205
rect 18604 6264 18656 6316
rect 19892 6264 19944 6316
rect 23296 6264 23348 6316
rect 14648 6128 14700 6180
rect 17868 6196 17920 6248
rect 19156 6196 19208 6248
rect 20076 6196 20128 6248
rect 21456 6196 21508 6248
rect 21640 6196 21692 6248
rect 15936 6128 15988 6180
rect 17592 6060 17644 6112
rect 19984 6128 20036 6180
rect 29828 6196 29880 6248
rect 24492 6128 24544 6180
rect 42800 6128 42852 6180
rect 20720 6060 20772 6112
rect 21088 6060 21140 6112
rect 22928 6103 22980 6112
rect 22928 6069 22937 6103
rect 22937 6069 22971 6103
rect 22971 6069 22980 6103
rect 22928 6060 22980 6069
rect 24584 6103 24636 6112
rect 24584 6069 24593 6103
rect 24593 6069 24627 6103
rect 24627 6069 24636 6103
rect 24584 6060 24636 6069
rect 25412 6060 25464 6112
rect 25688 6103 25740 6112
rect 25688 6069 25697 6103
rect 25697 6069 25731 6103
rect 25731 6069 25740 6103
rect 25688 6060 25740 6069
rect 26240 6103 26292 6112
rect 26240 6069 26249 6103
rect 26249 6069 26283 6103
rect 26283 6069 26292 6103
rect 26240 6060 26292 6069
rect 42984 6060 43036 6112
rect 43168 6060 43220 6112
rect 43812 6060 43864 6112
rect 44180 6103 44232 6112
rect 44180 6069 44189 6103
rect 44189 6069 44223 6103
rect 44223 6069 44232 6103
rect 44180 6060 44232 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1400 5899 1452 5908
rect 1400 5865 1409 5899
rect 1409 5865 1443 5899
rect 1443 5865 1452 5899
rect 1400 5856 1452 5865
rect 3056 5856 3108 5908
rect 3700 5856 3752 5908
rect 6460 5856 6512 5908
rect 8208 5856 8260 5908
rect 8760 5856 8812 5908
rect 9404 5856 9456 5908
rect 10600 5899 10652 5908
rect 10600 5865 10609 5899
rect 10609 5865 10643 5899
rect 10643 5865 10652 5899
rect 10600 5856 10652 5865
rect 11336 5856 11388 5908
rect 11796 5856 11848 5908
rect 12256 5899 12308 5908
rect 12256 5865 12265 5899
rect 12265 5865 12299 5899
rect 12299 5865 12308 5899
rect 12256 5856 12308 5865
rect 13544 5899 13596 5908
rect 2872 5788 2924 5840
rect 2964 5788 3016 5840
rect 1492 5652 1544 5704
rect 4068 5652 4120 5704
rect 5080 5584 5132 5636
rect 5724 5584 5776 5636
rect 7380 5584 7432 5636
rect 8024 5584 8076 5636
rect 11060 5788 11112 5840
rect 12072 5788 12124 5840
rect 8484 5652 8536 5704
rect 10232 5652 10284 5704
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 12348 5652 12400 5704
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 13544 5856 13596 5865
rect 15016 5856 15068 5908
rect 16396 5899 16448 5908
rect 16396 5865 16405 5899
rect 16405 5865 16439 5899
rect 16439 5865 16448 5899
rect 16396 5856 16448 5865
rect 16580 5856 16632 5908
rect 18328 5856 18380 5908
rect 18788 5856 18840 5908
rect 19248 5856 19300 5908
rect 19892 5899 19944 5908
rect 19892 5865 19901 5899
rect 19901 5865 19935 5899
rect 19935 5865 19944 5899
rect 19892 5856 19944 5865
rect 21180 5856 21232 5908
rect 23112 5899 23164 5908
rect 23112 5865 23121 5899
rect 23121 5865 23155 5899
rect 23155 5865 23164 5899
rect 23112 5856 23164 5865
rect 23296 5856 23348 5908
rect 27160 5899 27212 5908
rect 27160 5865 27169 5899
rect 27169 5865 27203 5899
rect 27203 5865 27212 5899
rect 27160 5856 27212 5865
rect 27804 5899 27856 5908
rect 27804 5865 27813 5899
rect 27813 5865 27847 5899
rect 27847 5865 27856 5899
rect 27804 5856 27856 5865
rect 27896 5856 27948 5908
rect 34520 5856 34572 5908
rect 13820 5788 13872 5840
rect 13176 5720 13228 5772
rect 15292 5720 15344 5772
rect 16028 5720 16080 5772
rect 18972 5788 19024 5840
rect 20352 5763 20404 5772
rect 15660 5652 15712 5704
rect 16764 5652 16816 5704
rect 17040 5652 17092 5704
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 20352 5729 20361 5763
rect 20361 5729 20395 5763
rect 20395 5729 20404 5763
rect 20352 5720 20404 5729
rect 23204 5720 23256 5772
rect 24584 5652 24636 5704
rect 42708 5652 42760 5704
rect 11612 5584 11664 5636
rect 14372 5627 14424 5636
rect 14372 5593 14381 5627
rect 14381 5593 14415 5627
rect 14415 5593 14424 5627
rect 14372 5584 14424 5593
rect 5632 5516 5684 5568
rect 5908 5559 5960 5568
rect 5908 5525 5917 5559
rect 5917 5525 5951 5559
rect 5951 5525 5960 5559
rect 5908 5516 5960 5525
rect 6092 5516 6144 5568
rect 7012 5516 7064 5568
rect 9772 5516 9824 5568
rect 11796 5559 11848 5568
rect 11796 5525 11805 5559
rect 11805 5525 11839 5559
rect 11839 5525 11848 5559
rect 11796 5516 11848 5525
rect 11888 5516 11940 5568
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 14464 5516 14516 5568
rect 15936 5559 15988 5568
rect 15936 5525 15945 5559
rect 15945 5525 15979 5559
rect 15979 5525 15988 5559
rect 15936 5516 15988 5525
rect 19340 5584 19392 5636
rect 22192 5584 22244 5636
rect 23020 5584 23072 5636
rect 18512 5516 18564 5568
rect 22008 5516 22060 5568
rect 22468 5516 22520 5568
rect 23664 5559 23716 5568
rect 23664 5525 23673 5559
rect 23673 5525 23707 5559
rect 23707 5525 23716 5559
rect 23664 5516 23716 5525
rect 24860 5516 24912 5568
rect 26148 5516 26200 5568
rect 30196 5516 30248 5568
rect 41696 5559 41748 5568
rect 41696 5525 41705 5559
rect 41705 5525 41739 5559
rect 41739 5525 41748 5559
rect 41696 5516 41748 5525
rect 42156 5516 42208 5568
rect 42340 5516 42392 5568
rect 42892 5559 42944 5568
rect 42892 5525 42901 5559
rect 42901 5525 42935 5559
rect 42935 5525 42944 5559
rect 42892 5516 42944 5525
rect 43536 5516 43588 5568
rect 45100 5516 45152 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1676 5312 1728 5364
rect 2136 5355 2188 5364
rect 2136 5321 2145 5355
rect 2145 5321 2179 5355
rect 2179 5321 2188 5355
rect 2136 5312 2188 5321
rect 5908 5312 5960 5364
rect 6368 5355 6420 5364
rect 6368 5321 6377 5355
rect 6377 5321 6411 5355
rect 6411 5321 6420 5355
rect 6368 5312 6420 5321
rect 8024 5355 8076 5364
rect 8024 5321 8033 5355
rect 8033 5321 8067 5355
rect 8067 5321 8076 5355
rect 8024 5312 8076 5321
rect 9864 5312 9916 5364
rect 10140 5312 10192 5364
rect 10784 5312 10836 5364
rect 848 5244 900 5296
rect 4068 5244 4120 5296
rect 5448 5244 5500 5296
rect 7012 5244 7064 5296
rect 10232 5244 10284 5296
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 8392 5176 8444 5228
rect 3976 5108 4028 5160
rect 8852 5108 8904 5160
rect 10784 5151 10836 5160
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 11796 5312 11848 5364
rect 12256 5244 12308 5296
rect 15660 5312 15712 5364
rect 16120 5355 16172 5364
rect 16120 5321 16129 5355
rect 16129 5321 16163 5355
rect 16163 5321 16172 5355
rect 16120 5312 16172 5321
rect 16856 5312 16908 5364
rect 17868 5355 17920 5364
rect 17868 5321 17877 5355
rect 17877 5321 17911 5355
rect 17911 5321 17920 5355
rect 17868 5312 17920 5321
rect 18144 5312 18196 5364
rect 18420 5312 18472 5364
rect 20628 5312 20680 5364
rect 23664 5312 23716 5364
rect 28080 5355 28132 5364
rect 28080 5321 28089 5355
rect 28089 5321 28123 5355
rect 28123 5321 28132 5355
rect 28080 5312 28132 5321
rect 28264 5312 28316 5364
rect 41420 5355 41472 5364
rect 41420 5321 41429 5355
rect 41429 5321 41463 5355
rect 41463 5321 41472 5355
rect 41420 5312 41472 5321
rect 16672 5244 16724 5296
rect 18328 5287 18380 5296
rect 18328 5253 18337 5287
rect 18337 5253 18371 5287
rect 18371 5253 18380 5287
rect 18328 5244 18380 5253
rect 19524 5287 19576 5296
rect 19524 5253 19533 5287
rect 19533 5253 19567 5287
rect 19567 5253 19576 5287
rect 19524 5244 19576 5253
rect 26608 5244 26660 5296
rect 42248 5244 42300 5296
rect 12716 5176 12768 5228
rect 14648 5219 14700 5228
rect 14188 5108 14240 5160
rect 14372 5151 14424 5160
rect 14372 5117 14381 5151
rect 14381 5117 14415 5151
rect 14415 5117 14424 5151
rect 14372 5108 14424 5117
rect 14648 5185 14657 5219
rect 14657 5185 14691 5219
rect 14691 5185 14700 5219
rect 14648 5176 14700 5185
rect 16304 5176 16356 5228
rect 22192 5176 22244 5228
rect 42892 5176 42944 5228
rect 45744 5176 45796 5228
rect 14924 5108 14976 5160
rect 15016 5108 15068 5160
rect 21916 5108 21968 5160
rect 23940 5108 23992 5160
rect 4528 5040 4580 5092
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 11060 5040 11112 5092
rect 11336 5040 11388 5092
rect 22928 5083 22980 5092
rect 22928 5049 22937 5083
rect 22937 5049 22971 5083
rect 22971 5049 22980 5083
rect 22928 5040 22980 5049
rect 23388 5040 23440 5092
rect 27896 5040 27948 5092
rect 5448 4972 5500 5024
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 5816 4972 5868 4981
rect 7104 4972 7156 5024
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 9036 5015 9088 5024
rect 9036 4981 9045 5015
rect 9045 4981 9079 5015
rect 9079 4981 9088 5015
rect 9036 4972 9088 4981
rect 13084 4972 13136 5024
rect 13728 4972 13780 5024
rect 15108 4972 15160 5024
rect 17040 4972 17092 5024
rect 17960 4972 18012 5024
rect 22284 4972 22336 5024
rect 24032 5015 24084 5024
rect 24032 4981 24041 5015
rect 24041 4981 24075 5015
rect 24075 4981 24084 5015
rect 24032 4972 24084 4981
rect 24676 4972 24728 5024
rect 25596 4972 25648 5024
rect 26332 5015 26384 5024
rect 26332 4981 26341 5015
rect 26341 4981 26375 5015
rect 26375 4981 26384 5015
rect 26332 4972 26384 4981
rect 26976 5015 27028 5024
rect 26976 4981 26985 5015
rect 26985 4981 27019 5015
rect 27019 4981 27028 5015
rect 26976 4972 27028 4981
rect 42616 5015 42668 5024
rect 42616 4981 42625 5015
rect 42625 4981 42659 5015
rect 42659 4981 42668 5015
rect 42616 4972 42668 4981
rect 43444 5015 43496 5024
rect 43444 4981 43453 5015
rect 43453 4981 43487 5015
rect 43487 4981 43496 5015
rect 43444 4972 43496 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1308 4768 1360 4820
rect 4620 4811 4672 4820
rect 4620 4777 4629 4811
rect 4629 4777 4663 4811
rect 4663 4777 4672 4811
rect 4620 4768 4672 4777
rect 8944 4768 8996 4820
rect 9128 4811 9180 4820
rect 9128 4777 9137 4811
rect 9137 4777 9171 4811
rect 9171 4777 9180 4811
rect 9128 4768 9180 4777
rect 9312 4768 9364 4820
rect 10508 4811 10560 4820
rect 10508 4777 10517 4811
rect 10517 4777 10551 4811
rect 10551 4777 10560 4811
rect 10508 4768 10560 4777
rect 11244 4811 11296 4820
rect 11244 4777 11253 4811
rect 11253 4777 11287 4811
rect 11287 4777 11296 4811
rect 11244 4768 11296 4777
rect 12624 4768 12676 4820
rect 14740 4811 14792 4820
rect 14740 4777 14749 4811
rect 14749 4777 14783 4811
rect 14783 4777 14792 4811
rect 14740 4768 14792 4777
rect 14924 4768 14976 4820
rect 16672 4811 16724 4820
rect 16672 4777 16681 4811
rect 16681 4777 16715 4811
rect 16715 4777 16724 4811
rect 16672 4768 16724 4777
rect 17316 4768 17368 4820
rect 18236 4768 18288 4820
rect 19984 4768 20036 4820
rect 23664 4811 23716 4820
rect 23664 4777 23673 4811
rect 23673 4777 23707 4811
rect 23707 4777 23716 4811
rect 23664 4768 23716 4777
rect 28816 4811 28868 4820
rect 28816 4777 28825 4811
rect 28825 4777 28859 4811
rect 28859 4777 28868 4811
rect 28816 4768 28868 4777
rect 35900 4811 35952 4820
rect 35900 4777 35909 4811
rect 35909 4777 35943 4811
rect 35943 4777 35952 4811
rect 37924 4811 37976 4820
rect 35900 4768 35952 4777
rect 37924 4777 37933 4811
rect 37933 4777 37967 4811
rect 37967 4777 37976 4811
rect 37924 4768 37976 4777
rect 40776 4811 40828 4820
rect 40776 4777 40785 4811
rect 40785 4777 40819 4811
rect 40819 4777 40828 4811
rect 40776 4768 40828 4777
rect 1584 4743 1636 4752
rect 1584 4709 1593 4743
rect 1593 4709 1627 4743
rect 1627 4709 1636 4743
rect 1584 4700 1636 4709
rect 10416 4700 10468 4752
rect 13452 4700 13504 4752
rect 13544 4700 13596 4752
rect 16212 4700 16264 4752
rect 22100 4743 22152 4752
rect 22100 4709 22109 4743
rect 22109 4709 22143 4743
rect 22143 4709 22152 4743
rect 22100 4700 22152 4709
rect 6552 4632 6604 4684
rect 6736 4632 6788 4684
rect 9496 4632 9548 4684
rect 13636 4632 13688 4684
rect 14740 4632 14792 4684
rect 19524 4632 19576 4684
rect 21272 4632 21324 4684
rect 28632 4700 28684 4752
rect 37096 4700 37148 4752
rect 42524 4700 42576 4752
rect 23572 4632 23624 4684
rect 1676 4564 1728 4616
rect 2044 4607 2096 4616
rect 2044 4573 2053 4607
rect 2053 4573 2087 4607
rect 2087 4573 2096 4607
rect 2044 4564 2096 4573
rect 5632 4564 5684 4616
rect 9036 4564 9088 4616
rect 14188 4564 14240 4616
rect 15200 4564 15252 4616
rect 3056 4496 3108 4548
rect 4712 4496 4764 4548
rect 12716 4496 12768 4548
rect 16396 4564 16448 4616
rect 20352 4564 20404 4616
rect 26976 4564 27028 4616
rect 39120 4607 39172 4616
rect 18512 4496 18564 4548
rect 5448 4428 5500 4480
rect 7932 4428 7984 4480
rect 13176 4428 13228 4480
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 14188 4428 14240 4437
rect 19984 4428 20036 4480
rect 21456 4471 21508 4480
rect 21456 4437 21465 4471
rect 21465 4437 21499 4471
rect 21499 4437 21508 4471
rect 21456 4428 21508 4437
rect 21548 4428 21600 4480
rect 24124 4496 24176 4548
rect 39120 4573 39129 4607
rect 39129 4573 39163 4607
rect 39163 4573 39172 4607
rect 39120 4564 39172 4573
rect 43168 4607 43220 4616
rect 43168 4573 43177 4607
rect 43177 4573 43211 4607
rect 43211 4573 43220 4607
rect 43168 4564 43220 4573
rect 27896 4496 27948 4548
rect 23112 4471 23164 4480
rect 23112 4437 23121 4471
rect 23121 4437 23155 4471
rect 23155 4437 23164 4471
rect 23112 4428 23164 4437
rect 24952 4471 25004 4480
rect 24952 4437 24961 4471
rect 24961 4437 24995 4471
rect 24995 4437 25004 4471
rect 24952 4428 25004 4437
rect 25044 4428 25096 4480
rect 26424 4428 26476 4480
rect 26608 4471 26660 4480
rect 26608 4437 26617 4471
rect 26617 4437 26651 4471
rect 26651 4437 26660 4471
rect 26608 4428 26660 4437
rect 27252 4471 27304 4480
rect 27252 4437 27261 4471
rect 27261 4437 27295 4471
rect 27295 4437 27304 4471
rect 27252 4428 27304 4437
rect 27712 4471 27764 4480
rect 27712 4437 27721 4471
rect 27721 4437 27755 4471
rect 27755 4437 27764 4471
rect 27712 4428 27764 4437
rect 33508 4428 33560 4480
rect 34796 4471 34848 4480
rect 34796 4437 34805 4471
rect 34805 4437 34839 4471
rect 34839 4437 34848 4471
rect 34796 4428 34848 4437
rect 35348 4471 35400 4480
rect 35348 4437 35357 4471
rect 35357 4437 35391 4471
rect 35391 4437 35400 4471
rect 35348 4428 35400 4437
rect 42984 4496 43036 4548
rect 44180 4496 44232 4548
rect 44824 4496 44876 4548
rect 36636 4428 36688 4480
rect 37280 4471 37332 4480
rect 37280 4437 37289 4471
rect 37289 4437 37323 4471
rect 37323 4437 37332 4471
rect 37280 4428 37332 4437
rect 38660 4471 38712 4480
rect 38660 4437 38669 4471
rect 38669 4437 38703 4471
rect 38703 4437 38712 4471
rect 38660 4428 38712 4437
rect 39856 4471 39908 4480
rect 39856 4437 39865 4471
rect 39865 4437 39899 4471
rect 39899 4437 39908 4471
rect 39856 4428 39908 4437
rect 41512 4428 41564 4480
rect 43168 4428 43220 4480
rect 43352 4471 43404 4480
rect 43352 4437 43361 4471
rect 43361 4437 43395 4471
rect 43395 4437 43404 4471
rect 43352 4428 43404 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 5816 4267 5868 4276
rect 5816 4233 5825 4267
rect 5825 4233 5859 4267
rect 5859 4233 5868 4267
rect 5816 4224 5868 4233
rect 9496 4267 9548 4276
rect 9496 4233 9505 4267
rect 9505 4233 9539 4267
rect 9539 4233 9548 4267
rect 9496 4224 9548 4233
rect 9680 4224 9732 4276
rect 21456 4224 21508 4276
rect 43536 4224 43588 4276
rect 1400 4156 1452 4208
rect 10416 4156 10468 4208
rect 10692 4199 10744 4208
rect 10692 4165 10701 4199
rect 10701 4165 10735 4199
rect 10735 4165 10744 4199
rect 10692 4156 10744 4165
rect 11428 4156 11480 4208
rect 11612 4199 11664 4208
rect 11612 4165 11621 4199
rect 11621 4165 11655 4199
rect 11655 4165 11664 4199
rect 11612 4156 11664 4165
rect 13360 4156 13412 4208
rect 14188 4156 14240 4208
rect 3884 4088 3936 4140
rect 7380 4088 7432 4140
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 8024 4088 8076 4140
rect 7932 4020 7984 4072
rect 1308 3952 1360 4004
rect 8484 3952 8536 4004
rect 9220 3952 9272 4004
rect 112 3884 164 3936
rect 1952 3884 2004 3936
rect 3240 3884 3292 3936
rect 5080 3884 5132 3936
rect 5724 3884 5776 3936
rect 6736 3927 6788 3936
rect 6736 3893 6745 3927
rect 6745 3893 6779 3927
rect 6779 3893 6788 3927
rect 6736 3884 6788 3893
rect 12808 4088 12860 4140
rect 14280 4088 14332 4140
rect 11428 4020 11480 4072
rect 15844 4088 15896 4140
rect 16580 4088 16632 4140
rect 17408 4131 17460 4140
rect 15384 4063 15436 4072
rect 12164 3995 12216 4004
rect 12164 3961 12173 3995
rect 12173 3961 12207 3995
rect 12207 3961 12216 3995
rect 12164 3952 12216 3961
rect 13544 3952 13596 4004
rect 15384 4029 15393 4063
rect 15393 4029 15427 4063
rect 15427 4029 15436 4063
rect 15384 4020 15436 4029
rect 17408 4097 17417 4131
rect 17417 4097 17451 4131
rect 17451 4097 17460 4131
rect 17408 4088 17460 4097
rect 18236 4088 18288 4140
rect 18328 4088 18380 4140
rect 18512 4088 18564 4140
rect 17592 4020 17644 4072
rect 14372 3952 14424 4004
rect 22744 4156 22796 4208
rect 25136 4156 25188 4208
rect 43812 4156 43864 4208
rect 45468 4156 45520 4208
rect 19156 4020 19208 4072
rect 21640 4088 21692 4140
rect 22376 4088 22428 4140
rect 27988 4088 28040 4140
rect 41696 4088 41748 4140
rect 43260 4088 43312 4140
rect 43996 4088 44048 4140
rect 19340 3995 19392 4004
rect 19340 3961 19349 3995
rect 19349 3961 19383 3995
rect 19383 3961 19392 3995
rect 19340 3952 19392 3961
rect 20260 3952 20312 4004
rect 24124 3952 24176 4004
rect 33048 4020 33100 4072
rect 36912 4020 36964 4072
rect 37372 3952 37424 4004
rect 44456 3952 44508 4004
rect 13820 3884 13872 3936
rect 14096 3884 14148 3936
rect 15292 3884 15344 3936
rect 19248 3884 19300 3936
rect 20444 3884 20496 3936
rect 21088 3927 21140 3936
rect 21088 3893 21097 3927
rect 21097 3893 21131 3927
rect 21131 3893 21140 3927
rect 21088 3884 21140 3893
rect 22928 3927 22980 3936
rect 22928 3893 22937 3927
rect 22937 3893 22971 3927
rect 22971 3893 22980 3927
rect 22928 3884 22980 3893
rect 23940 3884 23992 3936
rect 24584 3927 24636 3936
rect 24584 3893 24593 3927
rect 24593 3893 24627 3927
rect 24627 3893 24636 3927
rect 24584 3884 24636 3893
rect 25136 3927 25188 3936
rect 25136 3893 25145 3927
rect 25145 3893 25179 3927
rect 25179 3893 25188 3927
rect 25136 3884 25188 3893
rect 25320 3884 25372 3936
rect 27160 3884 27212 3936
rect 27988 3927 28040 3936
rect 27988 3893 27997 3927
rect 27997 3893 28031 3927
rect 28031 3893 28040 3927
rect 27988 3884 28040 3893
rect 28724 3927 28776 3936
rect 28724 3893 28733 3927
rect 28733 3893 28767 3927
rect 28767 3893 28776 3927
rect 28724 3884 28776 3893
rect 29368 3927 29420 3936
rect 29368 3893 29377 3927
rect 29377 3893 29411 3927
rect 29411 3893 29420 3927
rect 29368 3884 29420 3893
rect 30288 3884 30340 3936
rect 30748 3927 30800 3936
rect 30748 3893 30757 3927
rect 30757 3893 30791 3927
rect 30791 3893 30800 3927
rect 30748 3884 30800 3893
rect 31208 3927 31260 3936
rect 31208 3893 31217 3927
rect 31217 3893 31251 3927
rect 31251 3893 31260 3927
rect 31208 3884 31260 3893
rect 31668 3884 31720 3936
rect 33324 3884 33376 3936
rect 34612 3927 34664 3936
rect 34612 3893 34621 3927
rect 34621 3893 34655 3927
rect 34655 3893 34664 3927
rect 34612 3884 34664 3893
rect 35440 3884 35492 3936
rect 36084 3927 36136 3936
rect 36084 3893 36093 3927
rect 36093 3893 36127 3927
rect 36127 3893 36136 3927
rect 36084 3884 36136 3893
rect 36268 3884 36320 3936
rect 37188 3884 37240 3936
rect 38844 3927 38896 3936
rect 38844 3893 38853 3927
rect 38853 3893 38887 3927
rect 38887 3893 38896 3927
rect 38844 3884 38896 3893
rect 39764 3927 39816 3936
rect 39764 3893 39773 3927
rect 39773 3893 39807 3927
rect 39807 3893 39816 3927
rect 39764 3884 39816 3893
rect 39948 3884 40000 3936
rect 40408 3884 40460 3936
rect 44180 3884 44232 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 6644 3723 6696 3732
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 9496 3723 9548 3732
rect 9496 3689 9505 3723
rect 9505 3689 9539 3723
rect 9539 3689 9548 3723
rect 9496 3680 9548 3689
rect 9956 3723 10008 3732
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 10876 3680 10928 3732
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 11520 3680 11572 3732
rect 13360 3723 13412 3732
rect 13360 3689 13369 3723
rect 13369 3689 13403 3723
rect 13403 3689 13412 3723
rect 13360 3680 13412 3689
rect 13912 3680 13964 3732
rect 14648 3680 14700 3732
rect 18880 3680 18932 3732
rect 20168 3680 20220 3732
rect 20996 3680 21048 3732
rect 21364 3680 21416 3732
rect 664 3612 716 3664
rect 3976 3655 4028 3664
rect 3976 3621 3985 3655
rect 3985 3621 4019 3655
rect 4019 3621 4028 3655
rect 3976 3612 4028 3621
rect 10048 3612 10100 3664
rect 11704 3612 11756 3664
rect 14740 3655 14792 3664
rect 14740 3621 14749 3655
rect 14749 3621 14783 3655
rect 14783 3621 14792 3655
rect 14740 3612 14792 3621
rect 14832 3612 14884 3664
rect 7472 3544 7524 3596
rect 7656 3587 7708 3596
rect 7656 3553 7665 3587
rect 7665 3553 7699 3587
rect 7699 3553 7708 3587
rect 7656 3544 7708 3553
rect 8300 3544 8352 3596
rect 15016 3544 15068 3596
rect 1032 3476 1084 3528
rect 2964 3476 3016 3528
rect 4160 3476 4212 3528
rect 5724 3476 5776 3528
rect 6092 3476 6144 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 11244 3519 11296 3528
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 5172 3408 5224 3460
rect 11704 3408 11756 3460
rect 12624 3408 12676 3460
rect 13636 3476 13688 3528
rect 14372 3476 14424 3528
rect 15660 3476 15712 3528
rect 20444 3612 20496 3664
rect 20720 3612 20772 3664
rect 27528 3680 27580 3732
rect 37464 3723 37516 3732
rect 22652 3612 22704 3664
rect 27344 3612 27396 3664
rect 27436 3612 27488 3664
rect 30104 3612 30156 3664
rect 16488 3476 16540 3528
rect 19984 3544 20036 3596
rect 20076 3544 20128 3596
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 18972 3476 19024 3528
rect 20352 3519 20404 3528
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 20352 3476 20404 3485
rect 21272 3476 21324 3528
rect 22100 3476 22152 3528
rect 22744 3476 22796 3528
rect 17960 3408 18012 3460
rect 4620 3383 4672 3392
rect 4620 3349 4629 3383
rect 4629 3349 4663 3383
rect 4663 3349 4672 3383
rect 4620 3340 4672 3349
rect 16580 3340 16632 3392
rect 17868 3340 17920 3392
rect 19340 3408 19392 3460
rect 19432 3408 19484 3460
rect 18604 3340 18656 3392
rect 23572 3544 23624 3596
rect 25688 3544 25740 3596
rect 28356 3544 28408 3596
rect 37464 3689 37473 3723
rect 37473 3689 37507 3723
rect 37507 3689 37516 3723
rect 37464 3680 37516 3689
rect 43076 3612 43128 3664
rect 43904 3655 43956 3664
rect 43904 3621 43913 3655
rect 43913 3621 43947 3655
rect 43947 3621 43956 3655
rect 43904 3612 43956 3621
rect 23388 3519 23440 3528
rect 23388 3485 23397 3519
rect 23397 3485 23431 3519
rect 23431 3485 23440 3519
rect 23388 3476 23440 3485
rect 24032 3476 24084 3528
rect 24952 3476 25004 3528
rect 25228 3519 25280 3528
rect 25228 3485 25237 3519
rect 25237 3485 25271 3519
rect 25271 3485 25280 3519
rect 25228 3476 25280 3485
rect 27620 3476 27672 3528
rect 27988 3519 28040 3528
rect 27988 3485 27997 3519
rect 27997 3485 28031 3519
rect 28031 3485 28040 3519
rect 27988 3476 28040 3485
rect 28816 3476 28868 3528
rect 29552 3519 29604 3528
rect 29552 3485 29561 3519
rect 29561 3485 29595 3519
rect 29595 3485 29604 3519
rect 29552 3476 29604 3485
rect 43996 3544 44048 3596
rect 31024 3519 31076 3528
rect 31024 3485 31033 3519
rect 31033 3485 31067 3519
rect 31067 3485 31076 3519
rect 31024 3476 31076 3485
rect 31944 3519 31996 3528
rect 31944 3485 31953 3519
rect 31953 3485 31987 3519
rect 31987 3485 31996 3519
rect 31944 3476 31996 3485
rect 32956 3519 33008 3528
rect 32956 3485 32965 3519
rect 32965 3485 32999 3519
rect 32999 3485 33008 3519
rect 32956 3476 33008 3485
rect 33876 3519 33928 3528
rect 33876 3485 33885 3519
rect 33885 3485 33919 3519
rect 33919 3485 33928 3519
rect 33876 3476 33928 3485
rect 34520 3476 34572 3528
rect 35900 3476 35952 3528
rect 36636 3519 36688 3528
rect 36636 3485 36645 3519
rect 36645 3485 36679 3519
rect 36679 3485 36688 3519
rect 36636 3476 36688 3485
rect 37924 3476 37976 3528
rect 39120 3519 39172 3528
rect 39120 3485 39129 3519
rect 39129 3485 39163 3519
rect 39163 3485 39172 3519
rect 39120 3476 39172 3485
rect 39856 3519 39908 3528
rect 39856 3485 39865 3519
rect 39865 3485 39899 3519
rect 39899 3485 39908 3519
rect 39856 3476 39908 3485
rect 41420 3476 41472 3528
rect 42340 3519 42392 3528
rect 42340 3485 42349 3519
rect 42349 3485 42383 3519
rect 42383 3485 42392 3519
rect 42340 3476 42392 3485
rect 27068 3451 27120 3460
rect 27068 3417 27077 3451
rect 27077 3417 27111 3451
rect 27111 3417 27120 3451
rect 27068 3408 27120 3417
rect 27344 3408 27396 3460
rect 32404 3408 32456 3460
rect 37280 3408 37332 3460
rect 42984 3408 43036 3460
rect 44456 3408 44508 3460
rect 24584 3340 24636 3392
rect 24860 3340 24912 3392
rect 25688 3383 25740 3392
rect 25688 3349 25697 3383
rect 25697 3349 25731 3383
rect 25731 3349 25740 3383
rect 25688 3340 25740 3349
rect 26240 3340 26292 3392
rect 28172 3340 28224 3392
rect 29092 3340 29144 3392
rect 30012 3340 30064 3392
rect 30932 3340 30984 3392
rect 31852 3340 31904 3392
rect 32864 3340 32916 3392
rect 33784 3340 33836 3392
rect 34704 3340 34756 3392
rect 35624 3340 35676 3392
rect 36636 3340 36688 3392
rect 37648 3340 37700 3392
rect 38476 3340 38528 3392
rect 39488 3340 39540 3392
rect 40684 3383 40736 3392
rect 40684 3349 40693 3383
rect 40693 3349 40727 3383
rect 40727 3349 40736 3383
rect 40684 3340 40736 3349
rect 41328 3340 41380 3392
rect 42248 3340 42300 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4068 3136 4120 3188
rect 11888 3136 11940 3188
rect 12256 3136 12308 3188
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 14556 3136 14608 3188
rect 17776 3179 17828 3188
rect 3424 3000 3476 3052
rect 388 2932 440 2984
rect 2320 2932 2372 2984
rect 4712 3068 4764 3120
rect 4068 3000 4120 3052
rect 4896 3000 4948 3052
rect 5448 3000 5500 3052
rect 2596 2864 2648 2916
rect 4712 2932 4764 2984
rect 5540 2864 5592 2916
rect 13084 3068 13136 3120
rect 6736 3000 6788 3052
rect 8576 3043 8628 3052
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 8944 3000 8996 3052
rect 9680 3000 9732 3052
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 12256 3043 12308 3052
rect 8852 2975 8904 2984
rect 6920 2864 6972 2916
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 8852 2932 8904 2941
rect 9864 2932 9916 2984
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 12348 2932 12400 2984
rect 13268 3000 13320 3052
rect 14280 3000 14332 3052
rect 14648 3000 14700 3052
rect 16396 3068 16448 3120
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 17960 3136 18012 3188
rect 16120 3000 16172 3052
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 20536 3136 20588 3188
rect 20904 3136 20956 3188
rect 21824 3136 21876 3188
rect 22836 3179 22888 3188
rect 22836 3145 22845 3179
rect 22845 3145 22879 3179
rect 22879 3145 22888 3179
rect 22836 3136 22888 3145
rect 23112 3136 23164 3188
rect 23296 3136 23348 3188
rect 23848 3136 23900 3188
rect 24216 3136 24268 3188
rect 26884 3136 26936 3188
rect 27068 3179 27120 3188
rect 27068 3145 27077 3179
rect 27077 3145 27111 3179
rect 27111 3145 27120 3179
rect 27068 3136 27120 3145
rect 27528 3136 27580 3188
rect 32772 3136 32824 3188
rect 35532 3179 35584 3188
rect 35532 3145 35541 3179
rect 35541 3145 35575 3179
rect 35575 3145 35584 3179
rect 35532 3136 35584 3145
rect 37372 3179 37424 3188
rect 37372 3145 37381 3179
rect 37381 3145 37415 3179
rect 37415 3145 37424 3179
rect 37372 3136 37424 3145
rect 43996 3179 44048 3188
rect 43996 3145 44005 3179
rect 44005 3145 44039 3179
rect 44039 3145 44048 3179
rect 43996 3136 44048 3145
rect 20720 3068 20772 3120
rect 19064 3043 19116 3052
rect 13820 2932 13872 2984
rect 17040 2932 17092 2984
rect 19064 3009 19073 3043
rect 19073 3009 19107 3043
rect 19107 3009 19116 3043
rect 19064 3000 19116 3009
rect 19984 3043 20036 3052
rect 19984 3009 19993 3043
rect 19993 3009 20027 3043
rect 20027 3009 20036 3043
rect 19984 3000 20036 3009
rect 20628 3000 20680 3052
rect 20904 3000 20956 3052
rect 22376 3068 22428 3120
rect 21824 3000 21876 3052
rect 22192 3000 22244 3052
rect 22744 3000 22796 3052
rect 23020 3043 23072 3052
rect 23020 3009 23029 3043
rect 23029 3009 23063 3043
rect 23063 3009 23072 3043
rect 23020 3000 23072 3009
rect 23664 3000 23716 3052
rect 25044 3068 25096 3120
rect 25872 3068 25924 3120
rect 26148 3068 26200 3120
rect 27344 3068 27396 3120
rect 27436 3068 27488 3120
rect 27712 3068 27764 3120
rect 28448 3068 28500 3120
rect 29644 3068 29696 3120
rect 30288 3111 30340 3120
rect 30288 3077 30297 3111
rect 30297 3077 30331 3111
rect 30331 3077 30340 3111
rect 30288 3068 30340 3077
rect 30656 3068 30708 3120
rect 31208 3068 31260 3120
rect 32496 3068 32548 3120
rect 33048 3068 33100 3120
rect 34520 3068 34572 3120
rect 35992 3068 36044 3120
rect 37188 3068 37240 3120
rect 38016 3111 38068 3120
rect 38016 3077 38025 3111
rect 38025 3077 38059 3111
rect 38059 3077 38068 3111
rect 38016 3068 38068 3077
rect 39396 3068 39448 3120
rect 40224 3111 40276 3120
rect 40224 3077 40233 3111
rect 40233 3077 40267 3111
rect 40267 3077 40276 3111
rect 40224 3068 40276 3077
rect 42800 3111 42852 3120
rect 42800 3077 42809 3111
rect 42809 3077 42843 3111
rect 42843 3077 42852 3111
rect 42800 3068 42852 3077
rect 43168 3068 43220 3120
rect 43536 3068 43588 3120
rect 24584 2932 24636 2984
rect 24676 2932 24728 2984
rect 25780 3000 25832 3052
rect 26700 3000 26752 3052
rect 26792 2932 26844 2984
rect 27344 2932 27396 2984
rect 28724 3000 28776 3052
rect 28908 3000 28960 3052
rect 30196 3000 30248 3052
rect 31668 3000 31720 3052
rect 33508 3000 33560 3052
rect 34428 3000 34480 3052
rect 34796 3000 34848 3052
rect 35348 3000 35400 3052
rect 36268 3000 36320 3052
rect 36912 2932 36964 2984
rect 38292 3000 38344 3052
rect 38660 3000 38712 3052
rect 39120 3000 39172 3052
rect 39948 3000 40000 3052
rect 40040 3000 40092 3052
rect 40408 3043 40460 3052
rect 40408 3009 40417 3043
rect 40417 3009 40451 3043
rect 40451 3009 40460 3043
rect 40408 3000 40460 3009
rect 40776 3000 40828 3052
rect 41972 3000 42024 3052
rect 42616 3000 42668 3052
rect 9588 2796 9640 2848
rect 11060 2796 11112 2848
rect 11888 2796 11940 2848
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12440 2796 12492 2805
rect 12716 2864 12768 2916
rect 15752 2864 15804 2916
rect 18052 2864 18104 2916
rect 16672 2796 16724 2848
rect 16764 2796 16816 2848
rect 17592 2796 17644 2848
rect 19892 2864 19944 2916
rect 22560 2864 22612 2916
rect 33232 2907 33284 2916
rect 18696 2796 18748 2848
rect 25228 2796 25280 2848
rect 25780 2796 25832 2848
rect 26424 2796 26476 2848
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 33232 2873 33241 2907
rect 33241 2873 33275 2907
rect 33275 2873 33284 2907
rect 33232 2864 33284 2873
rect 34152 2864 34204 2916
rect 40408 2796 40460 2848
rect 41696 2796 41748 2848
rect 42800 2796 42852 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 5264 2592 5316 2644
rect 8300 2592 8352 2644
rect 8576 2592 8628 2644
rect 9496 2592 9548 2644
rect 19892 2592 19944 2644
rect 33692 2592 33744 2644
rect 2688 2567 2740 2576
rect 2688 2533 2697 2567
rect 2697 2533 2731 2567
rect 2731 2533 2740 2567
rect 2688 2524 2740 2533
rect 8116 2524 8168 2576
rect 11152 2524 11204 2576
rect 17776 2567 17828 2576
rect 17776 2533 17785 2567
rect 17785 2533 17819 2567
rect 17819 2533 17828 2567
rect 17776 2524 17828 2533
rect 5356 2456 5408 2508
rect 2780 2388 2832 2440
rect 4436 2388 4488 2440
rect 5080 2388 5132 2440
rect 6828 2388 6880 2440
rect 7012 2431 7064 2440
rect 7012 2397 7021 2431
rect 7021 2397 7055 2431
rect 7055 2397 7064 2431
rect 7012 2388 7064 2397
rect 2872 2363 2924 2372
rect 2872 2329 2881 2363
rect 2881 2329 2915 2363
rect 2915 2329 2924 2363
rect 2872 2320 2924 2329
rect 4068 2320 4120 2372
rect 9588 2456 9640 2508
rect 10140 2499 10192 2508
rect 10140 2465 10149 2499
rect 10149 2465 10183 2499
rect 10183 2465 10192 2499
rect 10140 2456 10192 2465
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 8484 2388 8536 2440
rect 9496 2388 9548 2440
rect 11428 2456 11480 2508
rect 11888 2456 11940 2508
rect 17500 2456 17552 2508
rect 12440 2388 12492 2440
rect 12992 2388 13044 2440
rect 14004 2388 14056 2440
rect 6368 2252 6420 2304
rect 15568 2388 15620 2440
rect 15476 2320 15528 2372
rect 10140 2252 10192 2304
rect 12072 2252 12124 2304
rect 12992 2252 13044 2304
rect 13912 2252 13964 2304
rect 14832 2252 14884 2304
rect 15200 2252 15252 2304
rect 15936 2388 15988 2440
rect 17224 2388 17276 2440
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 25964 2499 26016 2508
rect 25964 2465 25973 2499
rect 25973 2465 26007 2499
rect 26007 2465 26016 2499
rect 25964 2456 26016 2465
rect 20812 2388 20864 2440
rect 21732 2388 21784 2440
rect 23480 2388 23532 2440
rect 23756 2431 23808 2440
rect 23756 2397 23765 2431
rect 23765 2397 23799 2431
rect 23799 2397 23808 2431
rect 23756 2388 23808 2397
rect 24308 2388 24360 2440
rect 25596 2388 25648 2440
rect 25780 2431 25832 2440
rect 25780 2397 25789 2431
rect 25789 2397 25823 2431
rect 25823 2397 25832 2431
rect 25780 2388 25832 2397
rect 17408 2320 17460 2372
rect 21088 2320 21140 2372
rect 15844 2295 15896 2304
rect 15844 2261 15853 2295
rect 15853 2261 15887 2295
rect 15887 2261 15896 2295
rect 15844 2252 15896 2261
rect 15936 2252 15988 2304
rect 17776 2252 17828 2304
rect 19432 2252 19484 2304
rect 20536 2252 20588 2304
rect 21456 2252 21508 2304
rect 22468 2252 22520 2304
rect 23388 2252 23440 2304
rect 24308 2252 24360 2304
rect 25136 2295 25188 2304
rect 25136 2261 25145 2295
rect 25145 2261 25179 2295
rect 25179 2261 25188 2295
rect 25136 2252 25188 2261
rect 27344 2524 27396 2576
rect 28540 2524 28592 2576
rect 32680 2524 32732 2576
rect 35072 2524 35124 2576
rect 37096 2524 37148 2576
rect 27528 2456 27580 2508
rect 32220 2456 32272 2508
rect 33324 2456 33376 2508
rect 28356 2388 28408 2440
rect 29368 2388 29420 2440
rect 30380 2388 30432 2440
rect 34980 2456 35032 2508
rect 34060 2388 34112 2440
rect 26516 2320 26568 2372
rect 27252 2320 27304 2372
rect 29920 2320 29972 2372
rect 30288 2320 30340 2372
rect 30748 2320 30800 2372
rect 31300 2320 31352 2372
rect 28264 2252 28316 2304
rect 33140 2320 33192 2372
rect 34612 2320 34664 2372
rect 35072 2388 35124 2440
rect 36084 2388 36136 2440
rect 39764 2388 39816 2440
rect 42800 2388 42852 2440
rect 35440 2320 35492 2372
rect 37832 2320 37884 2372
rect 38844 2320 38896 2372
rect 40684 2320 40736 2372
rect 41052 2320 41104 2372
rect 41512 2320 41564 2372
rect 42616 2320 42668 2372
rect 43444 2320 43496 2372
rect 35532 2295 35584 2304
rect 35532 2261 35541 2295
rect 35541 2261 35575 2295
rect 35575 2261 35584 2295
rect 35532 2252 35584 2261
rect 40040 2295 40092 2304
rect 40040 2261 40049 2295
rect 40049 2261 40083 2295
rect 40083 2261 40092 2295
rect 40040 2252 40092 2261
rect 40132 2252 40184 2304
rect 41604 2295 41656 2304
rect 41604 2261 41613 2295
rect 41613 2261 41647 2295
rect 41647 2261 41656 2295
rect 41604 2252 41656 2261
rect 42892 2295 42944 2304
rect 42892 2261 42901 2295
rect 42901 2261 42935 2295
rect 42935 2261 42944 2295
rect 42892 2252 42944 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 7656 2048 7708 2100
rect 17316 2048 17368 2100
rect 20720 2048 20772 2100
rect 41604 2048 41656 2100
rect 5540 1980 5592 2032
rect 25688 1980 25740 2032
rect 31116 1980 31168 2032
rect 34980 1980 35032 2032
rect 5724 1912 5776 1964
rect 22928 1912 22980 1964
rect 27068 1912 27120 1964
rect 40040 1912 40092 1964
rect 6368 1844 6420 1896
rect 6828 1844 6880 1896
rect 25136 1844 25188 1896
rect 2872 1776 2924 1828
rect 11612 1776 11664 1828
rect 13820 1776 13872 1828
rect 24492 1776 24544 1828
rect 8116 1708 8168 1760
rect 11980 1708 12032 1760
rect 18420 1708 18472 1760
rect 35532 1708 35584 1760
rect 8024 1640 8076 1692
rect 23940 1640 23992 1692
rect 7012 1572 7064 1624
rect 7932 1572 7984 1624
rect 22008 1572 22060 1624
rect 17868 1504 17920 1556
rect 20260 1504 20312 1556
rect 11796 1368 11848 1420
rect 20444 1368 20496 1420
rect 20 1300 72 1352
rect 940 1300 992 1352
rect 15384 1300 15436 1352
rect 27528 1300 27580 1352
rect 17316 1232 17368 1284
rect 20168 1232 20220 1284
rect 20444 1232 20496 1284
rect 22192 1232 22244 1284
rect 6920 1164 6972 1216
rect 24124 1164 24176 1216
rect 10784 1096 10836 1148
rect 11244 1096 11296 1148
rect 17960 1096 18012 1148
rect 18144 1096 18196 1148
rect 25412 1096 25464 1148
rect 7288 1028 7340 1080
rect 8852 1028 8904 1080
rect 22284 1028 22336 1080
rect 2780 960 2832 1012
rect 22560 960 22612 1012
rect 7564 892 7616 944
rect 5540 824 5592 876
rect 16304 824 16356 876
rect 17960 892 18012 944
rect 23572 892 23624 944
rect 24768 824 24820 876
rect 3792 756 3844 808
rect 15108 756 15160 808
rect 4712 688 4764 740
rect 16856 688 16908 740
rect 9404 348 9456 400
rect 17868 348 17920 400
rect 13360 280 13412 332
rect 23204 280 23256 332
rect 16212 212 16264 264
rect 26332 212 26384 264
rect 11612 144 11664 196
rect 12256 144 12308 196
rect 25504 144 25556 196
rect 14372 76 14424 128
rect 26608 76 26660 128
rect 10692 8 10744 60
rect 25320 8 25372 60
<< metal2 >>
rect 202 39200 258 40000
rect 570 39200 626 40000
rect 938 39200 994 40000
rect 1398 39200 1454 40000
rect 1766 39200 1822 40000
rect 2134 39200 2190 40000
rect 2594 39200 2650 40000
rect 2962 39200 3018 40000
rect 3422 39200 3478 40000
rect 3790 39200 3846 40000
rect 3974 39672 4030 39681
rect 3974 39607 4030 39616
rect 216 37262 244 39200
rect 204 37256 256 37262
rect 204 37198 256 37204
rect 584 36922 612 39200
rect 572 36916 624 36922
rect 572 36858 624 36864
rect 952 36378 980 39200
rect 1412 37346 1440 39200
rect 1412 37318 1532 37346
rect 1504 37262 1532 37318
rect 1492 37256 1544 37262
rect 1492 37198 1544 37204
rect 1780 36922 1808 39200
rect 1768 36916 1820 36922
rect 1768 36858 1820 36864
rect 1308 36848 1360 36854
rect 1308 36790 1360 36796
rect 940 36372 992 36378
rect 940 36314 992 36320
rect 938 27432 994 27441
rect 938 27367 994 27376
rect 756 25424 808 25430
rect 756 25366 808 25372
rect 480 22704 532 22710
rect 480 22646 532 22652
rect 388 21140 440 21146
rect 388 21082 440 21088
rect 18 17096 74 17105
rect 18 17031 74 17040
rect 32 1358 60 17031
rect 400 14074 428 21082
rect 492 16998 520 22646
rect 570 21176 626 21185
rect 570 21111 626 21120
rect 480 16992 532 16998
rect 480 16934 532 16940
rect 388 14068 440 14074
rect 388 14010 440 14016
rect 584 10606 612 21111
rect 662 20632 718 20641
rect 662 20567 718 20576
rect 572 10600 624 10606
rect 572 10542 624 10548
rect 676 5273 704 20567
rect 768 17134 796 25366
rect 846 23488 902 23497
rect 846 23423 902 23432
rect 756 17128 808 17134
rect 756 17070 808 17076
rect 756 16992 808 16998
rect 756 16934 808 16940
rect 768 15638 796 16934
rect 860 16182 888 23423
rect 848 16176 900 16182
rect 848 16118 900 16124
rect 756 15632 808 15638
rect 756 15574 808 15580
rect 768 14890 796 15574
rect 756 14884 808 14890
rect 756 14826 808 14832
rect 768 11778 796 14826
rect 952 14618 980 27367
rect 1216 25356 1268 25362
rect 1216 25298 1268 25304
rect 1032 23792 1084 23798
rect 1032 23734 1084 23740
rect 1044 18834 1072 23734
rect 1124 23044 1176 23050
rect 1124 22986 1176 22992
rect 1032 18828 1084 18834
rect 1032 18770 1084 18776
rect 1136 18766 1164 22986
rect 1228 20602 1256 25298
rect 1320 20806 1348 36790
rect 2148 36378 2176 39200
rect 2228 37256 2280 37262
rect 2228 37198 2280 37204
rect 2608 37210 2636 39200
rect 2870 39128 2926 39137
rect 2870 39063 2926 39072
rect 2780 37868 2832 37874
rect 2780 37810 2832 37816
rect 2792 37466 2820 37810
rect 2780 37460 2832 37466
rect 2780 37402 2832 37408
rect 2780 37256 2832 37262
rect 2608 37204 2780 37210
rect 2608 37198 2832 37204
rect 2136 36372 2188 36378
rect 2136 36314 2188 36320
rect 2044 35624 2096 35630
rect 1398 35592 1454 35601
rect 2044 35566 2096 35572
rect 1398 35527 1454 35536
rect 1412 35086 1440 35527
rect 1584 35488 1636 35494
rect 1584 35430 1636 35436
rect 1596 35290 1624 35430
rect 2056 35290 2084 35566
rect 2240 35290 2268 37198
rect 2412 37188 2464 37194
rect 2608 37182 2820 37198
rect 2412 37130 2464 37136
rect 2424 35834 2452 37130
rect 2596 37120 2648 37126
rect 2596 37062 2648 37068
rect 2504 36712 2556 36718
rect 2504 36654 2556 36660
rect 2412 35828 2464 35834
rect 2412 35770 2464 35776
rect 2412 35488 2464 35494
rect 2412 35430 2464 35436
rect 1584 35284 1636 35290
rect 1584 35226 1636 35232
rect 2044 35284 2096 35290
rect 2044 35226 2096 35232
rect 2228 35284 2280 35290
rect 2228 35226 2280 35232
rect 1400 35080 1452 35086
rect 1400 35022 1452 35028
rect 1412 34762 1440 35022
rect 1412 34734 1532 34762
rect 1400 34604 1452 34610
rect 1400 34546 1452 34552
rect 1412 34377 1440 34546
rect 1398 34368 1454 34377
rect 1398 34303 1454 34312
rect 1504 34202 1532 34734
rect 1584 34400 1636 34406
rect 1584 34342 1636 34348
rect 1492 34196 1544 34202
rect 1492 34138 1544 34144
rect 1492 33516 1544 33522
rect 1492 33458 1544 33464
rect 1400 33312 1452 33318
rect 1504 33289 1532 33458
rect 1400 33254 1452 33260
rect 1490 33280 1546 33289
rect 1412 31822 1440 33254
rect 1490 33215 1546 33224
rect 1492 32428 1544 32434
rect 1492 32370 1544 32376
rect 1504 32065 1532 32370
rect 1490 32056 1546 32065
rect 1490 31991 1546 32000
rect 1596 31890 1624 34342
rect 1676 32224 1728 32230
rect 1676 32166 1728 32172
rect 1584 31884 1636 31890
rect 1584 31826 1636 31832
rect 1688 31822 1716 32166
rect 1768 32020 1820 32026
rect 1768 31962 1820 31968
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1780 31482 1808 31962
rect 1860 31680 1912 31686
rect 1860 31622 1912 31628
rect 1768 31476 1820 31482
rect 1768 31418 1820 31424
rect 1400 31340 1452 31346
rect 1400 31282 1452 31288
rect 1412 30841 1440 31282
rect 1398 30832 1454 30841
rect 1398 30767 1454 30776
rect 1400 30252 1452 30258
rect 1400 30194 1452 30200
rect 1412 29753 1440 30194
rect 1584 30048 1636 30054
rect 1584 29990 1636 29996
rect 1398 29744 1454 29753
rect 1398 29679 1454 29688
rect 1492 28552 1544 28558
rect 1490 28520 1492 28529
rect 1544 28520 1546 28529
rect 1490 28455 1546 28464
rect 1400 28416 1452 28422
rect 1400 28358 1452 28364
rect 1412 28150 1440 28358
rect 1400 28144 1452 28150
rect 1400 28086 1452 28092
rect 1596 28014 1624 29990
rect 1676 28076 1728 28082
rect 1676 28018 1728 28024
rect 1584 28008 1636 28014
rect 1584 27950 1636 27956
rect 1584 27872 1636 27878
rect 1584 27814 1636 27820
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1412 27305 1440 27406
rect 1398 27296 1454 27305
rect 1398 27231 1454 27240
rect 1412 27130 1440 27231
rect 1400 27124 1452 27130
rect 1400 27066 1452 27072
rect 1596 26586 1624 27814
rect 1688 27674 1716 28018
rect 1676 27668 1728 27674
rect 1676 27610 1728 27616
rect 1872 27606 1900 31622
rect 1860 27600 1912 27606
rect 1860 27542 1912 27548
rect 2424 27470 2452 35430
rect 2516 33862 2544 36654
rect 2504 33856 2556 33862
rect 2504 33798 2556 33804
rect 2516 31754 2544 33798
rect 2608 32502 2636 37062
rect 2700 35766 2728 37182
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2688 35760 2740 35766
rect 2688 35702 2740 35708
rect 2792 35698 2820 36751
rect 2780 35692 2832 35698
rect 2780 35634 2832 35640
rect 2792 34746 2820 35634
rect 2884 35086 2912 39063
rect 2976 36922 3004 39200
rect 3146 37904 3202 37913
rect 3146 37839 3202 37848
rect 3056 37800 3108 37806
rect 3056 37742 3108 37748
rect 3068 37466 3096 37742
rect 3056 37460 3108 37466
rect 3056 37402 3108 37408
rect 2964 36916 3016 36922
rect 2964 36858 3016 36864
rect 3160 36174 3188 37839
rect 3436 36378 3464 39200
rect 3514 38584 3570 38593
rect 3514 38519 3570 38528
rect 3528 37466 3556 38519
rect 3516 37460 3568 37466
rect 3516 37402 3568 37408
rect 3698 37360 3754 37369
rect 3698 37295 3700 37304
rect 3752 37295 3754 37304
rect 3700 37266 3752 37272
rect 3804 37262 3832 39200
rect 3988 37738 4016 39607
rect 4158 39200 4214 40000
rect 4618 39200 4674 40000
rect 4986 39200 5042 40000
rect 5446 39200 5502 40000
rect 5814 39200 5870 40000
rect 6182 39200 6238 40000
rect 6642 39200 6698 40000
rect 7010 39200 7066 40000
rect 7378 39200 7434 40000
rect 7838 39200 7894 40000
rect 8206 39200 8262 40000
rect 8666 39200 8722 40000
rect 9034 39200 9090 40000
rect 9402 39200 9458 40000
rect 9862 39200 9918 40000
rect 10230 39200 10286 40000
rect 10690 39200 10746 40000
rect 11058 39200 11114 40000
rect 11426 39200 11482 40000
rect 11886 39200 11942 40000
rect 12254 39200 12310 40000
rect 12622 39200 12678 40000
rect 13082 39200 13138 40000
rect 13450 39200 13506 40000
rect 13910 39200 13966 40000
rect 14278 39200 14334 40000
rect 14646 39200 14702 40000
rect 14752 39222 15056 39250
rect 3976 37732 4028 37738
rect 4172 37720 4200 39200
rect 3976 37674 4028 37680
rect 4080 37692 4200 37720
rect 4080 37380 4108 37692
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4080 37352 4200 37380
rect 3792 37256 3844 37262
rect 3792 37198 3844 37204
rect 4172 36922 4200 37352
rect 4160 36916 4212 36922
rect 4160 36858 4212 36864
rect 3884 36780 3936 36786
rect 3884 36722 3936 36728
rect 3424 36372 3476 36378
rect 3424 36314 3476 36320
rect 3148 36168 3200 36174
rect 3148 36110 3200 36116
rect 2964 36032 3016 36038
rect 2964 35974 3016 35980
rect 2976 35630 3004 35974
rect 3160 35834 3188 36110
rect 3240 36100 3292 36106
rect 3240 36042 3292 36048
rect 3148 35828 3200 35834
rect 3148 35770 3200 35776
rect 2964 35624 3016 35630
rect 2964 35566 3016 35572
rect 2872 35080 2924 35086
rect 2872 35022 2924 35028
rect 2780 34740 2832 34746
rect 2780 34682 2832 34688
rect 2884 34202 2912 35022
rect 3252 34610 3280 36042
rect 3514 35048 3570 35057
rect 3514 34983 3570 34992
rect 3240 34604 3292 34610
rect 3240 34546 3292 34552
rect 3528 34542 3556 34983
rect 3896 34950 3924 36722
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4632 36378 4660 39200
rect 4710 37496 4766 37505
rect 4710 37431 4766 37440
rect 4724 37398 4752 37431
rect 4712 37392 4764 37398
rect 4712 37334 4764 37340
rect 5000 37262 5028 39200
rect 5354 37632 5410 37641
rect 5354 37567 5410 37576
rect 5172 37460 5224 37466
rect 5172 37402 5224 37408
rect 5080 37324 5132 37330
rect 5080 37266 5132 37272
rect 4804 37256 4856 37262
rect 4988 37256 5040 37262
rect 4804 37198 4856 37204
rect 4908 37204 4988 37210
rect 4908 37198 5040 37204
rect 4816 36922 4844 37198
rect 4908 37182 5028 37198
rect 4804 36916 4856 36922
rect 4804 36858 4856 36864
rect 4712 36780 4764 36786
rect 4712 36722 4764 36728
rect 4620 36372 4672 36378
rect 4620 36314 4672 36320
rect 4620 36236 4672 36242
rect 4620 36178 4672 36184
rect 4066 36136 4122 36145
rect 4066 36071 4122 36080
rect 4080 36038 4108 36071
rect 4068 36032 4120 36038
rect 4068 35974 4120 35980
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4632 35018 4660 36178
rect 4620 35012 4672 35018
rect 4620 34954 4672 34960
rect 3884 34944 3936 34950
rect 3884 34886 3936 34892
rect 3516 34536 3568 34542
rect 3516 34478 3568 34484
rect 2872 34196 2924 34202
rect 2872 34138 2924 34144
rect 3606 33824 3662 33833
rect 3606 33759 3662 33768
rect 3422 32600 3478 32609
rect 3422 32535 3478 32544
rect 2596 32496 2648 32502
rect 2596 32438 2648 32444
rect 3436 31754 3464 32535
rect 2516 31726 2636 31754
rect 2412 27464 2464 27470
rect 2412 27406 2464 27412
rect 1860 26784 1912 26790
rect 1860 26726 1912 26732
rect 2228 26784 2280 26790
rect 2228 26726 2280 26732
rect 1584 26580 1636 26586
rect 1584 26522 1636 26528
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 26217 1440 26318
rect 1398 26208 1454 26217
rect 1398 26143 1454 26152
rect 1400 25832 1452 25838
rect 1400 25774 1452 25780
rect 1412 25294 1440 25774
rect 1492 25696 1544 25702
rect 1492 25638 1544 25644
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1412 24993 1440 25230
rect 1398 24984 1454 24993
rect 1398 24919 1454 24928
rect 1400 24132 1452 24138
rect 1400 24074 1452 24080
rect 1412 23866 1440 24074
rect 1400 23860 1452 23866
rect 1400 23802 1452 23808
rect 1504 23769 1532 25638
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1596 24274 1624 25094
rect 1768 24404 1820 24410
rect 1768 24346 1820 24352
rect 1584 24268 1636 24274
rect 1584 24210 1636 24216
rect 1676 24200 1728 24206
rect 1676 24142 1728 24148
rect 1490 23760 1546 23769
rect 1490 23695 1492 23704
rect 1544 23695 1546 23704
rect 1492 23666 1544 23672
rect 1504 23635 1532 23666
rect 1688 23322 1716 24142
rect 1676 23316 1728 23322
rect 1676 23258 1728 23264
rect 1584 23180 1636 23186
rect 1584 23122 1636 23128
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 22681 1440 23054
rect 1490 22808 1546 22817
rect 1490 22743 1546 22752
rect 1398 22672 1454 22681
rect 1398 22607 1454 22616
rect 1400 22432 1452 22438
rect 1400 22374 1452 22380
rect 1308 20800 1360 20806
rect 1308 20742 1360 20748
rect 1216 20596 1268 20602
rect 1216 20538 1268 20544
rect 1124 18760 1176 18766
rect 1124 18702 1176 18708
rect 1412 17678 1440 22374
rect 1504 21554 1532 22743
rect 1596 22642 1624 23122
rect 1780 22778 1808 24346
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 1584 22636 1636 22642
rect 1584 22578 1636 22584
rect 1596 22094 1624 22578
rect 1596 22066 1808 22094
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1492 21548 1544 21554
rect 1492 21490 1544 21496
rect 1492 21412 1544 21418
rect 1492 21354 1544 21360
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1306 16144 1362 16153
rect 1306 16079 1308 16088
rect 1360 16079 1362 16088
rect 1308 16050 1360 16056
rect 1412 15570 1440 16594
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1306 14920 1362 14929
rect 1306 14855 1362 14864
rect 940 14612 992 14618
rect 940 14554 992 14560
rect 1030 14104 1086 14113
rect 1030 14039 1086 14048
rect 848 13456 900 13462
rect 848 13398 900 13404
rect 860 12434 888 13398
rect 860 12406 980 12434
rect 846 11792 902 11801
rect 768 11750 846 11778
rect 846 11727 902 11736
rect 860 5302 888 11727
rect 848 5296 900 5302
rect 662 5264 718 5273
rect 848 5238 900 5244
rect 662 5199 718 5208
rect 112 3936 164 3942
rect 112 3878 164 3884
rect 20 1352 72 1358
rect 20 1294 72 1300
rect 124 800 152 3878
rect 664 3664 716 3670
rect 664 3606 716 3612
rect 388 2984 440 2990
rect 388 2926 440 2932
rect 400 800 428 2926
rect 676 800 704 3606
rect 952 2553 980 12406
rect 1044 9450 1072 14039
rect 1216 13320 1268 13326
rect 1216 13262 1268 13268
rect 1124 12708 1176 12714
rect 1124 12650 1176 12656
rect 1032 9444 1084 9450
rect 1032 9386 1084 9392
rect 1136 6361 1164 12650
rect 1228 8022 1256 13262
rect 1320 11830 1348 14855
rect 1504 13394 1532 21354
rect 1596 17882 1624 21830
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 1688 17678 1716 21830
rect 1780 19145 1808 22066
rect 1872 21962 1900 26726
rect 2136 26376 2188 26382
rect 2136 26318 2188 26324
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 1964 22250 1992 25230
rect 2044 24676 2096 24682
rect 2044 24618 2096 24624
rect 2056 23497 2084 24618
rect 2042 23488 2098 23497
rect 2042 23423 2098 23432
rect 2148 23186 2176 26318
rect 2136 23180 2188 23186
rect 2136 23122 2188 23128
rect 2136 22976 2188 22982
rect 2136 22918 2188 22924
rect 2044 22636 2096 22642
rect 2044 22578 2096 22584
rect 2056 22386 2084 22578
rect 2148 22574 2176 22918
rect 2136 22568 2188 22574
rect 2136 22510 2188 22516
rect 2056 22358 2176 22386
rect 1964 22222 2084 22250
rect 1952 22160 2004 22166
rect 1952 22102 2004 22108
rect 1860 21956 1912 21962
rect 1860 21898 1912 21904
rect 1964 21729 1992 22102
rect 1950 21720 2006 21729
rect 1950 21655 2006 21664
rect 2056 21146 2084 22222
rect 2044 21140 2096 21146
rect 2044 21082 2096 21088
rect 2148 21026 2176 22358
rect 2240 22030 2268 26726
rect 2412 26580 2464 26586
rect 2412 26522 2464 26528
rect 2320 25696 2372 25702
rect 2320 25638 2372 25644
rect 2332 23882 2360 25638
rect 2424 24614 2452 26522
rect 2504 26240 2556 26246
rect 2504 26182 2556 26188
rect 2412 24608 2464 24614
rect 2410 24576 2412 24585
rect 2464 24576 2466 24585
rect 2410 24511 2466 24520
rect 2412 24064 2464 24070
rect 2410 24032 2412 24041
rect 2464 24032 2466 24041
rect 2410 23967 2466 23976
rect 2332 23854 2452 23882
rect 2320 22568 2372 22574
rect 2320 22510 2372 22516
rect 2228 22024 2280 22030
rect 2228 21966 2280 21972
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 1964 20998 2176 21026
rect 1964 20942 1992 20998
rect 1952 20936 2004 20942
rect 1872 20896 1952 20924
rect 1872 19378 1900 20896
rect 1952 20878 2004 20884
rect 2136 20936 2188 20942
rect 2136 20878 2188 20884
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 1952 19984 2004 19990
rect 1952 19926 2004 19932
rect 1964 19514 1992 19926
rect 2056 19922 2084 20334
rect 2148 20058 2176 20878
rect 2136 20052 2188 20058
rect 2136 19994 2188 20000
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2044 19780 2096 19786
rect 2044 19722 2096 19728
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 2056 19394 2084 19722
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1964 19366 2084 19394
rect 2136 19372 2188 19378
rect 1964 19174 1992 19366
rect 2136 19314 2188 19320
rect 2042 19272 2098 19281
rect 2042 19207 2098 19216
rect 1952 19168 2004 19174
rect 1766 19136 1822 19145
rect 1952 19110 2004 19116
rect 1766 19071 1822 19080
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1674 17232 1730 17241
rect 1674 17167 1676 17176
rect 1728 17167 1730 17176
rect 1676 17138 1728 17144
rect 1780 16794 1808 17818
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1596 16130 1624 16526
rect 1674 16280 1730 16289
rect 1674 16215 1676 16224
rect 1728 16215 1730 16224
rect 1676 16186 1728 16192
rect 1596 16102 1716 16130
rect 1584 16040 1636 16046
rect 1582 16008 1584 16017
rect 1636 16008 1638 16017
rect 1582 15943 1638 15952
rect 1688 15484 1716 16102
rect 1780 15706 1808 16730
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1768 15496 1820 15502
rect 1688 15456 1768 15484
rect 1768 15438 1820 15444
rect 1674 14512 1730 14521
rect 1674 14447 1730 14456
rect 1688 14414 1716 14447
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1584 13796 1636 13802
rect 1584 13738 1636 13744
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 1400 13252 1452 13258
rect 1400 13194 1452 13200
rect 1492 13252 1544 13258
rect 1492 13194 1544 13200
rect 1308 11824 1360 11830
rect 1308 11766 1360 11772
rect 1216 8016 1268 8022
rect 1216 7958 1268 7964
rect 1122 6352 1178 6361
rect 1122 6287 1178 6296
rect 1320 4826 1348 11766
rect 1412 9178 1440 13194
rect 1504 12850 1532 13194
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 1504 11354 1532 12786
rect 1596 12646 1624 13738
rect 1780 13705 1808 15438
rect 1872 14498 1900 17478
rect 1964 16574 1992 19110
rect 2056 18970 2084 19207
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2042 18864 2098 18873
rect 2042 18799 2098 18808
rect 2056 18766 2084 18799
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 2148 17626 2176 19314
rect 2240 17746 2268 21830
rect 2332 20466 2360 22510
rect 2320 20460 2372 20466
rect 2320 20402 2372 20408
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2332 19446 2360 20266
rect 2320 19440 2372 19446
rect 2320 19382 2372 19388
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2148 17598 2268 17626
rect 2134 17096 2190 17105
rect 2134 17031 2136 17040
rect 2188 17031 2190 17040
rect 2136 17002 2188 17008
rect 1964 16546 2084 16574
rect 1872 14470 1992 14498
rect 1766 13696 1822 13705
rect 1766 13631 1822 13640
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1688 12753 1716 12786
rect 1674 12744 1730 12753
rect 1674 12679 1730 12688
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 11558 1624 12582
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1582 10704 1638 10713
rect 1582 10639 1584 10648
rect 1636 10639 1638 10648
rect 1584 10610 1636 10616
rect 1582 10568 1638 10577
rect 1582 10503 1584 10512
rect 1636 10503 1638 10512
rect 1584 10474 1636 10480
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1504 8974 1532 9551
rect 1492 8968 1544 8974
rect 1398 8936 1454 8945
rect 1492 8910 1544 8916
rect 1398 8871 1454 8880
rect 1412 8498 1440 8871
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1596 7546 1624 10202
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1688 9178 1716 9998
rect 1780 9738 1808 13466
rect 1860 12368 1912 12374
rect 1858 12336 1860 12345
rect 1912 12336 1914 12345
rect 1858 12271 1914 12280
rect 1964 12238 1992 14470
rect 2056 13462 2084 16546
rect 2134 16416 2190 16425
rect 2134 16351 2190 16360
rect 2148 16250 2176 16351
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2148 15473 2176 15642
rect 2134 15464 2190 15473
rect 2134 15399 2190 15408
rect 2148 15366 2176 15399
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 1872 10305 1900 11834
rect 1858 10296 1914 10305
rect 1858 10231 1914 10240
rect 1780 9710 1900 9738
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1780 9042 1808 9522
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1780 8537 1808 8842
rect 1872 8634 1900 9710
rect 1964 9654 1992 12038
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1964 8809 1992 9318
rect 1950 8800 2006 8809
rect 1950 8735 2006 8744
rect 2056 8634 2084 13262
rect 2148 12986 2176 14962
rect 2240 13734 2268 17598
rect 2332 17202 2360 19382
rect 2424 19378 2452 23854
rect 2516 21554 2544 26182
rect 2608 22166 2636 31726
rect 3252 31726 3464 31754
rect 2870 31512 2926 31521
rect 2870 31447 2926 31456
rect 2780 27872 2832 27878
rect 2780 27814 2832 27820
rect 2688 27600 2740 27606
rect 2688 27542 2740 27548
rect 2700 24410 2728 27542
rect 2792 27538 2820 27814
rect 2780 27532 2832 27538
rect 2780 27474 2832 27480
rect 2884 25702 2912 31447
rect 3056 27328 3108 27334
rect 3056 27270 3108 27276
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 2964 25696 3016 25702
rect 2964 25638 3016 25644
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 2688 24404 2740 24410
rect 2688 24346 2740 24352
rect 2792 23474 2820 24686
rect 2976 24596 3004 25638
rect 3068 24750 3096 27270
rect 3252 25702 3280 31726
rect 3514 30288 3570 30297
rect 3514 30223 3570 30232
rect 3528 29034 3556 30223
rect 3516 29028 3568 29034
rect 3516 28970 3568 28976
rect 3422 27976 3478 27985
rect 3422 27911 3478 27920
rect 3240 25696 3292 25702
rect 3240 25638 3292 25644
rect 3148 25424 3200 25430
rect 3148 25366 3200 25372
rect 3160 25158 3188 25366
rect 3148 25152 3200 25158
rect 3148 25094 3200 25100
rect 3160 24954 3188 25094
rect 3148 24948 3200 24954
rect 3148 24890 3200 24896
rect 3436 24818 3464 27911
rect 3516 25696 3568 25702
rect 3516 25638 3568 25644
rect 3148 24812 3200 24818
rect 3148 24754 3200 24760
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3056 24744 3108 24750
rect 3056 24686 3108 24692
rect 2976 24568 3096 24596
rect 2872 24064 2924 24070
rect 2872 24006 2924 24012
rect 2884 23905 2912 24006
rect 2870 23896 2926 23905
rect 2870 23831 2872 23840
rect 2924 23831 2926 23840
rect 2872 23802 2924 23808
rect 2884 23771 2912 23802
rect 2964 23588 3016 23594
rect 2964 23530 3016 23536
rect 2700 23446 2820 23474
rect 2872 23520 2924 23526
rect 2976 23497 3004 23530
rect 2872 23462 2924 23468
rect 2962 23488 3018 23497
rect 2700 22642 2728 23446
rect 2884 22778 2912 23462
rect 2962 23423 3018 23432
rect 2872 22772 2924 22778
rect 2792 22732 2872 22760
rect 2688 22636 2740 22642
rect 2688 22578 2740 22584
rect 2596 22160 2648 22166
rect 2792 22114 2820 22732
rect 2872 22714 2924 22720
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2596 22102 2648 22108
rect 2700 22086 2820 22114
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2516 20584 2544 21490
rect 2608 21049 2636 21626
rect 2594 21040 2650 21049
rect 2594 20975 2650 20984
rect 2516 20556 2636 20584
rect 2608 20466 2636 20556
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2516 20074 2544 20402
rect 2700 20262 2728 22086
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2792 20369 2820 21966
rect 2884 21457 2912 22578
rect 3068 22137 3096 24568
rect 3054 22128 3110 22137
rect 2964 22092 3016 22098
rect 3160 22098 3188 24754
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3240 23588 3292 23594
rect 3240 23530 3292 23536
rect 3252 23322 3280 23530
rect 3240 23316 3292 23322
rect 3240 23258 3292 23264
rect 3436 22930 3464 23666
rect 3344 22902 3464 22930
rect 3240 22160 3292 22166
rect 3240 22102 3292 22108
rect 3054 22063 3110 22072
rect 3148 22092 3200 22098
rect 2964 22034 3016 22040
rect 3148 22034 3200 22040
rect 2870 21448 2926 21457
rect 2870 21383 2926 21392
rect 2870 20904 2926 20913
rect 2870 20839 2926 20848
rect 2778 20360 2834 20369
rect 2778 20295 2834 20304
rect 2688 20256 2740 20262
rect 2884 20244 2912 20839
rect 2688 20198 2740 20204
rect 2792 20216 2912 20244
rect 2516 20046 2728 20074
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2516 19514 2544 19926
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2700 19394 2728 20046
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2516 19366 2728 19394
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2318 13968 2374 13977
rect 2318 13903 2320 13912
rect 2372 13903 2374 13912
rect 2320 13874 2372 13880
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2320 13456 2372 13462
rect 2320 13398 2372 13404
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2240 12918 2268 13398
rect 2332 13258 2360 13398
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2228 12912 2280 12918
rect 2228 12854 2280 12860
rect 2424 12434 2452 14894
rect 2516 13462 2544 19366
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2700 18834 2728 19246
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2700 18193 2728 18566
rect 2686 18184 2742 18193
rect 2686 18119 2742 18128
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2608 17354 2636 18022
rect 2608 17326 2728 17354
rect 2792 17338 2820 20216
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 2884 18154 2912 19858
rect 2872 18148 2924 18154
rect 2872 18090 2924 18096
rect 2976 17921 3004 22034
rect 3148 21956 3200 21962
rect 3148 21898 3200 21904
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 3068 21146 3096 21490
rect 3056 21140 3108 21146
rect 3056 21082 3108 21088
rect 3056 20868 3108 20874
rect 3160 20856 3188 21898
rect 3108 20828 3188 20856
rect 3056 20810 3108 20816
rect 3148 20324 3200 20330
rect 3148 20266 3200 20272
rect 3056 20256 3108 20262
rect 3056 20198 3108 20204
rect 2962 17912 3018 17921
rect 2962 17847 3018 17856
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2608 16114 2636 17138
rect 2700 16561 2728 17326
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2884 16794 2912 17614
rect 3068 17610 3096 20198
rect 3160 18970 3188 20266
rect 3252 20058 3280 22102
rect 3344 21146 3372 22902
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3436 20448 3464 22170
rect 3528 22030 3556 25638
rect 3620 25430 3648 33759
rect 3896 29073 3924 34886
rect 4724 34649 4752 36722
rect 4908 35834 4936 37182
rect 4988 36168 5040 36174
rect 4988 36110 5040 36116
rect 5000 36009 5028 36110
rect 4986 36000 5042 36009
rect 4986 35935 5042 35944
rect 5092 35850 5120 37266
rect 4896 35828 4948 35834
rect 4896 35770 4948 35776
rect 5000 35822 5120 35850
rect 4710 34640 4766 34649
rect 4710 34575 4766 34584
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 3882 29064 3938 29073
rect 3882 28999 3938 29008
rect 4896 29028 4948 29034
rect 4896 28970 4948 28976
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4068 26988 4120 26994
rect 4068 26930 4120 26936
rect 4080 26761 4108 26930
rect 4066 26752 4122 26761
rect 4066 26687 4122 26696
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 3792 26308 3844 26314
rect 3792 26250 3844 26256
rect 3608 25424 3660 25430
rect 3608 25366 3660 25372
rect 3700 24064 3752 24070
rect 3700 24006 3752 24012
rect 3608 23588 3660 23594
rect 3608 23530 3660 23536
rect 3516 22024 3568 22030
rect 3516 21966 3568 21972
rect 3516 21888 3568 21894
rect 3620 21865 3648 23530
rect 3712 22710 3740 24006
rect 3804 23118 3832 26250
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 3884 25152 3936 25158
rect 3884 25094 3936 25100
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3700 22704 3752 22710
rect 3700 22646 3752 22652
rect 3804 22098 3832 22918
rect 3896 22642 3924 25094
rect 4158 24712 4214 24721
rect 4158 24647 4160 24656
rect 4212 24647 4214 24656
rect 4160 24618 4212 24624
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4066 24440 4122 24449
rect 4214 24432 4522 24452
rect 4066 24375 4122 24384
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3988 22953 4016 24006
rect 4080 23866 4108 24375
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4724 23497 4752 24550
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 4066 23488 4122 23497
rect 4710 23488 4766 23497
rect 4066 23423 4122 23432
rect 4080 23050 4108 23423
rect 4214 23420 4522 23440
rect 4710 23423 4766 23432
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4528 23248 4580 23254
rect 4528 23190 4580 23196
rect 4068 23044 4120 23050
rect 4068 22986 4120 22992
rect 4540 22964 4568 23190
rect 3974 22944 4030 22953
rect 4540 22936 4660 22964
rect 3974 22879 4030 22888
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 4068 22432 4120 22438
rect 4068 22374 4120 22380
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 3792 22092 3844 22098
rect 3792 22034 3844 22040
rect 3516 21830 3568 21836
rect 3606 21856 3662 21865
rect 3344 20420 3464 20448
rect 3240 20052 3292 20058
rect 3240 19994 3292 20000
rect 3344 19854 3372 20420
rect 3424 20324 3476 20330
rect 3424 20266 3476 20272
rect 3332 19848 3384 19854
rect 3238 19816 3294 19825
rect 3332 19790 3384 19796
rect 3238 19751 3294 19760
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3252 18766 3280 19751
rect 3332 19712 3384 19718
rect 3330 19680 3332 19689
rect 3384 19680 3386 19689
rect 3330 19615 3386 19624
rect 3436 19378 3464 20266
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3422 19272 3478 19281
rect 3422 19207 3478 19216
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 3146 18456 3202 18465
rect 3146 18391 3202 18400
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2686 16552 2742 16561
rect 2686 16487 2742 16496
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2700 14074 2728 16487
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2778 13968 2834 13977
rect 2778 13903 2834 13912
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2148 12406 2452 12434
rect 2148 10810 2176 12406
rect 2516 12306 2544 13126
rect 2608 13002 2636 13806
rect 2792 13394 2820 13903
rect 2870 13832 2926 13841
rect 2870 13767 2926 13776
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2884 13326 2912 13767
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2608 12974 2728 13002
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2608 12646 2636 12786
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2228 11620 2280 11626
rect 2228 11562 2280 11568
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 10169 2176 10610
rect 2134 10160 2190 10169
rect 2134 10095 2190 10104
rect 2240 9994 2268 11562
rect 2332 11150 2360 12038
rect 2410 11928 2466 11937
rect 2410 11863 2466 11872
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2424 10810 2452 11863
rect 2516 11694 2544 12106
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2148 9178 2176 9930
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2240 8786 2268 9658
rect 2148 8758 2268 8786
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1766 8528 1822 8537
rect 1766 8463 1822 8472
rect 2042 8392 2098 8401
rect 2042 8327 2098 8336
rect 2056 8090 2084 8327
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 7313 1440 7346
rect 1398 7304 1454 7313
rect 1398 7239 1454 7248
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 5914 1440 6258
rect 1504 6225 1532 6734
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 6322 1624 6598
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1490 6216 1546 6225
rect 1490 6151 1546 6160
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1308 4820 1360 4826
rect 1308 4762 1360 4768
rect 1412 4214 1440 5170
rect 1504 5001 1532 5646
rect 1490 4992 1546 5001
rect 1490 4927 1546 4936
rect 1596 4758 1624 6054
rect 1688 5370 1716 6258
rect 2148 6186 2176 8758
rect 2226 8664 2282 8673
rect 2332 8634 2360 10066
rect 2424 9722 2452 10610
rect 2516 10606 2544 11630
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2608 10282 2636 12378
rect 2700 12322 2728 12974
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2700 12294 2820 12322
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2516 10254 2636 10282
rect 2700 10266 2728 12174
rect 2792 12102 2820 12294
rect 2884 12238 2912 12854
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2976 11914 3004 12718
rect 3056 12096 3108 12102
rect 3160 12073 3188 18391
rect 3344 18086 3372 19110
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3332 17604 3384 17610
rect 3332 17546 3384 17552
rect 3238 17232 3294 17241
rect 3238 17167 3294 17176
rect 3252 16697 3280 17167
rect 3344 16998 3372 17546
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3238 16688 3294 16697
rect 3238 16623 3294 16632
rect 3344 16522 3372 16934
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3252 14414 3280 15438
rect 3344 15434 3372 16458
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 3240 14408 3292 14414
rect 3436 14385 3464 19207
rect 3528 16833 3556 21830
rect 3606 21791 3662 21800
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3514 16824 3570 16833
rect 3514 16759 3570 16768
rect 3620 15609 3648 20402
rect 3712 20233 3740 22034
rect 4080 21842 4108 22374
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 3988 21814 4108 21842
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 3698 20224 3754 20233
rect 3698 20159 3754 20168
rect 3698 20088 3754 20097
rect 3698 20023 3754 20032
rect 3712 19378 3740 20023
rect 3804 19922 3832 21490
rect 3884 21344 3936 21350
rect 3884 21286 3936 21292
rect 3896 21185 3924 21286
rect 3882 21176 3938 21185
rect 3882 21111 3938 21120
rect 3882 21040 3938 21049
rect 3882 20975 3938 20984
rect 3896 20806 3924 20975
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 3792 19916 3844 19922
rect 3792 19858 3844 19864
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3700 18896 3752 18902
rect 3700 18838 3752 18844
rect 3712 18601 3740 18838
rect 3804 18630 3832 19246
rect 3792 18624 3844 18630
rect 3698 18592 3754 18601
rect 3988 18612 4016 21814
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 3792 18566 3844 18572
rect 3896 18584 4016 18612
rect 3698 18527 3754 18536
rect 3698 18048 3754 18057
rect 3698 17983 3754 17992
rect 3712 17746 3740 17983
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3712 17338 3740 17478
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3804 16454 3832 18566
rect 3896 17270 3924 18584
rect 3974 18320 4030 18329
rect 3974 18255 3976 18264
rect 4028 18255 4030 18264
rect 3976 18226 4028 18232
rect 4080 17762 4108 21626
rect 4632 21434 4660 22936
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4724 22030 4752 22714
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4816 21593 4844 24006
rect 4908 23322 4936 28970
rect 5000 25498 5028 35822
rect 5184 35748 5212 37402
rect 5368 37398 5396 37567
rect 5356 37392 5408 37398
rect 5356 37334 5408 37340
rect 5460 36938 5488 39200
rect 5460 36922 5580 36938
rect 5460 36916 5592 36922
rect 5460 36910 5540 36916
rect 5540 36858 5592 36864
rect 5828 36378 5856 39200
rect 6196 37262 6224 39200
rect 6184 37256 6236 37262
rect 6184 37198 6236 37204
rect 6656 36922 6684 39200
rect 6644 36916 6696 36922
rect 6644 36858 6696 36864
rect 6460 36780 6512 36786
rect 6460 36722 6512 36728
rect 5816 36372 5868 36378
rect 5816 36314 5868 36320
rect 5540 36100 5592 36106
rect 5540 36042 5592 36048
rect 5092 35720 5212 35748
rect 5092 25498 5120 35720
rect 5552 34950 5580 36042
rect 6472 35562 6500 36722
rect 7024 36378 7052 39200
rect 7392 37262 7420 39200
rect 7656 37664 7708 37670
rect 7656 37606 7708 37612
rect 7668 37466 7696 37606
rect 7656 37460 7708 37466
rect 7656 37402 7708 37408
rect 7380 37256 7432 37262
rect 7380 37198 7432 37204
rect 7392 36378 7420 37198
rect 7852 36922 7880 39200
rect 8116 37392 8168 37398
rect 8114 37360 8116 37369
rect 8168 37360 8170 37369
rect 8114 37295 8170 37304
rect 7840 36916 7892 36922
rect 7840 36858 7892 36864
rect 8220 36394 8248 39200
rect 8680 37262 8708 39200
rect 8668 37256 8720 37262
rect 8668 37198 8720 37204
rect 9048 36922 9076 39200
rect 9416 36922 9444 39200
rect 9496 37936 9548 37942
rect 9496 37878 9548 37884
rect 9508 37466 9536 37878
rect 9496 37460 9548 37466
rect 9496 37402 9548 37408
rect 9876 37262 9904 39200
rect 9588 37256 9640 37262
rect 9588 37198 9640 37204
rect 9864 37256 9916 37262
rect 9864 37198 9916 37204
rect 9036 36916 9088 36922
rect 9036 36858 9088 36864
rect 9404 36916 9456 36922
rect 9404 36858 9456 36864
rect 8668 36780 8720 36786
rect 8668 36722 8720 36728
rect 9496 36780 9548 36786
rect 9496 36722 9548 36728
rect 8220 36378 8340 36394
rect 7012 36372 7064 36378
rect 7012 36314 7064 36320
rect 7380 36372 7432 36378
rect 8220 36372 8352 36378
rect 8220 36366 8300 36372
rect 7380 36314 7432 36320
rect 8300 36314 8352 36320
rect 6920 36168 6972 36174
rect 6920 36110 6972 36116
rect 7380 36168 7432 36174
rect 7380 36110 7432 36116
rect 6460 35556 6512 35562
rect 6460 35498 6512 35504
rect 6368 35012 6420 35018
rect 6368 34954 6420 34960
rect 5540 34944 5592 34950
rect 5540 34886 5592 34892
rect 5172 34604 5224 34610
rect 5172 34546 5224 34552
rect 4988 25492 5040 25498
rect 4988 25434 5040 25440
rect 5080 25492 5132 25498
rect 5080 25434 5132 25440
rect 5000 23905 5028 25434
rect 5080 24608 5132 24614
rect 5080 24550 5132 24556
rect 5092 24138 5120 24550
rect 5080 24132 5132 24138
rect 5080 24074 5132 24080
rect 4986 23896 5042 23905
rect 4986 23831 5042 23840
rect 4988 23792 5040 23798
rect 4988 23734 5040 23740
rect 5080 23792 5132 23798
rect 5080 23734 5132 23740
rect 5000 23322 5028 23734
rect 4896 23316 4948 23322
rect 4896 23258 4948 23264
rect 4988 23316 5040 23322
rect 4988 23258 5040 23264
rect 4894 23216 4950 23225
rect 4894 23151 4950 23160
rect 4802 21584 4858 21593
rect 4802 21519 4858 21528
rect 4632 21406 4844 21434
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4632 21146 4660 21286
rect 4620 21140 4672 21146
rect 4620 21082 4672 21088
rect 4436 21072 4488 21078
rect 4250 21040 4306 21049
rect 4724 21026 4752 21286
rect 4488 21020 4752 21026
rect 4436 21014 4752 21020
rect 4448 20998 4752 21014
rect 4816 21010 4844 21406
rect 4804 21004 4856 21010
rect 4250 20975 4306 20984
rect 4264 20466 4292 20975
rect 4804 20946 4856 20952
rect 4342 20904 4398 20913
rect 4342 20839 4344 20848
rect 4396 20839 4398 20848
rect 4344 20810 4396 20816
rect 4356 20602 4384 20810
rect 4712 20800 4764 20806
rect 4712 20742 4764 20748
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4528 20392 4580 20398
rect 4526 20360 4528 20369
rect 4580 20360 4582 20369
rect 4526 20295 4582 20304
rect 4618 20224 4674 20233
rect 4214 20156 4522 20176
rect 4618 20159 4674 20168
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4250 19952 4306 19961
rect 4250 19887 4306 19896
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 4172 19242 4200 19654
rect 4264 19242 4292 19887
rect 4526 19408 4582 19417
rect 4632 19394 4660 20159
rect 4724 20058 4752 20742
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4724 19417 4752 19790
rect 4582 19366 4660 19394
rect 4710 19408 4766 19417
rect 4526 19343 4582 19352
rect 4710 19343 4766 19352
rect 4344 19304 4396 19310
rect 4396 19264 4752 19292
rect 4344 19246 4396 19252
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4526 18864 4582 18873
rect 4526 18799 4582 18808
rect 4540 18766 4568 18799
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4158 18592 4214 18601
rect 4158 18527 4214 18536
rect 4172 18426 4200 18527
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4632 18306 4660 19110
rect 4724 18970 4752 19264
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4448 18290 4660 18306
rect 4436 18284 4660 18290
rect 4488 18278 4660 18284
rect 4436 18226 4488 18232
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4080 17734 4200 17762
rect 4632 17746 4660 18278
rect 4068 17672 4120 17678
rect 3988 17620 4068 17626
rect 3988 17614 4120 17620
rect 3988 17598 4108 17614
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3988 17134 4016 17598
rect 4066 17368 4122 17377
rect 4066 17303 4122 17312
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3988 16590 4016 17070
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 4080 16250 4108 17303
rect 4172 17270 4200 17734
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4632 17626 4660 17682
rect 4448 17598 4660 17626
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 4448 17202 4476 17598
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4528 16108 4580 16114
rect 4632 16096 4660 17598
rect 4724 16658 4752 18634
rect 4816 17542 4844 20198
rect 4908 19922 4936 23151
rect 4988 22976 5040 22982
rect 4988 22918 5040 22924
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 5000 18358 5028 22918
rect 5092 22778 5120 23734
rect 5184 23497 5212 34546
rect 6092 26512 6144 26518
rect 6092 26454 6144 26460
rect 5724 25696 5776 25702
rect 5724 25638 5776 25644
rect 5448 25492 5500 25498
rect 5448 25434 5500 25440
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5170 23488 5226 23497
rect 5170 23423 5226 23432
rect 5172 22976 5224 22982
rect 5172 22918 5224 22924
rect 5080 22772 5132 22778
rect 5080 22714 5132 22720
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5092 21962 5120 22510
rect 5184 22273 5212 22918
rect 5170 22264 5226 22273
rect 5170 22199 5226 22208
rect 5276 22098 5304 24754
rect 5356 23044 5408 23050
rect 5356 22986 5408 22992
rect 5368 22574 5396 22986
rect 5356 22568 5408 22574
rect 5356 22510 5408 22516
rect 5264 22092 5316 22098
rect 5264 22034 5316 22040
rect 5080 21956 5132 21962
rect 5080 21898 5132 21904
rect 5172 21956 5224 21962
rect 5172 21898 5224 21904
rect 5184 21486 5212 21898
rect 5354 21720 5410 21729
rect 5354 21655 5410 21664
rect 5368 21622 5396 21655
rect 5356 21616 5408 21622
rect 5356 21558 5408 21564
rect 5460 21554 5488 25434
rect 5736 25294 5764 25638
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5908 25288 5960 25294
rect 5908 25230 5960 25236
rect 5816 24608 5868 24614
rect 5816 24550 5868 24556
rect 5724 24200 5776 24206
rect 5724 24142 5776 24148
rect 5630 23624 5686 23633
rect 5630 23559 5632 23568
rect 5684 23559 5686 23568
rect 5632 23530 5684 23536
rect 5540 23248 5592 23254
rect 5538 23216 5540 23225
rect 5592 23216 5594 23225
rect 5538 23151 5594 23160
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5552 22234 5580 22578
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5632 22160 5684 22166
rect 5632 22102 5684 22108
rect 5540 21956 5592 21962
rect 5540 21898 5592 21904
rect 5448 21548 5500 21554
rect 5448 21490 5500 21496
rect 5172 21480 5224 21486
rect 5172 21422 5224 21428
rect 5264 21480 5316 21486
rect 5460 21457 5488 21490
rect 5264 21422 5316 21428
rect 5446 21448 5502 21457
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 4988 18352 5040 18358
rect 4988 18294 5040 18300
rect 5092 17610 5120 21082
rect 5184 20466 5212 21422
rect 5276 21350 5304 21422
rect 5446 21383 5502 21392
rect 5264 21344 5316 21350
rect 5552 21298 5580 21898
rect 5264 21286 5316 21292
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4986 17504 5042 17513
rect 4986 17439 5042 17448
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4580 16068 4660 16096
rect 4528 16050 4580 16056
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15706 3924 15846
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3606 15600 3662 15609
rect 3606 15535 3662 15544
rect 4618 15600 4674 15609
rect 4618 15535 4620 15544
rect 4672 15535 4674 15544
rect 4620 15506 4672 15512
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4710 15464 4766 15473
rect 4066 15056 4122 15065
rect 4540 15026 4568 15438
rect 4710 15399 4766 15408
rect 4066 14991 4122 15000
rect 4528 15020 4580 15026
rect 4080 14618 4108 14991
rect 4580 14980 4660 15008
rect 4528 14962 4580 14968
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3608 14408 3660 14414
rect 3240 14350 3292 14356
rect 3422 14376 3478 14385
rect 3252 14278 3280 14350
rect 3608 14350 3660 14356
rect 3422 14311 3478 14320
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3056 12038 3108 12044
rect 3146 12064 3202 12073
rect 2792 11886 3004 11914
rect 3068 11914 3096 12038
rect 3146 11999 3202 12008
rect 3068 11886 3188 11914
rect 2792 10470 2820 11886
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2884 11393 2912 11630
rect 2870 11384 2926 11393
rect 2976 11354 3004 11698
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2870 11319 2926 11328
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2688 10260 2740 10266
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2226 8599 2282 8608
rect 2320 8628 2372 8634
rect 2240 8498 2268 8599
rect 2320 8570 2372 8576
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2424 6390 2452 9522
rect 2516 6458 2544 10254
rect 2688 10202 2740 10208
rect 2596 10192 2648 10198
rect 2594 10160 2596 10169
rect 2648 10160 2650 10169
rect 2594 10095 2650 10104
rect 2884 9874 2912 11222
rect 2792 9846 2912 9874
rect 2594 8256 2650 8265
rect 2594 8191 2650 8200
rect 2608 8090 2636 8191
rect 2686 8120 2742 8129
rect 2596 8084 2648 8090
rect 2686 8055 2742 8064
rect 2596 8026 2648 8032
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2136 6180 2188 6186
rect 2136 6122 2188 6128
rect 2148 5370 2176 6122
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 1584 4752 1636 4758
rect 1584 4694 1636 4700
rect 2042 4720 2098 4729
rect 2042 4655 2098 4664
rect 2056 4622 2084 4655
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 1400 4208 1452 4214
rect 1400 4150 1452 4156
rect 1308 4004 1360 4010
rect 1308 3946 1360 3952
rect 1032 3528 1084 3534
rect 1032 3470 1084 3476
rect 938 2544 994 2553
rect 938 2479 994 2488
rect 940 1352 992 1358
rect 940 1294 992 1300
rect 110 0 166 800
rect 386 0 442 800
rect 662 0 718 800
rect 952 377 980 1294
rect 1044 800 1072 3470
rect 1320 800 1348 3946
rect 1412 3777 1440 4150
rect 1398 3768 1454 3777
rect 1398 3703 1454 3712
rect 1688 800 1716 4558
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1964 800 1992 3878
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2332 2394 2360 2926
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2240 2366 2360 2394
rect 2240 800 2268 2366
rect 2608 800 2636 2858
rect 2700 2582 2728 8055
rect 2792 6730 2820 9846
rect 2870 9752 2926 9761
rect 2870 9687 2926 9696
rect 2884 8974 2912 9687
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2884 6934 2912 7346
rect 2872 6928 2924 6934
rect 2872 6870 2924 6876
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2792 6322 2820 6666
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2884 5846 2912 6666
rect 2976 6458 3004 11290
rect 3068 6662 3096 11494
rect 3160 11150 3188 11886
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3146 10840 3202 10849
rect 3146 10775 3202 10784
rect 3160 8498 3188 10775
rect 3252 10674 3280 13670
rect 3332 13456 3384 13462
rect 3332 13398 3384 13404
rect 3344 12782 3372 13398
rect 3528 13161 3556 13874
rect 3620 13870 3648 14350
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3712 13308 3740 14282
rect 3804 13410 3832 14418
rect 3884 14272 3936 14278
rect 3882 14240 3884 14249
rect 3936 14240 3938 14249
rect 3882 14175 3938 14184
rect 3988 14090 4016 14554
rect 4344 14544 4396 14550
rect 4342 14512 4344 14521
rect 4396 14512 4398 14521
rect 4342 14447 4398 14456
rect 4632 14414 4660 14980
rect 4724 14482 4752 15399
rect 4816 14550 4844 17206
rect 5000 15638 5028 17439
rect 5184 16114 5212 19994
rect 5276 16182 5304 21286
rect 5460 21270 5580 21298
rect 5460 21026 5488 21270
rect 5368 21010 5488 21026
rect 5368 21004 5500 21010
rect 5368 20998 5448 21004
rect 5368 19854 5396 20998
rect 5448 20946 5500 20952
rect 5540 20936 5592 20942
rect 5446 20904 5502 20913
rect 5540 20878 5592 20884
rect 5446 20839 5502 20848
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5354 19680 5410 19689
rect 5354 19615 5410 19624
rect 5368 19417 5396 19615
rect 5354 19408 5410 19417
rect 5354 19343 5410 19352
rect 5368 18442 5396 19343
rect 5460 18873 5488 20839
rect 5552 20777 5580 20878
rect 5538 20768 5594 20777
rect 5538 20703 5594 20712
rect 5538 20632 5594 20641
rect 5538 20567 5594 20576
rect 5552 20466 5580 20567
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5552 19446 5580 19654
rect 5644 19514 5672 22102
rect 5736 22098 5764 24142
rect 5724 22092 5776 22098
rect 5724 22034 5776 22040
rect 5724 21072 5776 21078
rect 5724 21014 5776 21020
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5736 19446 5764 21014
rect 5828 20505 5856 24550
rect 5920 22778 5948 25230
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 6012 23118 6040 24006
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 5908 22772 5960 22778
rect 5908 22714 5960 22720
rect 6012 22438 6040 23054
rect 6104 22438 6132 26454
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6288 24138 6316 24550
rect 6276 24132 6328 24138
rect 6276 24074 6328 24080
rect 6184 23588 6236 23594
rect 6184 23530 6236 23536
rect 6196 22817 6224 23530
rect 6288 23322 6316 24074
rect 6276 23316 6328 23322
rect 6276 23258 6328 23264
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6182 22808 6238 22817
rect 6182 22743 6238 22752
rect 6288 22710 6316 22918
rect 6276 22704 6328 22710
rect 6276 22646 6328 22652
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6274 22536 6330 22545
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 6092 22432 6144 22438
rect 6092 22374 6144 22380
rect 6012 22234 6040 22374
rect 6000 22228 6052 22234
rect 6000 22170 6052 22176
rect 6196 22098 6224 22510
rect 6274 22471 6330 22480
rect 6184 22094 6236 22098
rect 5920 22092 6236 22094
rect 5920 22066 6184 22092
rect 5920 21690 5948 22066
rect 6184 22034 6236 22040
rect 6288 21978 6316 22471
rect 6012 21950 6316 21978
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5814 20496 5870 20505
rect 5814 20431 5816 20440
rect 5868 20431 5870 20440
rect 5816 20402 5868 20408
rect 5816 19780 5868 19786
rect 5816 19722 5868 19728
rect 5828 19514 5856 19722
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5540 19440 5592 19446
rect 5540 19382 5592 19388
rect 5724 19440 5776 19446
rect 5724 19382 5776 19388
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5446 18864 5502 18873
rect 5644 18834 5672 19246
rect 5446 18799 5502 18808
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5368 18414 5580 18442
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5354 18048 5410 18057
rect 5354 17983 5410 17992
rect 5264 16176 5316 16182
rect 5264 16118 5316 16124
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4620 14408 4672 14414
rect 4066 14376 4122 14385
rect 4620 14350 4672 14356
rect 4066 14311 4122 14320
rect 3896 14062 4016 14090
rect 3896 13530 3924 14062
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3882 13424 3938 13433
rect 3804 13382 3882 13410
rect 3882 13359 3884 13368
rect 3936 13359 3938 13368
rect 3884 13330 3936 13336
rect 3792 13320 3844 13326
rect 3712 13280 3792 13308
rect 3882 13288 3938 13297
rect 3844 13268 3882 13274
rect 3792 13262 3882 13268
rect 3804 13246 3882 13262
rect 3882 13223 3938 13232
rect 3792 13184 3844 13190
rect 3514 13152 3570 13161
rect 3792 13126 3844 13132
rect 3514 13087 3570 13096
rect 3514 13016 3570 13025
rect 3514 12951 3516 12960
rect 3568 12951 3570 12960
rect 3516 12922 3568 12928
rect 3608 12912 3660 12918
rect 3608 12854 3660 12860
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3514 12744 3570 12753
rect 3344 10810 3372 12718
rect 3514 12679 3570 12688
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3436 11762 3464 12174
rect 3528 11762 3556 12679
rect 3620 11898 3648 12854
rect 3700 12640 3752 12646
rect 3804 12617 3832 13126
rect 3884 12640 3936 12646
rect 3700 12582 3752 12588
rect 3790 12608 3846 12617
rect 3712 12306 3740 12582
rect 3884 12582 3936 12588
rect 3790 12543 3846 12552
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3516 11756 3568 11762
rect 3712 11744 3740 12242
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3516 11698 3568 11704
rect 3620 11716 3740 11744
rect 3436 11354 3464 11698
rect 3620 11370 3648 11716
rect 3804 11529 3832 12174
rect 3896 12170 3924 12582
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3988 11898 4016 13806
rect 4080 13326 4108 14311
rect 4528 13932 4580 13938
rect 4632 13920 4660 14350
rect 4580 13892 4660 13920
rect 4528 13874 4580 13880
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4172 13161 4200 13398
rect 4632 13326 4660 13892
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4158 13152 4214 13161
rect 4158 13087 4214 13096
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4528 12844 4580 12850
rect 4632 12832 4660 13262
rect 4580 12804 4660 12832
rect 4528 12786 4580 12792
rect 4080 12434 4108 12786
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4080 12406 4200 12434
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3790 11520 3846 11529
rect 3790 11455 3846 11464
rect 3896 11370 3924 11698
rect 3988 11665 4016 11698
rect 3974 11656 4030 11665
rect 4080 11626 4108 12038
rect 4172 11898 4200 12406
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4264 11762 4292 12242
rect 4540 12209 4568 12242
rect 4526 12200 4582 12209
rect 4526 12135 4582 12144
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 3974 11591 4030 11600
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3528 11342 3648 11370
rect 3712 11342 3924 11370
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3252 8974 3280 10610
rect 3436 9518 3464 11086
rect 3528 9602 3556 11342
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3620 10033 3648 10066
rect 3606 10024 3662 10033
rect 3606 9959 3662 9968
rect 3606 9752 3662 9761
rect 3606 9687 3608 9696
rect 3660 9687 3662 9696
rect 3608 9658 3660 9664
rect 3528 9574 3648 9602
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3514 9480 3570 9489
rect 3620 9450 3648 9574
rect 3514 9415 3516 9424
rect 3568 9415 3570 9424
rect 3608 9444 3660 9450
rect 3516 9386 3568 9392
rect 3608 9386 3660 9392
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2976 5846 3004 6394
rect 3068 5914 3096 6598
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2792 1018 2820 2382
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 2884 1834 2912 2314
rect 2872 1828 2924 1834
rect 2872 1770 2924 1776
rect 2884 1465 2912 1770
rect 2976 1601 3004 3470
rect 3068 2689 3096 4490
rect 3054 2680 3110 2689
rect 3054 2615 3110 2624
rect 3068 2145 3096 2615
rect 3054 2136 3110 2145
rect 3054 2071 3110 2080
rect 2962 1592 3018 1601
rect 2962 1527 3018 1536
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 2976 1306 3004 1527
rect 2884 1278 3004 1306
rect 2780 1012 2832 1018
rect 2780 954 2832 960
rect 2792 921 2820 954
rect 2778 912 2834 921
rect 2778 847 2834 856
rect 2884 800 2912 1278
rect 3160 921 3188 8434
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3252 8090 3280 8298
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3344 7002 3372 8842
rect 3422 8664 3478 8673
rect 3422 8599 3424 8608
rect 3476 8599 3478 8608
rect 3424 8570 3476 8576
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3620 7546 3648 7686
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3712 6730 3740 11342
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3804 10538 3832 10610
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3804 9654 3832 10474
rect 3896 10130 3924 11018
rect 3988 10470 4016 11494
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4172 10849 4200 10950
rect 4158 10840 4214 10849
rect 4158 10775 4214 10784
rect 4264 10674 4292 11154
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4540 10606 4568 11018
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10180 4016 10406
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4632 10198 4660 12804
rect 4712 12844 4764 12850
rect 4764 12804 4844 12832
rect 4712 12786 4764 12792
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 11762 4752 12582
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4710 11112 4766 11121
rect 4710 11047 4766 11056
rect 4620 10192 4672 10198
rect 3988 10152 4200 10180
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 4172 10062 4200 10152
rect 4620 10134 4672 10140
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9761 3924 9862
rect 3882 9752 3938 9761
rect 3882 9687 3938 9696
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3882 9616 3938 9625
rect 3882 9551 3938 9560
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3804 8090 3832 8910
rect 3896 8412 3924 9551
rect 3988 8566 4016 9930
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3896 8384 4016 8412
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3804 7546 3832 8026
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3804 6440 3832 7482
rect 3896 6914 3924 8230
rect 3988 8106 4016 8384
rect 4080 8294 4108 9998
rect 4540 9994 4568 10066
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4356 9586 4384 9658
rect 4540 9625 4568 9930
rect 4526 9616 4582 9625
rect 4344 9580 4396 9586
rect 4526 9551 4582 9560
rect 4620 9580 4672 9586
rect 4344 9522 4396 9528
rect 4620 9522 4672 9528
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4632 8974 4660 9522
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4724 8498 4752 11047
rect 4816 8634 4844 12804
rect 5000 12481 5028 13874
rect 5276 13841 5304 13874
rect 5262 13832 5318 13841
rect 5262 13767 5318 13776
rect 5368 13530 5396 17983
rect 5460 17678 5488 18294
rect 5552 17785 5580 18414
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5538 17776 5594 17785
rect 5538 17711 5594 17720
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5552 17524 5580 17614
rect 5460 17496 5580 17524
rect 5460 16522 5488 17496
rect 5644 17338 5672 18226
rect 5736 17338 5764 19382
rect 5828 17746 5856 19450
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5920 18902 5948 19110
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 6012 18057 6040 21950
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6184 20392 6236 20398
rect 6184 20334 6236 20340
rect 6196 19990 6224 20334
rect 6184 19984 6236 19990
rect 6184 19926 6236 19932
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6104 19417 6132 19790
rect 6090 19408 6146 19417
rect 6090 19343 6146 19352
rect 6092 19236 6144 19242
rect 6092 19178 6144 19184
rect 5998 18048 6054 18057
rect 5998 17983 6054 17992
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 6104 17626 6132 19178
rect 6196 17814 6224 19926
rect 6288 18290 6316 21830
rect 6380 21010 6408 34954
rect 6736 34944 6788 34950
rect 6736 34886 6788 34892
rect 6644 26852 6696 26858
rect 6644 26794 6696 26800
rect 6656 26586 6684 26794
rect 6644 26580 6696 26586
rect 6644 26522 6696 26528
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6460 24064 6512 24070
rect 6460 24006 6512 24012
rect 6472 23730 6500 24006
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6472 22642 6500 23666
rect 6656 23633 6684 25094
rect 6642 23624 6698 23633
rect 6642 23559 6698 23568
rect 6550 23488 6606 23497
rect 6550 23423 6606 23432
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6472 21010 6500 22374
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 6380 19990 6408 20538
rect 6368 19984 6420 19990
rect 6368 19926 6420 19932
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6276 18284 6328 18290
rect 6276 18226 6328 18232
rect 6380 18086 6408 19790
rect 6472 19378 6500 20810
rect 6564 20602 6592 23423
rect 6644 23316 6696 23322
rect 6644 23258 6696 23264
rect 6656 22574 6684 23258
rect 6644 22568 6696 22574
rect 6644 22510 6696 22516
rect 6642 21856 6698 21865
rect 6642 21791 6698 21800
rect 6656 21622 6684 21791
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 6656 20602 6684 20946
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6656 20369 6684 20402
rect 6642 20360 6698 20369
rect 6642 20295 6698 20304
rect 6550 20088 6606 20097
rect 6550 20023 6606 20032
rect 6644 20052 6696 20058
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6564 19258 6592 20023
rect 6644 19994 6696 20000
rect 6472 19230 6592 19258
rect 6656 19242 6684 19994
rect 6748 19922 6776 34886
rect 6828 34536 6880 34542
rect 6828 34478 6880 34484
rect 6840 26586 6868 34478
rect 6932 26897 6960 36110
rect 7392 27169 7420 36110
rect 8024 36032 8076 36038
rect 8024 35974 8076 35980
rect 7472 27668 7524 27674
rect 7472 27610 7524 27616
rect 7378 27160 7434 27169
rect 7378 27095 7434 27104
rect 6918 26888 6974 26897
rect 6918 26823 6974 26832
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6840 22094 6868 26522
rect 6918 26208 6974 26217
rect 6918 26143 6974 26152
rect 6932 26042 6960 26143
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7012 24064 7064 24070
rect 7012 24006 7064 24012
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 6932 22234 6960 23190
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 6840 22066 6960 22094
rect 6932 21894 6960 22066
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 6826 20768 6882 20777
rect 6826 20703 6882 20712
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 6644 19236 6696 19242
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 5828 17598 6132 17626
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5724 16992 5776 16998
rect 5538 16960 5594 16969
rect 5724 16934 5776 16940
rect 5538 16895 5594 16904
rect 5448 16516 5500 16522
rect 5448 16458 5500 16464
rect 5552 14521 5580 16895
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 5644 15366 5672 16458
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5538 14512 5594 14521
rect 5538 14447 5594 14456
rect 5439 14408 5491 14414
rect 5439 14350 5491 14356
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 4986 12472 5042 12481
rect 4986 12407 5042 12416
rect 5460 12374 5488 14350
rect 5552 13705 5580 14447
rect 5644 14006 5672 14894
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5538 13696 5594 13705
rect 5538 13631 5594 13640
rect 5736 12434 5764 16934
rect 5828 16810 5856 17598
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5920 16998 5948 17274
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5828 16782 5948 16810
rect 5920 14822 5948 16782
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5828 14249 5856 14758
rect 5814 14240 5870 14249
rect 5814 14175 5870 14184
rect 5920 12889 5948 14758
rect 5906 12880 5962 12889
rect 5906 12815 5962 12824
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12442 5948 12582
rect 5908 12436 5960 12442
rect 5736 12406 5856 12434
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5828 12322 5856 12406
rect 5908 12378 5960 12384
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4908 11393 4936 12038
rect 4986 11656 5042 11665
rect 4986 11591 4988 11600
rect 5040 11591 5042 11600
rect 4988 11562 5040 11568
rect 4894 11384 4950 11393
rect 4894 11319 4950 11328
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 3988 8078 4108 8106
rect 4080 6984 4108 8078
rect 4342 7848 4398 7857
rect 4342 7783 4398 7792
rect 4356 7750 4384 7783
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4618 7032 4674 7041
rect 4080 6956 4568 6984
rect 4618 6967 4674 6976
rect 4804 6996 4856 7002
rect 3896 6886 4108 6914
rect 3712 6412 3832 6440
rect 3882 6488 3938 6497
rect 4080 6458 4108 6886
rect 4434 6896 4490 6905
rect 4434 6831 4436 6840
rect 4488 6831 4490 6840
rect 4436 6802 4488 6808
rect 4540 6610 4568 6956
rect 4632 6769 4660 6967
rect 4804 6938 4856 6944
rect 4618 6760 4674 6769
rect 4618 6695 4674 6704
rect 4540 6582 4660 6610
rect 4068 6452 4120 6458
rect 3882 6423 3884 6432
rect 3330 6216 3386 6225
rect 3330 6151 3386 6160
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3146 912 3202 921
rect 3146 847 3202 856
rect 3252 800 3280 3878
rect 3344 1329 3372 6151
rect 3712 5914 3740 6412
rect 3936 6423 3938 6432
rect 3884 6394 3936 6400
rect 3988 6412 4068 6440
rect 3988 6338 4016 6412
rect 4068 6394 4120 6400
rect 3804 6310 4016 6338
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3422 3088 3478 3097
rect 3422 3023 3424 3032
rect 3476 3023 3478 3032
rect 3424 2994 3476 3000
rect 3330 1320 3386 1329
rect 3330 1255 3386 1264
rect 3804 814 3832 6310
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4632 5794 4660 6582
rect 4540 5766 4660 5794
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3974 5536 4030 5545
rect 3974 5471 4030 5480
rect 3988 5166 4016 5471
rect 4080 5409 4108 5646
rect 4066 5400 4122 5409
rect 4066 5335 4122 5344
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 4080 4457 4108 5238
rect 4540 5098 4568 5766
rect 4618 5536 4674 5545
rect 4618 5471 4674 5480
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4632 4826 4660 5471
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4724 4554 4752 4966
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4066 4448 4122 4457
rect 4816 4434 4844 6938
rect 4908 6254 4936 10406
rect 5000 8498 5028 10610
rect 5092 10198 5120 12106
rect 5276 11694 5304 12310
rect 5540 12300 5592 12306
rect 5828 12294 5948 12322
rect 5540 12242 5592 12248
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5184 10470 5212 11290
rect 5460 11150 5488 12106
rect 5552 11218 5580 12242
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5722 11928 5778 11937
rect 5722 11863 5724 11872
rect 5776 11863 5778 11872
rect 5724 11834 5776 11840
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5092 7886 5120 9862
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5184 7954 5212 9522
rect 5276 8430 5304 10678
rect 5368 10674 5396 10950
rect 5552 10742 5580 11018
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5368 9994 5396 10610
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5460 10130 5488 10542
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 10266 5580 10406
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5460 9518 5488 10066
rect 5538 9616 5594 9625
rect 5538 9551 5594 9560
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5356 9376 5408 9382
rect 5354 9344 5356 9353
rect 5408 9344 5410 9353
rect 5354 9279 5410 9288
rect 5460 9178 5488 9454
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5460 8294 5488 8910
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 5000 6984 5028 7754
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5092 7313 5120 7482
rect 5276 7342 5304 8230
rect 5552 8106 5580 9551
rect 5644 8974 5672 11494
rect 5828 11286 5856 12174
rect 5816 11280 5868 11286
rect 5816 11222 5868 11228
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10810 5764 10950
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5736 10130 5764 10746
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5828 10062 5856 10610
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5828 9654 5856 9998
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5828 9194 5856 9590
rect 5736 9166 5856 9194
rect 5736 9110 5764 9166
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5460 8078 5580 8106
rect 5264 7336 5316 7342
rect 5078 7304 5134 7313
rect 5264 7278 5316 7284
rect 5078 7239 5134 7248
rect 5000 6956 5120 6984
rect 5092 6916 5120 6956
rect 5000 6888 5120 6916
rect 5170 6896 5226 6905
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 5000 5953 5028 6888
rect 5170 6831 5172 6840
rect 5224 6831 5226 6840
rect 5172 6802 5224 6808
rect 5078 6760 5134 6769
rect 5078 6695 5134 6704
rect 4986 5944 5042 5953
rect 4986 5879 5042 5888
rect 5092 5642 5120 6695
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 4894 4992 4950 5001
rect 4894 4927 4950 4936
rect 4066 4383 4122 4392
rect 4632 4406 4844 4434
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3896 3233 3924 4082
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3976 3664 4028 3670
rect 3974 3632 3976 3641
rect 4028 3632 4030 3641
rect 4632 3618 4660 4406
rect 4710 3904 4766 3913
rect 4710 3839 4766 3848
rect 3974 3567 4030 3576
rect 4540 3590 4660 3618
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3882 3224 3938 3233
rect 3882 3159 3938 3168
rect 4066 3224 4122 3233
rect 4066 3159 4068 3168
rect 4120 3159 4122 3168
rect 4068 3130 4120 3136
rect 4068 3052 4120 3058
rect 3988 3012 4068 3040
rect 3988 2774 4016 3012
rect 4068 2994 4120 3000
rect 4172 2904 4200 3470
rect 4540 3210 4568 3590
rect 4618 3496 4674 3505
rect 4618 3431 4674 3440
rect 4632 3398 4660 3431
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4540 3182 4660 3210
rect 3896 2746 4016 2774
rect 4080 2876 4200 2904
rect 3792 808 3844 814
rect 938 368 994 377
rect 938 303 994 312
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 1950 0 2006 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2870 0 2926 800
rect 3238 0 3294 800
rect 3514 0 3570 800
rect 3896 800 3924 2746
rect 4080 2530 4108 2876
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4080 2502 4200 2530
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4080 2009 4108 2314
rect 4066 2000 4122 2009
rect 4066 1935 4122 1944
rect 4172 898 4200 2502
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 4172 870 4292 898
rect 4172 800 4200 870
rect 3792 750 3844 756
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4264 105 4292 870
rect 4448 800 4476 2382
rect 4632 1193 4660 3182
rect 4724 3126 4752 3839
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4908 3058 4936 4927
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4618 1184 4674 1193
rect 4618 1119 4674 1128
rect 4250 96 4306 105
rect 4250 31 4306 40
rect 4434 0 4490 800
rect 4724 746 4752 2926
rect 5092 2446 5120 3878
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5184 2825 5212 3402
rect 5170 2816 5226 2825
rect 5170 2751 5226 2760
rect 5276 2650 5304 7278
rect 5354 6760 5410 6769
rect 5354 6695 5410 6704
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5368 2514 5396 6695
rect 5460 5302 5488 8078
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5552 7410 5580 7686
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 4486 5488 4966
rect 5552 4593 5580 7346
rect 5644 5574 5672 8434
rect 5920 8362 5948 12294
rect 6012 11257 6040 16934
rect 6104 13530 6132 17138
rect 6196 14346 6224 17614
rect 6274 16824 6330 16833
rect 6274 16759 6330 16768
rect 6288 14550 6316 16759
rect 6380 15978 6408 18022
rect 6472 17678 6500 19230
rect 6644 19178 6696 19184
rect 6550 18592 6606 18601
rect 6550 18527 6606 18536
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6564 16998 6592 18527
rect 6748 17882 6776 19722
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6734 17776 6790 17785
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6368 15972 6420 15978
rect 6368 15914 6420 15920
rect 6472 15337 6500 16050
rect 6656 15502 6684 17750
rect 6734 17711 6736 17720
rect 6788 17711 6790 17720
rect 6736 17682 6788 17688
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6748 16794 6776 16934
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6840 16590 6868 20703
rect 6932 18222 6960 21830
rect 7024 20777 7052 24006
rect 7010 20768 7066 20777
rect 7010 20703 7066 20712
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 6734 16008 6790 16017
rect 6734 15943 6790 15952
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6458 15328 6514 15337
rect 6458 15263 6514 15272
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6458 14512 6514 14521
rect 6458 14447 6514 14456
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 6288 13938 6316 14350
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6104 12986 6132 13466
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6196 12918 6224 13466
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6380 12646 6408 14282
rect 6472 14278 6500 14447
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6472 12850 6500 13942
rect 6564 13705 6592 15370
rect 6748 14822 6776 15943
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6840 14482 6868 15438
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6734 14376 6790 14385
rect 6734 14311 6790 14320
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6550 13696 6606 13705
rect 6550 13631 6606 13640
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6092 12232 6144 12238
rect 6288 12209 6316 12378
rect 6092 12174 6144 12180
rect 6274 12200 6330 12209
rect 5998 11248 6054 11257
rect 5998 11183 6054 11192
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 6012 10146 6040 11018
rect 6104 10266 6132 12174
rect 6274 12135 6330 12144
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6196 10266 6224 11766
rect 6288 11393 6316 12135
rect 6380 11762 6408 12378
rect 6564 12073 6592 13194
rect 6550 12064 6606 12073
rect 6550 11999 6606 12008
rect 6550 11792 6606 11801
rect 6368 11756 6420 11762
rect 6550 11727 6606 11736
rect 6368 11698 6420 11704
rect 6274 11384 6330 11393
rect 6274 11319 6330 11328
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6288 10849 6316 11086
rect 6380 11082 6408 11698
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6472 11098 6500 11562
rect 6564 11218 6592 11727
rect 6656 11354 6684 13874
rect 6748 12850 6776 14311
rect 6840 14006 6868 14418
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6932 13462 6960 15846
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6642 11112 6698 11121
rect 6368 11076 6420 11082
rect 6472 11070 6592 11098
rect 6368 11018 6420 11024
rect 6366 10976 6422 10985
rect 6366 10911 6422 10920
rect 6274 10840 6330 10849
rect 6274 10775 6330 10784
rect 6288 10606 6316 10775
rect 6380 10674 6408 10911
rect 6458 10840 6514 10849
rect 6458 10775 6514 10784
rect 6472 10742 6500 10775
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6012 10118 6132 10146
rect 6104 9625 6132 10118
rect 6090 9616 6146 9625
rect 6000 9580 6052 9586
rect 6090 9551 6146 9560
rect 6000 9522 6052 9528
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 6012 8242 6040 9522
rect 6288 9382 6316 10406
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 9586 6408 9930
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6090 9208 6146 9217
rect 6090 9143 6146 9152
rect 6104 8974 6132 9143
rect 6196 9110 6224 9318
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6182 8936 6238 8945
rect 5920 8214 6040 8242
rect 5814 6624 5870 6633
rect 5814 6559 5870 6568
rect 5828 6458 5856 6559
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 4622 5672 5510
rect 5632 4616 5684 4622
rect 5538 4584 5594 4593
rect 5632 4558 5684 4564
rect 5538 4519 5594 4528
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5736 3942 5764 5578
rect 5920 5574 5948 8214
rect 6104 6866 6132 8910
rect 6182 8871 6184 8880
rect 6236 8871 6238 8880
rect 6184 8842 6236 8848
rect 6182 8392 6238 8401
rect 6182 8327 6238 8336
rect 6196 8090 6224 8327
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6288 7002 6316 9318
rect 6380 7206 6408 9522
rect 6472 9058 6500 9998
rect 6564 9722 6592 11070
rect 6642 11047 6644 11056
rect 6696 11047 6698 11056
rect 6644 11018 6696 11024
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6656 10130 6684 10678
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6656 9217 6684 9930
rect 6642 9208 6698 9217
rect 6748 9178 6776 12582
rect 6840 11694 6868 12854
rect 7024 12434 7052 20538
rect 7116 19718 7144 24550
rect 7208 23526 7236 25094
rect 7196 23520 7248 23526
rect 7196 23462 7248 23468
rect 7196 22976 7248 22982
rect 7196 22918 7248 22924
rect 7208 22506 7236 22918
rect 7196 22500 7248 22506
rect 7196 22442 7248 22448
rect 7194 22128 7250 22137
rect 7194 22063 7250 22072
rect 7208 20074 7236 22063
rect 7300 20874 7328 25094
rect 7484 24834 7512 27610
rect 8036 27130 8064 35974
rect 8680 35494 8708 36722
rect 9404 35556 9456 35562
rect 9404 35498 9456 35504
rect 8668 35488 8720 35494
rect 8668 35430 8720 35436
rect 8484 27328 8536 27334
rect 8484 27270 8536 27276
rect 8024 27124 8076 27130
rect 8024 27066 8076 27072
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 7668 25702 7696 25842
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7564 25492 7616 25498
rect 7564 25434 7616 25440
rect 7392 24806 7512 24834
rect 7288 20868 7340 20874
rect 7288 20810 7340 20816
rect 7208 20046 7328 20074
rect 7300 19922 7328 20046
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7194 19816 7250 19825
rect 7194 19751 7250 19760
rect 7208 19718 7236 19751
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7300 18737 7328 19858
rect 7286 18728 7342 18737
rect 7286 18663 7342 18672
rect 7102 17912 7158 17921
rect 7102 17847 7158 17856
rect 7116 17746 7144 17847
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 7104 17604 7156 17610
rect 7104 17546 7156 17552
rect 7116 17202 7144 17546
rect 7392 17218 7420 24806
rect 7472 24676 7524 24682
rect 7472 24618 7524 24624
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7300 17190 7420 17218
rect 7116 16794 7144 17138
rect 7208 16794 7236 17138
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7116 15026 7144 16730
rect 7194 16552 7250 16561
rect 7194 16487 7250 16496
rect 7208 15502 7236 16487
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 6932 12406 7052 12434
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6642 9143 6698 9152
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6472 9030 6684 9058
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6366 7032 6422 7041
rect 6276 6996 6328 7002
rect 6366 6967 6422 6976
rect 6276 6938 6328 6944
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6104 5574 6132 6802
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 5920 5370 5948 5510
rect 6380 5370 6408 6967
rect 6472 5914 6500 8910
rect 6550 7712 6606 7721
rect 6656 7698 6684 9030
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6748 8090 6776 8910
rect 6840 8566 6868 11630
rect 6932 10033 6960 12406
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7208 12209 7236 12310
rect 7194 12200 7250 12209
rect 7194 12135 7250 12144
rect 7300 11642 7328 17190
rect 7378 16688 7434 16697
rect 7378 16623 7434 16632
rect 7392 16454 7420 16623
rect 7484 16590 7512 24618
rect 7576 22642 7604 25434
rect 7748 24336 7800 24342
rect 7748 24278 7800 24284
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7668 23186 7696 24006
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7760 22778 7788 24278
rect 7932 24132 7984 24138
rect 7932 24074 7984 24080
rect 7944 23798 7972 24074
rect 7932 23792 7984 23798
rect 7932 23734 7984 23740
rect 7930 23488 7986 23497
rect 7930 23423 7986 23432
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7748 22772 7800 22778
rect 7748 22714 7800 22720
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7576 22234 7604 22578
rect 7564 22228 7616 22234
rect 7564 22170 7616 22176
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7576 20602 7604 21966
rect 7564 20596 7616 20602
rect 7564 20538 7616 20544
rect 7654 20360 7710 20369
rect 7654 20295 7710 20304
rect 7562 18184 7618 18193
rect 7562 18119 7618 18128
rect 7576 17377 7604 18119
rect 7562 17368 7618 17377
rect 7562 17303 7618 17312
rect 7562 16688 7618 16697
rect 7562 16623 7618 16632
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7392 15910 7420 16390
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7576 15026 7604 16623
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7668 14906 7696 20295
rect 7852 18358 7880 23190
rect 7944 22642 7972 23423
rect 8036 23118 8064 27066
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 8312 25294 8340 26182
rect 8392 25696 8444 25702
rect 8392 25638 8444 25644
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 8312 24818 8340 25230
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8404 24750 8432 25638
rect 8496 25226 8524 27270
rect 8576 26784 8628 26790
rect 8574 26752 8576 26761
rect 8628 26752 8630 26761
rect 8574 26687 8630 26696
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8484 25220 8536 25226
rect 8484 25162 8536 25168
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8300 24608 8352 24614
rect 8404 24596 8432 24686
rect 8352 24568 8432 24596
rect 8300 24550 8352 24556
rect 8128 24138 8156 24550
rect 8116 24132 8168 24138
rect 8116 24074 8168 24080
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 7932 22636 7984 22642
rect 7932 22578 7984 22584
rect 7932 22024 7984 22030
rect 7930 21992 7932 22001
rect 7984 21992 7986 22001
rect 7930 21927 7986 21936
rect 8036 21486 8064 23054
rect 8128 23050 8156 24074
rect 8312 24041 8340 24550
rect 8298 24032 8354 24041
rect 8298 23967 8354 23976
rect 8312 23526 8340 23967
rect 8300 23520 8352 23526
rect 8300 23462 8352 23468
rect 8312 23322 8340 23462
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8496 23202 8524 25162
rect 8588 24818 8616 25774
rect 8680 24857 8708 35430
rect 9036 27328 9088 27334
rect 9036 27270 9088 27276
rect 9048 27062 9076 27270
rect 9036 27056 9088 27062
rect 9036 26998 9088 27004
rect 8760 26308 8812 26314
rect 8760 26250 8812 26256
rect 8666 24848 8722 24857
rect 8576 24812 8628 24818
rect 8666 24783 8722 24792
rect 8576 24754 8628 24760
rect 8588 24070 8616 24754
rect 8576 24064 8628 24070
rect 8576 24006 8628 24012
rect 8588 23746 8616 24006
rect 8588 23718 8708 23746
rect 8772 23730 8800 26250
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8852 23792 8904 23798
rect 8852 23734 8904 23740
rect 8576 23588 8628 23594
rect 8576 23530 8628 23536
rect 8312 23174 8524 23202
rect 8116 23044 8168 23050
rect 8116 22986 8168 22992
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 8024 21072 8076 21078
rect 8024 21014 8076 21020
rect 7932 20868 7984 20874
rect 7932 20810 7984 20816
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 7944 17610 7972 20810
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 7944 16182 7972 17546
rect 8036 16969 8064 21014
rect 8128 20641 8156 21966
rect 8312 21894 8340 23174
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 8404 21418 8432 22918
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8300 21412 8352 21418
rect 8300 21354 8352 21360
rect 8392 21412 8444 21418
rect 8392 21354 8444 21360
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 8114 20632 8170 20641
rect 8114 20567 8170 20576
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 8022 16960 8078 16969
rect 8022 16895 8078 16904
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7576 14878 7696 14906
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7378 12880 7434 12889
rect 7378 12815 7434 12824
rect 7024 11614 7328 11642
rect 7024 10470 7052 11614
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6918 10024 6974 10033
rect 6918 9959 6974 9968
rect 6918 9616 6974 9625
rect 6918 9551 6974 9560
rect 6932 8566 6960 9551
rect 7024 9081 7052 10406
rect 7116 9110 7144 11494
rect 7392 10690 7420 12815
rect 7484 12374 7512 14010
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7208 10662 7420 10690
rect 7104 9104 7156 9110
rect 7010 9072 7066 9081
rect 7104 9046 7156 9052
rect 7010 9007 7066 9016
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 7024 8498 7052 9007
rect 7102 8936 7158 8945
rect 7102 8871 7158 8880
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7116 8378 7144 8871
rect 7208 8634 7236 10662
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7380 10600 7432 10606
rect 7484 10588 7512 12106
rect 7576 11558 7604 14878
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7668 11393 7696 14758
rect 7760 14521 7788 14962
rect 8128 14929 8156 19178
rect 8220 18834 8248 21286
rect 8312 20942 8340 21354
rect 8404 21146 8432 21354
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8404 20097 8432 20810
rect 8390 20088 8446 20097
rect 8390 20023 8446 20032
rect 8496 19446 8524 21966
rect 8588 19961 8616 23530
rect 8680 22930 8708 23718
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8772 23225 8800 23666
rect 8864 23594 8892 23734
rect 8852 23588 8904 23594
rect 8852 23530 8904 23536
rect 8758 23216 8814 23225
rect 8758 23151 8814 23160
rect 8772 23118 8800 23151
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8864 23050 8892 23530
rect 8852 23044 8904 23050
rect 8852 22986 8904 22992
rect 8680 22902 8892 22930
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8574 19952 8630 19961
rect 8574 19887 8630 19896
rect 8680 19689 8708 22374
rect 8772 19802 8800 22646
rect 8864 21146 8892 22902
rect 8956 21962 8984 24550
rect 9048 24274 9076 25434
rect 9036 24268 9088 24274
rect 9036 24210 9088 24216
rect 9048 23798 9076 24210
rect 9232 24177 9260 25638
rect 9218 24168 9274 24177
rect 9218 24103 9274 24112
rect 9036 23792 9088 23798
rect 9036 23734 9088 23740
rect 9048 23254 9076 23734
rect 9232 23662 9260 24103
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9036 23248 9088 23254
rect 9036 23190 9088 23196
rect 9232 23186 9260 23598
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9034 22944 9090 22953
rect 9034 22879 9090 22888
rect 9048 22642 9076 22879
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 9048 22094 9076 22578
rect 9048 22066 9260 22094
rect 8944 21956 8996 21962
rect 8944 21898 8996 21904
rect 9128 21888 9180 21894
rect 9034 21856 9090 21865
rect 9128 21830 9180 21836
rect 9034 21791 9090 21800
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 8864 20874 8892 21082
rect 8852 20868 8904 20874
rect 8852 20810 8904 20816
rect 8942 20496 8998 20505
rect 8942 20431 8998 20440
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8864 19990 8892 20334
rect 8852 19984 8904 19990
rect 8852 19926 8904 19932
rect 8852 19848 8904 19854
rect 8772 19796 8852 19802
rect 8772 19790 8904 19796
rect 8772 19774 8892 19790
rect 8760 19712 8812 19718
rect 8666 19680 8722 19689
rect 8760 19654 8812 19660
rect 8666 19615 8722 19624
rect 8772 19446 8800 19654
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 8666 18728 8722 18737
rect 8666 18663 8722 18672
rect 8574 18184 8630 18193
rect 8574 18119 8630 18128
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8496 16794 8524 17138
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8220 16454 8248 16662
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8588 16114 8616 18119
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8390 15328 8446 15337
rect 8390 15263 8446 15272
rect 8208 15088 8260 15094
rect 8206 15056 8208 15065
rect 8260 15056 8262 15065
rect 8206 14991 8262 15000
rect 8114 14920 8170 14929
rect 8024 14884 8076 14890
rect 8114 14855 8170 14864
rect 8024 14826 8076 14832
rect 7746 14512 7802 14521
rect 7746 14447 7802 14456
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7760 12170 7788 12650
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7654 11384 7710 11393
rect 7654 11319 7710 11328
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7576 10810 7604 11086
rect 7760 10810 7788 11766
rect 7852 11665 7880 14282
rect 7944 14074 7972 14282
rect 8036 14278 8064 14826
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 7932 13796 7984 13802
rect 7932 13738 7984 13744
rect 7944 13025 7972 13738
rect 7930 13016 7986 13025
rect 7930 12951 7986 12960
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7838 11656 7894 11665
rect 7838 11591 7894 11600
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7484 10560 7604 10588
rect 7380 10542 7432 10548
rect 7300 9994 7328 10542
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7392 9722 7420 10542
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7300 8974 7328 9590
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7288 8968 7340 8974
rect 7392 8945 7420 9522
rect 7484 9382 7512 10202
rect 7576 10010 7604 10560
rect 7760 10130 7788 10746
rect 7944 10130 7972 12786
rect 8036 11218 8064 13942
rect 8220 13394 8248 14010
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8312 13190 8340 14486
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8404 12434 8432 15263
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8496 12918 8524 15098
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8588 13870 8616 14282
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8588 12481 8616 13194
rect 8574 12472 8630 12481
rect 8404 12406 8524 12434
rect 8574 12407 8630 12416
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8128 11898 8156 12310
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8220 10849 8248 12106
rect 8206 10840 8262 10849
rect 8206 10775 8262 10784
rect 8312 10742 8340 12310
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11898 8432 12174
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8022 10296 8078 10305
rect 8022 10231 8078 10240
rect 8036 10130 8064 10231
rect 7748 10124 7800 10130
rect 7932 10124 7984 10130
rect 7800 10084 7880 10112
rect 7748 10066 7800 10072
rect 7576 9982 7788 10010
rect 7760 9926 7788 9982
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7668 9518 7696 9862
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7668 9382 7696 9454
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7484 9178 7512 9318
rect 7760 9217 7788 9862
rect 7852 9450 7880 10084
rect 7932 10066 7984 10072
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8022 10024 8078 10033
rect 8022 9959 8078 9968
rect 8036 9625 8064 9959
rect 8022 9616 8078 9625
rect 7932 9580 7984 9586
rect 8022 9551 8078 9560
rect 8208 9580 8260 9586
rect 7932 9522 7984 9528
rect 8208 9522 8260 9528
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7746 9208 7802 9217
rect 7472 9172 7524 9178
rect 7746 9143 7802 9152
rect 7472 9114 7524 9120
rect 7484 9024 7512 9114
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7840 9104 7892 9110
rect 7944 9092 7972 9522
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7892 9064 7972 9092
rect 7840 9046 7892 9052
rect 7484 8996 7604 9024
rect 7288 8910 7340 8916
rect 7378 8936 7434 8945
rect 7378 8871 7434 8880
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 7024 8350 7144 8378
rect 6932 8090 6960 8298
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6748 7818 6776 8026
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6656 7670 6776 7698
rect 6550 7647 6606 7656
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5828 4282 5856 4966
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 5092 800 5120 2382
rect 5460 898 5488 2994
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5552 2038 5580 2858
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5736 1970 5764 3470
rect 5724 1964 5776 1970
rect 5724 1906 5776 1912
rect 5460 882 5580 898
rect 5460 876 5592 882
rect 5460 870 5540 876
rect 5460 800 5488 870
rect 5540 818 5592 824
rect 5736 800 5764 1906
rect 6104 898 6132 3470
rect 6380 2310 6408 5306
rect 6472 2774 6500 5850
rect 6564 4690 6592 7647
rect 6642 7168 6698 7177
rect 6642 7103 6698 7112
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6656 3738 6684 7103
rect 6748 4690 6776 7670
rect 6840 7410 6868 7822
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6748 3369 6776 3878
rect 6734 3360 6790 3369
rect 6734 3295 6790 3304
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6472 2746 6592 2774
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 6368 1896 6420 1902
rect 6564 1873 6592 2746
rect 6368 1838 6420 1844
rect 6550 1864 6606 1873
rect 6104 870 6224 898
rect 6104 800 6132 870
rect 4712 740 4764 746
rect 4712 682 4764 688
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6196 241 6224 870
rect 6380 800 6408 1838
rect 6550 1799 6606 1808
rect 6748 1170 6776 2994
rect 6932 2922 6960 6666
rect 7024 6610 7052 8350
rect 7208 8276 7236 8434
rect 7116 8248 7236 8276
rect 7116 6798 7144 8248
rect 7194 7984 7250 7993
rect 7194 7919 7250 7928
rect 7208 7886 7236 7919
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7208 6866 7236 7822
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7024 6582 7144 6610
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7024 5302 7052 5510
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 7116 5030 7144 6582
rect 7208 6458 7236 6802
rect 7300 6798 7328 8774
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7392 5642 7420 8366
rect 7484 8090 7512 8842
rect 7576 8090 7604 8996
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7484 7274 7512 8026
rect 7576 7750 7604 8026
rect 7668 7886 7696 9046
rect 8036 9042 8064 9318
rect 8114 9208 8170 9217
rect 8114 9143 8170 9152
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7746 8800 7802 8809
rect 7746 8735 7802 8744
rect 7760 8362 7788 8735
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7654 7304 7710 7313
rect 7472 7268 7524 7274
rect 7654 7239 7710 7248
rect 7472 7210 7524 7216
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7470 6760 7526 6769
rect 7470 6695 7526 6704
rect 7484 6662 7512 6695
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7470 6488 7526 6497
rect 7470 6423 7526 6432
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4146 7420 4966
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7484 3602 7512 6423
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 7010 2680 7066 2689
rect 7010 2615 7066 2624
rect 7024 2446 7052 2615
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 6840 1902 6868 2382
rect 6828 1896 6880 1902
rect 6828 1838 6880 1844
rect 7012 1624 7064 1630
rect 7012 1566 7064 1572
rect 6920 1216 6972 1222
rect 6656 1164 6920 1170
rect 6656 1158 6972 1164
rect 6656 1142 6960 1158
rect 6656 800 6684 1142
rect 7024 800 7052 1566
rect 7288 1080 7340 1086
rect 7288 1022 7340 1028
rect 7300 800 7328 1022
rect 7576 950 7604 6870
rect 7668 3602 7696 7239
rect 7852 6914 7880 8502
rect 8036 8480 8064 8978
rect 8128 8838 8156 9143
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8220 8566 8248 9522
rect 8312 9382 8340 10406
rect 8404 10010 8432 11562
rect 8496 10810 8524 12406
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8680 10538 8708 18663
rect 8864 18086 8892 19774
rect 8956 19514 8984 20431
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 9048 18834 9076 21791
rect 9140 21418 9168 21830
rect 9128 21412 9180 21418
rect 9128 21354 9180 21360
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 9140 20466 9168 20538
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 8942 18456 8998 18465
rect 8942 18391 8998 18400
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8852 17196 8904 17202
rect 8772 17156 8852 17184
rect 8772 15638 8800 17156
rect 8956 17184 8984 18391
rect 9048 18222 9076 18770
rect 9140 18426 9168 19722
rect 9232 18426 9260 22066
rect 9324 21010 9352 23054
rect 9416 21010 9444 35498
rect 9508 35494 9536 36722
rect 9600 36378 9628 37198
rect 9876 36378 9904 37198
rect 10244 36650 10272 39200
rect 10324 37800 10376 37806
rect 10324 37742 10376 37748
rect 10416 37800 10468 37806
rect 10416 37742 10468 37748
rect 10232 36644 10284 36650
rect 10232 36586 10284 36592
rect 9588 36372 9640 36378
rect 9588 36314 9640 36320
rect 9864 36372 9916 36378
rect 9864 36314 9916 36320
rect 10140 36168 10192 36174
rect 10140 36110 10192 36116
rect 10152 35562 10180 36110
rect 10140 35556 10192 35562
rect 10140 35498 10192 35504
rect 9496 35488 9548 35494
rect 9496 35430 9548 35436
rect 9508 28937 9536 35430
rect 9494 28928 9550 28937
rect 9494 28863 9550 28872
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9600 27130 9628 27270
rect 9588 27124 9640 27130
rect 9588 27066 9640 27072
rect 9496 26512 9548 26518
rect 9494 26480 9496 26489
rect 9548 26480 9550 26489
rect 9494 26415 9550 26424
rect 9600 26382 9628 27066
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9600 25498 9628 26318
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 9784 24818 9812 25638
rect 9876 24954 9904 26182
rect 10060 25906 10088 26726
rect 10048 25900 10100 25906
rect 10048 25842 10100 25848
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9588 24336 9640 24342
rect 9588 24278 9640 24284
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9508 21554 9536 23462
rect 9600 22094 9628 24278
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9692 22545 9720 24142
rect 9678 22536 9734 22545
rect 9678 22471 9734 22480
rect 9600 22066 9720 22094
rect 9692 21554 9720 22066
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9784 21185 9812 24754
rect 9876 24426 9904 24890
rect 10060 24886 10088 25842
rect 10140 25832 10192 25838
rect 10140 25774 10192 25780
rect 10048 24880 10100 24886
rect 10048 24822 10100 24828
rect 9956 24608 10008 24614
rect 9954 24576 9956 24585
rect 10008 24576 10010 24585
rect 9954 24511 10010 24520
rect 9876 24398 9996 24426
rect 9864 24336 9916 24342
rect 9864 24278 9916 24284
rect 9876 23186 9904 24278
rect 9968 23882 9996 24398
rect 10060 24313 10088 24822
rect 10046 24304 10102 24313
rect 10046 24239 10102 24248
rect 10060 24138 10088 24239
rect 10152 24138 10180 25774
rect 10048 24132 10100 24138
rect 10048 24074 10100 24080
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 10152 24041 10180 24074
rect 10138 24032 10194 24041
rect 10138 23967 10194 23976
rect 9968 23854 10180 23882
rect 10046 23760 10102 23769
rect 9956 23724 10008 23730
rect 10046 23695 10102 23704
rect 9956 23666 10008 23672
rect 9864 23180 9916 23186
rect 9864 23122 9916 23128
rect 9770 21176 9826 21185
rect 9770 21111 9826 21120
rect 9784 21026 9812 21111
rect 9312 21004 9364 21010
rect 9312 20946 9364 20952
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9692 20998 9812 21026
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8904 17156 8984 17184
rect 8852 17138 8904 17144
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9140 16794 9168 17070
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9324 16658 9352 20402
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 9416 19553 9444 19858
rect 9402 19544 9458 19553
rect 9402 19479 9458 19488
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9034 16552 9090 16561
rect 9034 16487 9090 16496
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8772 13190 8800 15574
rect 8864 15162 8892 16390
rect 8944 16176 8996 16182
rect 8944 16118 8996 16124
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8956 14958 8984 16118
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8956 14618 8984 14894
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8758 12336 8814 12345
rect 8758 12271 8814 12280
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8404 9982 8524 10010
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 7944 8452 8064 8480
rect 7944 7954 7972 8452
rect 8312 8430 8340 8910
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8404 8362 8432 9862
rect 8496 9518 8524 9982
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8482 9208 8538 9217
rect 8482 9143 8538 9152
rect 8666 9208 8722 9217
rect 8666 9143 8722 9152
rect 8496 8974 8524 9143
rect 8680 9110 8708 9143
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8588 8616 8616 8978
rect 8772 8634 8800 12271
rect 8864 11778 8892 13330
rect 8942 12608 8998 12617
rect 8942 12543 8998 12552
rect 8956 12306 8984 12543
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 9048 12102 9076 16487
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9140 16017 9168 16050
rect 9126 16008 9182 16017
rect 9126 15943 9182 15952
rect 9218 15736 9274 15745
rect 9218 15671 9274 15680
rect 9232 14657 9260 15671
rect 9218 14648 9274 14657
rect 9218 14583 9274 14592
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9140 12306 9168 13670
rect 9232 12646 9260 14583
rect 9324 14006 9352 16594
rect 9416 16250 9444 19246
rect 9600 19242 9628 20538
rect 9692 20058 9720 20998
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9784 20466 9812 20810
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9678 19680 9734 19689
rect 9678 19615 9734 19624
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9402 15192 9458 15201
rect 9402 15127 9458 15136
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8864 11750 8984 11778
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8864 9432 8892 11630
rect 8956 11014 8984 11750
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8942 10296 8998 10305
rect 8942 10231 8944 10240
rect 8996 10231 8998 10240
rect 8944 10202 8996 10208
rect 9048 10112 9076 11630
rect 9324 11218 9352 12106
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9140 10577 9168 11018
rect 9310 10840 9366 10849
rect 9310 10775 9366 10784
rect 9126 10568 9182 10577
rect 9126 10503 9182 10512
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 9048 10084 9168 10112
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 9034 10024 9090 10033
rect 8956 9897 8984 9998
rect 9034 9959 9036 9968
rect 9088 9959 9090 9968
rect 9036 9930 9088 9936
rect 8942 9888 8998 9897
rect 8942 9823 8998 9832
rect 9140 9722 9168 10084
rect 9232 9897 9260 10134
rect 9218 9888 9274 9897
rect 9218 9823 9274 9832
rect 9324 9722 9352 10775
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 8864 9404 8984 9432
rect 8850 9344 8906 9353
rect 8850 9279 8906 9288
rect 8760 8628 8812 8634
rect 8588 8588 8708 8616
rect 8680 8480 8708 8588
rect 8760 8570 8812 8576
rect 8588 8452 8708 8480
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7760 6886 7880 6914
rect 7760 6322 7788 6886
rect 7944 6662 7972 7754
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6458 7972 6598
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7944 4486 7972 6394
rect 8036 6186 8064 8230
rect 8128 6322 8156 8298
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8220 8106 8248 8230
rect 8220 8078 8524 8106
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8312 7546 8340 7958
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8220 7041 8248 7346
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8206 7032 8262 7041
rect 8206 6967 8262 6976
rect 8312 6882 8340 7278
rect 8220 6854 8340 6882
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8128 6118 8156 6258
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8220 5914 8248 6854
rect 8298 6760 8354 6769
rect 8298 6695 8354 6704
rect 8312 6662 8340 6695
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 8036 5370 8064 5578
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8404 5234 8432 7686
rect 8496 5710 8524 8078
rect 8588 6934 8616 8452
rect 8668 8356 8720 8362
rect 8864 8344 8892 9279
rect 8956 9024 8984 9404
rect 9140 9353 9168 9658
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9126 9344 9182 9353
rect 9126 9279 9182 9288
rect 9036 9172 9088 9178
rect 9324 9160 9352 9522
rect 9416 9353 9444 15127
rect 9508 14822 9536 18566
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9508 11801 9536 13398
rect 9494 11792 9550 11801
rect 9494 11727 9550 11736
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9508 9518 9536 10678
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9402 9344 9458 9353
rect 9402 9279 9458 9288
rect 9088 9132 9352 9160
rect 9036 9114 9088 9120
rect 9312 9036 9364 9042
rect 8956 8996 9168 9024
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 8668 8298 8720 8304
rect 8772 8316 8892 8344
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 6390 8616 6598
rect 8680 6458 8708 8298
rect 8772 7426 8800 8316
rect 8942 7848 8998 7857
rect 8942 7783 8998 7792
rect 8850 7712 8906 7721
rect 8850 7647 8906 7656
rect 8864 7546 8892 7647
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8772 7398 8892 7426
rect 8956 7410 8984 7783
rect 9048 7721 9076 8842
rect 9140 8430 9168 8996
rect 9312 8978 9364 8984
rect 9324 8498 9352 8978
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9034 7712 9090 7721
rect 9034 7647 9090 7656
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8574 6080 8630 6089
rect 8574 6015 8630 6024
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7760 2122 7788 4082
rect 7944 4078 7972 4422
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7668 2106 7788 2122
rect 7656 2100 7788 2106
rect 7708 2094 7788 2100
rect 7656 2042 7708 2048
rect 7564 944 7616 950
rect 7564 886 7616 892
rect 7668 800 7696 2042
rect 7944 1630 7972 3470
rect 8036 1698 8064 4082
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8312 2650 8340 3538
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8116 2576 8168 2582
rect 8312 2530 8340 2586
rect 8116 2518 8168 2524
rect 8128 1766 8156 2518
rect 8220 2502 8340 2530
rect 8220 2446 8248 2502
rect 8496 2446 8524 3946
rect 8588 3058 8616 6015
rect 8772 5914 8800 6870
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8864 5166 8892 7398
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9140 7002 9168 8230
rect 9416 8022 9444 8910
rect 9508 8498 9536 9454
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9600 8378 9628 18906
rect 9692 18902 9720 19615
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9680 18896 9732 18902
rect 9680 18838 9732 18844
rect 9784 17542 9812 19110
rect 9876 17882 9904 23122
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9784 16658 9812 17478
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9876 14618 9904 17070
rect 9968 15366 9996 23666
rect 10060 23594 10088 23695
rect 10048 23588 10100 23594
rect 10048 23530 10100 23536
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 10060 21894 10088 22986
rect 10152 22420 10180 23854
rect 10244 23050 10272 26726
rect 10336 26042 10364 37742
rect 10428 37466 10456 37742
rect 10416 37460 10468 37466
rect 10416 37402 10468 37408
rect 10704 36922 10732 39200
rect 11072 37262 11100 39200
rect 11152 37868 11204 37874
rect 11152 37810 11204 37816
rect 11060 37256 11112 37262
rect 11060 37198 11112 37204
rect 10692 36916 10744 36922
rect 10692 36858 10744 36864
rect 10968 36780 11020 36786
rect 10968 36722 11020 36728
rect 10876 36712 10928 36718
rect 10876 36654 10928 36660
rect 10784 36576 10836 36582
rect 10784 36518 10836 36524
rect 10796 31754 10824 36518
rect 10888 36038 10916 36654
rect 10876 36032 10928 36038
rect 10876 35974 10928 35980
rect 10888 32473 10916 35974
rect 10980 35494 11008 36722
rect 11072 36378 11100 37198
rect 11060 36372 11112 36378
rect 11060 36314 11112 36320
rect 10968 35488 11020 35494
rect 10968 35430 11020 35436
rect 10980 34610 11008 35430
rect 10968 34604 11020 34610
rect 10968 34546 11020 34552
rect 10874 32464 10930 32473
rect 10874 32399 10930 32408
rect 10704 31726 10824 31754
rect 10414 27704 10470 27713
rect 10414 27639 10470 27648
rect 10428 26586 10456 27639
rect 10508 26920 10560 26926
rect 10508 26862 10560 26868
rect 10416 26580 10468 26586
rect 10416 26522 10468 26528
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10336 23254 10364 25978
rect 10428 23905 10456 26522
rect 10520 26314 10548 26862
rect 10508 26308 10560 26314
rect 10508 26250 10560 26256
rect 10600 26308 10652 26314
rect 10600 26250 10652 26256
rect 10520 25498 10548 26250
rect 10508 25492 10560 25498
rect 10508 25434 10560 25440
rect 10612 24857 10640 26250
rect 10598 24848 10654 24857
rect 10598 24783 10600 24792
rect 10652 24783 10654 24792
rect 10600 24754 10652 24760
rect 10414 23896 10470 23905
rect 10414 23831 10470 23840
rect 10428 23798 10456 23831
rect 10416 23792 10468 23798
rect 10416 23734 10468 23740
rect 10416 23588 10468 23594
rect 10416 23530 10468 23536
rect 10508 23588 10560 23594
rect 10508 23530 10560 23536
rect 10428 23338 10456 23530
rect 10520 23497 10548 23530
rect 10506 23488 10562 23497
rect 10506 23423 10562 23432
rect 10428 23310 10548 23338
rect 10324 23248 10376 23254
rect 10324 23190 10376 23196
rect 10232 23044 10284 23050
rect 10232 22986 10284 22992
rect 10324 22976 10376 22982
rect 10230 22944 10286 22953
rect 10324 22918 10376 22924
rect 10230 22879 10286 22888
rect 10244 22710 10272 22879
rect 10232 22704 10284 22710
rect 10232 22646 10284 22652
rect 10336 22545 10364 22918
rect 10416 22704 10468 22710
rect 10414 22672 10416 22681
rect 10468 22672 10470 22681
rect 10414 22607 10470 22616
rect 10322 22536 10378 22545
rect 10322 22471 10378 22480
rect 10416 22500 10468 22506
rect 10416 22442 10468 22448
rect 10152 22392 10364 22420
rect 10138 22264 10194 22273
rect 10138 22199 10194 22208
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10152 17649 10180 22199
rect 10230 22128 10286 22137
rect 10336 22098 10364 22392
rect 10428 22098 10456 22442
rect 10520 22386 10548 23310
rect 10600 22976 10652 22982
rect 10600 22918 10652 22924
rect 10612 22642 10640 22918
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10520 22358 10640 22386
rect 10230 22063 10286 22072
rect 10324 22092 10376 22098
rect 10244 21350 10272 22063
rect 10324 22034 10376 22040
rect 10416 22092 10468 22098
rect 10416 22034 10468 22040
rect 10322 21992 10378 22001
rect 10322 21927 10378 21936
rect 10336 21690 10364 21927
rect 10612 21894 10640 22358
rect 10704 22098 10732 31726
rect 10876 27940 10928 27946
rect 10876 27882 10928 27888
rect 10888 26790 10916 27882
rect 11060 27872 11112 27878
rect 11060 27814 11112 27820
rect 10968 27328 11020 27334
rect 10968 27270 11020 27276
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10980 24721 11008 27270
rect 11072 24954 11100 27814
rect 11164 25498 11192 37810
rect 11440 36922 11468 39200
rect 11428 36916 11480 36922
rect 11428 36858 11480 36864
rect 11900 36378 11928 39200
rect 12268 37330 12296 39200
rect 12440 37732 12492 37738
rect 12440 37674 12492 37680
rect 12256 37324 12308 37330
rect 12256 37266 12308 37272
rect 11980 36780 12032 36786
rect 11980 36722 12032 36728
rect 11888 36372 11940 36378
rect 11888 36314 11940 36320
rect 11992 35494 12020 36722
rect 12256 35556 12308 35562
rect 12256 35498 12308 35504
rect 11980 35488 12032 35494
rect 11980 35430 12032 35436
rect 11992 34542 12020 35430
rect 11980 34536 12032 34542
rect 11980 34478 12032 34484
rect 11336 26988 11388 26994
rect 11336 26930 11388 26936
rect 11152 25492 11204 25498
rect 11152 25434 11204 25440
rect 11060 24948 11112 24954
rect 11060 24890 11112 24896
rect 10966 24712 11022 24721
rect 11022 24670 11100 24698
rect 10966 24647 11022 24656
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 10784 23180 10836 23186
rect 10784 23122 10836 23128
rect 10796 22760 10824 23122
rect 10888 22982 10916 23666
rect 10968 23248 11020 23254
rect 10968 23190 11020 23196
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10876 22772 10928 22778
rect 10796 22732 10876 22760
rect 10876 22714 10928 22720
rect 10782 22672 10838 22681
rect 10782 22607 10784 22616
rect 10836 22607 10838 22616
rect 10784 22578 10836 22584
rect 10796 22438 10824 22578
rect 10876 22500 10928 22506
rect 10876 22442 10928 22448
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10796 22137 10824 22170
rect 10782 22128 10838 22137
rect 10692 22092 10744 22098
rect 10782 22063 10838 22072
rect 10692 22034 10744 22040
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10324 21684 10376 21690
rect 10324 21626 10376 21632
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 10138 17640 10194 17649
rect 10138 17575 10194 17584
rect 10140 16720 10192 16726
rect 10244 16697 10272 21286
rect 10428 20398 10456 21354
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10322 19544 10378 19553
rect 10322 19479 10378 19488
rect 10140 16662 10192 16668
rect 10230 16688 10286 16697
rect 10152 16130 10180 16662
rect 10230 16623 10286 16632
rect 10244 16522 10272 16623
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 10152 16102 10272 16130
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9864 13864 9916 13870
rect 9862 13832 9864 13841
rect 9916 13832 9918 13841
rect 9680 13796 9732 13802
rect 9862 13767 9918 13776
rect 9680 13738 9732 13744
rect 9692 13530 9720 13738
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9678 13424 9734 13433
rect 9678 13359 9734 13368
rect 9692 12986 9720 13359
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9968 12850 9996 15302
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9862 12472 9918 12481
rect 9862 12407 9918 12416
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9692 8906 9720 11154
rect 9784 11121 9812 11494
rect 9770 11112 9826 11121
rect 9770 11047 9826 11056
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9784 9722 9812 10474
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9600 8350 9720 8378
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9494 7984 9550 7993
rect 9494 7919 9550 7928
rect 9508 7868 9536 7919
rect 9416 7840 9536 7868
rect 9416 7256 9444 7840
rect 9588 7744 9640 7750
rect 9494 7712 9550 7721
rect 9588 7686 9640 7692
rect 9494 7647 9550 7656
rect 9508 7546 9536 7647
rect 9600 7585 9628 7686
rect 9586 7576 9642 7585
rect 9496 7540 9548 7546
rect 9586 7511 9642 7520
rect 9496 7482 9548 7488
rect 9496 7268 9548 7274
rect 9416 7228 9496 7256
rect 9496 7210 9548 7216
rect 9494 7032 9550 7041
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9220 6996 9272 7002
rect 9494 6967 9550 6976
rect 9220 6938 9272 6944
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 9048 5030 9076 6258
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8956 4457 8984 4762
rect 9048 4622 9076 4966
rect 9126 4856 9182 4865
rect 9126 4791 9128 4800
rect 9180 4791 9182 4800
rect 9128 4762 9180 4768
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8942 4448 8998 4457
rect 8942 4383 8998 4392
rect 9232 4010 9260 6938
rect 9402 6896 9458 6905
rect 9402 6831 9404 6840
rect 9456 6831 9458 6840
rect 9404 6802 9456 6808
rect 9310 6216 9366 6225
rect 9310 6151 9366 6160
rect 9324 4826 9352 6151
rect 9402 5944 9458 5953
rect 9402 5879 9404 5888
rect 9456 5879 9458 5888
rect 9404 5850 9456 5856
rect 9312 4820 9364 4826
rect 9508 4808 9536 6967
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9600 6769 9628 6802
rect 9586 6760 9642 6769
rect 9586 6695 9642 6704
rect 9586 6216 9642 6225
rect 9586 6151 9642 6160
rect 9312 4762 9364 4768
rect 9416 4780 9536 4808
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8208 2440 8260 2446
rect 8484 2440 8536 2446
rect 8208 2382 8260 2388
rect 8312 2400 8484 2428
rect 8116 1760 8168 1766
rect 8116 1702 8168 1708
rect 8024 1692 8076 1698
rect 8024 1634 8076 1640
rect 7932 1624 7984 1630
rect 7932 1566 7984 1572
rect 8036 1442 8064 1634
rect 7944 1414 8064 1442
rect 7944 800 7972 1414
rect 8312 800 8340 2400
rect 8484 2382 8536 2388
rect 8588 800 8616 2586
rect 8864 1086 8892 2926
rect 8852 1080 8904 1086
rect 8852 1022 8904 1028
rect 8956 898 8984 2994
rect 9324 898 9352 3470
rect 9416 2774 9444 4780
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9508 4282 9536 4626
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9494 3768 9550 3777
rect 9494 3703 9496 3712
rect 9548 3703 9550 3712
rect 9496 3674 9548 3680
rect 9600 2854 9628 6151
rect 9692 5545 9720 8350
rect 9784 7002 9812 9522
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9770 6352 9826 6361
rect 9770 6287 9772 6296
rect 9824 6287 9826 6296
rect 9772 6258 9824 6264
rect 9772 5568 9824 5574
rect 9678 5536 9734 5545
rect 9772 5510 9824 5516
rect 9678 5471 9734 5480
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9692 3058 9720 4218
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9416 2746 9536 2774
rect 9508 2650 9536 2746
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9784 2553 9812 5510
rect 9876 5370 9904 12407
rect 9954 11248 10010 11257
rect 9954 11183 10010 11192
rect 9968 9897 9996 11183
rect 9954 9888 10010 9897
rect 9954 9823 10010 9832
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9968 9110 9996 9658
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9968 8537 9996 8570
rect 9954 8528 10010 8537
rect 9954 8463 10010 8472
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9968 8265 9996 8366
rect 9954 8256 10010 8265
rect 9954 8191 10010 8200
rect 9954 8120 10010 8129
rect 9954 8055 9956 8064
rect 10008 8055 10010 8064
rect 9956 8026 10008 8032
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9968 6730 9996 7890
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 9968 6633 9996 6666
rect 9954 6624 10010 6633
rect 9954 6559 10010 6568
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9968 3738 9996 6559
rect 10060 6458 10088 14282
rect 10152 10742 10180 15846
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10152 10198 10180 10678
rect 10244 10577 10272 16102
rect 10336 13705 10364 19479
rect 10428 18698 10456 20334
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10520 18630 10548 21830
rect 10612 18834 10640 21830
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10704 21146 10732 21490
rect 10782 21448 10838 21457
rect 10782 21383 10838 21392
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10796 20942 10824 21383
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10782 20496 10838 20505
rect 10692 20460 10744 20466
rect 10782 20431 10838 20440
rect 10692 20402 10744 20408
rect 10704 20058 10732 20402
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10690 19816 10746 19825
rect 10690 19751 10746 19760
rect 10704 19553 10732 19751
rect 10690 19544 10746 19553
rect 10690 19479 10746 19488
rect 10690 19408 10746 19417
rect 10690 19343 10746 19352
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10428 13870 10456 16934
rect 10520 14006 10548 17682
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 10612 16998 10640 17274
rect 10704 17270 10732 19343
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10322 13696 10378 13705
rect 10322 13631 10378 13640
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10336 11830 10364 12922
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10428 10674 10456 13194
rect 10520 12458 10548 13942
rect 10612 13870 10640 16934
rect 10690 16824 10746 16833
rect 10690 16759 10746 16768
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10598 13016 10654 13025
rect 10598 12951 10654 12960
rect 10612 12782 10640 12951
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10520 12430 10640 12458
rect 10506 12336 10562 12345
rect 10506 12271 10562 12280
rect 10520 11762 10548 12271
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10520 11558 10548 11698
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10612 10810 10640 12430
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10230 10568 10286 10577
rect 10230 10503 10286 10512
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 10232 9512 10284 9518
rect 10152 9460 10232 9466
rect 10152 9454 10284 9460
rect 10152 9438 10272 9454
rect 10152 9081 10180 9438
rect 10232 9104 10284 9110
rect 10138 9072 10194 9081
rect 10232 9046 10284 9052
rect 10138 9007 10194 9016
rect 10152 8974 10180 9007
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10152 7206 10180 8434
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10244 6662 10272 9046
rect 10336 7886 10364 9687
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10428 7698 10456 9998
rect 10520 9722 10548 10746
rect 10600 10260 10652 10266
rect 10704 10248 10732 16759
rect 10796 16046 10824 20431
rect 10888 19242 10916 22442
rect 10980 22234 11008 23190
rect 11072 22506 11100 24670
rect 11060 22500 11112 22506
rect 11060 22442 11112 22448
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 11164 22166 11192 25434
rect 11244 25424 11296 25430
rect 11244 25366 11296 25372
rect 11152 22160 11204 22166
rect 11058 22128 11114 22137
rect 11152 22102 11204 22108
rect 11058 22063 11114 22072
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10876 19236 10928 19242
rect 10876 19178 10928 19184
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 10888 17678 10916 18634
rect 10980 18601 11008 21830
rect 11072 19922 11100 22063
rect 11152 20392 11204 20398
rect 11152 20334 11204 20340
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 10966 18592 11022 18601
rect 10966 18527 11022 18536
rect 11072 18086 11100 18634
rect 11164 18154 11192 20334
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11256 17882 11284 25366
rect 11348 25294 11376 26930
rect 11520 26852 11572 26858
rect 11520 26794 11572 26800
rect 11704 26852 11756 26858
rect 11704 26794 11756 26800
rect 11532 26518 11560 26794
rect 11520 26512 11572 26518
rect 11520 26454 11572 26460
rect 11520 25696 11572 25702
rect 11518 25664 11520 25673
rect 11572 25664 11574 25673
rect 11518 25599 11574 25608
rect 11428 25492 11480 25498
rect 11428 25434 11480 25440
rect 11336 25288 11388 25294
rect 11336 25230 11388 25236
rect 11440 25129 11468 25434
rect 11426 25120 11482 25129
rect 11426 25055 11482 25064
rect 11518 24984 11574 24993
rect 11518 24919 11574 24928
rect 11532 24410 11560 24919
rect 11612 24676 11664 24682
rect 11612 24618 11664 24624
rect 11520 24404 11572 24410
rect 11520 24346 11572 24352
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11348 23866 11376 24142
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11348 22681 11376 23190
rect 11334 22672 11390 22681
rect 11334 22607 11390 22616
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11348 21146 11376 21626
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11334 18864 11390 18873
rect 11334 18799 11390 18808
rect 11348 18290 11376 18799
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11440 18154 11468 24006
rect 11624 23866 11652 24618
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11716 23798 11744 26794
rect 12072 26376 12124 26382
rect 12072 26318 12124 26324
rect 12084 26042 12112 26318
rect 12072 26036 12124 26042
rect 12072 25978 12124 25984
rect 12084 25770 12112 25978
rect 12072 25764 12124 25770
rect 12072 25706 12124 25712
rect 11888 25288 11940 25294
rect 11888 25230 11940 25236
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11704 23792 11756 23798
rect 11704 23734 11756 23740
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11532 23186 11560 23530
rect 11610 23352 11666 23361
rect 11610 23287 11666 23296
rect 11520 23180 11572 23186
rect 11520 23122 11572 23128
rect 11532 20534 11560 23122
rect 11624 21962 11652 23287
rect 11612 21956 11664 21962
rect 11612 21898 11664 21904
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11624 21078 11652 21626
rect 11716 21593 11744 23734
rect 11808 22982 11836 24074
rect 11796 22976 11848 22982
rect 11796 22918 11848 22924
rect 11808 21706 11836 22918
rect 11900 22658 11928 25230
rect 12164 24608 12216 24614
rect 12164 24550 12216 24556
rect 12072 24404 12124 24410
rect 12072 24346 12124 24352
rect 12084 24206 12112 24346
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12084 23730 12112 24142
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11992 22778 12020 23598
rect 12176 23361 12204 24550
rect 12162 23352 12218 23361
rect 12162 23287 12218 23296
rect 12164 23248 12216 23254
rect 12164 23190 12216 23196
rect 12176 22778 12204 23190
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 11900 22630 12204 22658
rect 11888 22500 11940 22506
rect 11888 22442 11940 22448
rect 11900 22094 11928 22442
rect 11900 22066 12020 22094
rect 11888 21888 11940 21894
rect 11886 21856 11888 21865
rect 11940 21856 11942 21865
rect 11886 21791 11942 21800
rect 11808 21678 11928 21706
rect 11796 21616 11848 21622
rect 11702 21584 11758 21593
rect 11796 21558 11848 21564
rect 11702 21519 11758 21528
rect 11612 21072 11664 21078
rect 11612 21014 11664 21020
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11532 18834 11560 19246
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11336 18148 11388 18154
rect 11336 18090 11388 18096
rect 11428 18148 11480 18154
rect 11428 18090 11480 18096
rect 11348 17921 11376 18090
rect 11334 17912 11390 17921
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11244 17876 11296 17882
rect 11334 17847 11390 17856
rect 11244 17818 11296 17824
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10888 16726 10916 17614
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 10874 16552 10930 16561
rect 10874 16487 10930 16496
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10888 15892 10916 16487
rect 10796 15864 10916 15892
rect 10796 14872 10824 15864
rect 10874 15736 10930 15745
rect 10874 15671 10930 15680
rect 10888 15570 10916 15671
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10796 14844 10916 14872
rect 10782 14512 10838 14521
rect 10782 14447 10838 14456
rect 10796 14414 10824 14447
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10796 13977 10824 14350
rect 10782 13968 10838 13977
rect 10782 13903 10838 13912
rect 10888 13734 10916 14844
rect 11072 14226 11100 17818
rect 11348 17762 11376 17847
rect 11256 17734 11376 17762
rect 11150 17096 11206 17105
rect 11150 17031 11206 17040
rect 11164 15502 11192 17031
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11256 15162 11284 17734
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11334 16416 11390 16425
rect 11334 16351 11390 16360
rect 11348 16250 11376 16351
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11440 15434 11468 17546
rect 11532 16658 11560 18770
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11624 16522 11652 20810
rect 11716 20602 11744 21519
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11808 19922 11836 21558
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 11702 18592 11758 18601
rect 11702 18527 11758 18536
rect 11612 16516 11664 16522
rect 11612 16458 11664 16464
rect 11610 16280 11666 16289
rect 11610 16215 11612 16224
rect 11664 16215 11666 16224
rect 11612 16186 11664 16192
rect 11624 15570 11652 16186
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11428 15428 11480 15434
rect 11428 15370 11480 15376
rect 11716 15201 11744 18527
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11702 15192 11758 15201
rect 11244 15156 11296 15162
rect 11702 15127 11758 15136
rect 11244 15098 11296 15104
rect 11610 14920 11666 14929
rect 11610 14855 11612 14864
rect 11664 14855 11666 14864
rect 11612 14826 11664 14832
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11164 14346 11192 14486
rect 11244 14408 11296 14414
rect 11520 14408 11572 14414
rect 11244 14350 11296 14356
rect 11440 14368 11520 14396
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11072 14198 11192 14226
rect 11058 14104 11114 14113
rect 11058 14039 11114 14048
rect 11072 14006 11100 14039
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 11164 13802 11192 14198
rect 11256 13870 11284 14350
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10796 11014 10824 13262
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12889 10916 13194
rect 10874 12880 10930 12889
rect 10874 12815 10930 12824
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10782 10704 10838 10713
rect 10782 10639 10838 10648
rect 10652 10220 10732 10248
rect 10600 10202 10652 10208
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10336 7670 10456 7698
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10048 6452 10100 6458
rect 10336 6440 10364 7670
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10048 6394 10100 6400
rect 10152 6412 10364 6440
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10060 3670 10088 6258
rect 10152 5370 10180 6412
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10230 6216 10286 6225
rect 10230 6151 10286 6160
rect 10244 6118 10272 6151
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10232 5704 10284 5710
rect 10230 5672 10232 5681
rect 10284 5672 10286 5681
rect 10230 5607 10286 5616
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10152 4593 10180 5306
rect 10232 5296 10284 5302
rect 10336 5284 10364 6258
rect 10284 5256 10364 5284
rect 10232 5238 10284 5244
rect 10428 4758 10456 7414
rect 10520 7041 10548 8910
rect 10612 8634 10640 9930
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10704 8514 10732 9658
rect 10796 9110 10824 10639
rect 10888 9382 10916 10746
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10784 9104 10836 9110
rect 10784 9046 10836 9052
rect 10888 8673 10916 9318
rect 10980 9042 11008 12310
rect 11072 10305 11100 12786
rect 11164 12714 11192 13738
rect 11256 13326 11284 13806
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11058 10296 11114 10305
rect 11058 10231 11114 10240
rect 11164 10169 11192 12106
rect 11256 11694 11284 13262
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11348 11937 11376 12582
rect 11440 12481 11468 14368
rect 11520 14350 11572 14356
rect 11518 14240 11574 14249
rect 11518 14175 11574 14184
rect 11426 12472 11482 12481
rect 11426 12407 11482 12416
rect 11334 11928 11390 11937
rect 11334 11863 11390 11872
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11256 11150 11284 11630
rect 11532 11558 11560 14175
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11426 11248 11482 11257
rect 11426 11183 11482 11192
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11334 11112 11390 11121
rect 11256 10606 11284 11086
rect 11334 11047 11390 11056
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11150 10160 11206 10169
rect 11150 10095 11206 10104
rect 11348 9194 11376 11047
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11164 9166 11376 9194
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 11072 8673 11100 9114
rect 10874 8664 10930 8673
rect 10874 8599 10930 8608
rect 11058 8664 11114 8673
rect 11058 8599 11114 8608
rect 10612 8486 10732 8514
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10874 8528 10930 8537
rect 10506 7032 10562 7041
rect 10612 7002 10640 8486
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10506 6967 10562 6976
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10704 6866 10732 7890
rect 10796 7886 10824 8502
rect 11164 8514 11192 9166
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 10874 8463 10930 8472
rect 10980 8486 11192 8514
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 7449 10824 7686
rect 10782 7440 10838 7449
rect 10782 7375 10838 7384
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10506 6760 10562 6769
rect 10704 6730 10732 6802
rect 10506 6695 10562 6704
rect 10692 6724 10744 6730
rect 10520 6390 10548 6695
rect 10692 6666 10744 6672
rect 10598 6624 10654 6633
rect 10598 6559 10654 6568
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10520 4826 10548 6326
rect 10612 5914 10640 6559
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10600 5704 10652 5710
rect 10598 5672 10600 5681
rect 10652 5672 10654 5681
rect 10598 5607 10654 5616
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10138 4584 10194 4593
rect 10138 4519 10194 4528
rect 10520 4298 10548 4762
rect 10428 4270 10548 4298
rect 10428 4214 10456 4270
rect 10704 4214 10732 6258
rect 10796 5370 10824 7278
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10784 5160 10836 5166
rect 10782 5128 10784 5137
rect 10836 5128 10838 5137
rect 10782 5063 10838 5072
rect 10782 4584 10838 4593
rect 10782 4519 10838 4528
rect 10416 4208 10468 4214
rect 10692 4208 10744 4214
rect 10416 4150 10468 4156
rect 10506 4176 10562 4185
rect 10692 4150 10744 4156
rect 10506 4111 10562 4120
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10520 3058 10548 4111
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9770 2544 9826 2553
rect 9588 2508 9640 2514
rect 9770 2479 9826 2488
rect 9588 2450 9640 2456
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 8864 870 8984 898
rect 9232 870 9352 898
rect 8864 800 8892 870
rect 9232 800 9260 870
rect 6182 232 6238 241
rect 6182 167 6238 176
rect 6366 0 6422 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9324 762 9352 870
rect 9508 800 9536 2382
rect 9600 2281 9628 2450
rect 9586 2272 9642 2281
rect 9586 2207 9642 2216
rect 9876 800 9904 2926
rect 10138 2544 10194 2553
rect 10138 2479 10140 2488
rect 10192 2479 10194 2488
rect 10140 2450 10192 2456
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10152 800 10180 2246
rect 10612 898 10640 3470
rect 10796 3058 10824 4519
rect 10888 3738 10916 8463
rect 10980 6934 11008 8486
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 11072 6458 11100 8366
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11164 7177 11192 7822
rect 11150 7168 11206 7177
rect 11150 7103 11206 7112
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11072 6202 11100 6258
rect 10980 6174 11100 6202
rect 10980 5545 11008 6174
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5953 11100 6054
rect 11058 5944 11114 5953
rect 11058 5879 11114 5888
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 10966 5536 11022 5545
rect 10966 5471 11022 5480
rect 11072 5098 11100 5782
rect 11164 5273 11192 6598
rect 11150 5264 11206 5273
rect 11150 5199 11206 5208
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 11256 4826 11284 8842
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11348 6066 11376 8774
rect 11440 8634 11468 11183
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11532 10062 11560 10542
rect 11624 10266 11652 10610
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11518 9888 11574 9897
rect 11518 9823 11574 9832
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11532 7954 11560 9823
rect 11610 9616 11666 9625
rect 11610 9551 11666 9560
rect 11624 9518 11652 9551
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11624 9042 11652 9454
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11716 8922 11744 13126
rect 11808 11830 11836 17206
rect 11900 12374 11928 21678
rect 11992 21350 12020 22066
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 12084 21486 12112 21966
rect 12176 21554 12204 22630
rect 12268 21622 12296 35498
rect 12452 30546 12480 37674
rect 12636 37126 12664 39200
rect 12716 38004 12768 38010
rect 12716 37946 12768 37952
rect 12728 37398 12756 37946
rect 12716 37392 12768 37398
rect 12716 37334 12768 37340
rect 12624 37120 12676 37126
rect 12624 37062 12676 37068
rect 13096 36922 13124 39200
rect 13464 37330 13492 39200
rect 13452 37324 13504 37330
rect 13452 37266 13504 37272
rect 13360 37256 13412 37262
rect 13360 37198 13412 37204
rect 13084 36916 13136 36922
rect 13084 36858 13136 36864
rect 12624 36780 12676 36786
rect 12624 36722 12676 36728
rect 12636 35494 12664 36722
rect 13176 36168 13228 36174
rect 13176 36110 13228 36116
rect 13188 35494 13216 36110
rect 12624 35488 12676 35494
rect 12624 35430 12676 35436
rect 13176 35488 13228 35494
rect 13176 35430 13228 35436
rect 12636 31754 12664 35430
rect 12992 34604 13044 34610
rect 12992 34546 13044 34552
rect 12636 31726 12756 31754
rect 12452 30518 12664 30546
rect 12636 26518 12664 30518
rect 12728 27033 12756 31726
rect 12714 27024 12770 27033
rect 12714 26959 12770 26968
rect 12624 26512 12676 26518
rect 12622 26480 12624 26489
rect 12676 26480 12678 26489
rect 12622 26415 12678 26424
rect 12714 25936 12770 25945
rect 12714 25871 12770 25880
rect 12530 25664 12586 25673
rect 12530 25599 12586 25608
rect 12544 25498 12572 25599
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12624 25424 12676 25430
rect 12624 25366 12676 25372
rect 12440 25356 12492 25362
rect 12440 25298 12492 25304
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 12360 24886 12388 25094
rect 12348 24880 12400 24886
rect 12348 24822 12400 24828
rect 12360 23798 12388 24822
rect 12348 23792 12400 23798
rect 12348 23734 12400 23740
rect 12348 23520 12400 23526
rect 12346 23488 12348 23497
rect 12400 23488 12402 23497
rect 12346 23423 12402 23432
rect 12348 23112 12400 23118
rect 12452 23100 12480 25298
rect 12530 25256 12586 25265
rect 12530 25191 12586 25200
rect 12400 23072 12480 23100
rect 12348 23054 12400 23060
rect 12346 22944 12402 22953
rect 12346 22879 12402 22888
rect 12360 22030 12388 22879
rect 12452 22642 12480 23072
rect 12544 22953 12572 25191
rect 12530 22944 12586 22953
rect 12530 22879 12586 22888
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12438 22128 12494 22137
rect 12438 22063 12494 22072
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12452 21876 12480 22063
rect 12360 21848 12480 21876
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 12164 21412 12216 21418
rect 12164 21354 12216 21360
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 12084 20777 12112 20878
rect 12070 20768 12126 20777
rect 12070 20703 12126 20712
rect 12176 18873 12204 21354
rect 12360 19938 12388 21848
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12268 19910 12388 19938
rect 12162 18864 12218 18873
rect 12162 18799 12218 18808
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11992 16402 12020 18362
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 12084 16590 12112 17818
rect 12176 17746 12204 18090
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12268 17338 12296 19910
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12360 18034 12388 19790
rect 12452 18222 12480 21490
rect 12544 20777 12572 22714
rect 12636 22658 12664 25366
rect 12728 23594 12756 25871
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12716 23588 12768 23594
rect 12716 23530 12768 23536
rect 12820 22982 12848 24550
rect 12898 23624 12954 23633
rect 12898 23559 12900 23568
rect 12952 23559 12954 23568
rect 12900 23530 12952 23536
rect 12900 23248 12952 23254
rect 12900 23190 12952 23196
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12820 22778 12848 22918
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 12636 22630 12848 22658
rect 12912 22642 12940 23190
rect 12624 22500 12676 22506
rect 12624 22442 12676 22448
rect 12636 21962 12664 22442
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12728 22030 12756 22374
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12624 21956 12676 21962
rect 12624 21898 12676 21904
rect 12636 21690 12664 21898
rect 12820 21894 12848 22630
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 12912 22001 12940 22102
rect 12898 21992 12954 22001
rect 12898 21927 12954 21936
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12530 20768 12586 20777
rect 12530 20703 12586 20712
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12360 18006 12572 18034
rect 12438 17776 12494 17785
rect 12438 17711 12440 17720
rect 12492 17711 12494 17720
rect 12440 17682 12492 17688
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12360 17270 12388 17546
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12544 17066 12572 18006
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12452 16658 12480 17002
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 11992 16374 12112 16402
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11992 14006 12020 14282
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11886 11520 11942 11529
rect 11886 11455 11942 11464
rect 11900 10690 11928 11455
rect 11992 10810 12020 12650
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11900 10662 12020 10690
rect 11886 10024 11942 10033
rect 11796 9988 11848 9994
rect 11886 9959 11942 9968
rect 11796 9930 11848 9936
rect 11808 9489 11836 9930
rect 11794 9480 11850 9489
rect 11794 9415 11850 9424
rect 11900 9382 11928 9959
rect 11992 9761 12020 10662
rect 11978 9752 12034 9761
rect 11978 9687 12034 9696
rect 11978 9616 12034 9625
rect 11978 9551 12034 9560
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11992 9178 12020 9551
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11624 8906 11744 8922
rect 11612 8900 11744 8906
rect 11664 8894 11744 8900
rect 11796 8900 11848 8906
rect 11612 8842 11664 8848
rect 11796 8842 11848 8848
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11428 7744 11480 7750
rect 11426 7712 11428 7721
rect 11480 7712 11482 7721
rect 11426 7647 11482 7656
rect 11532 7585 11560 7890
rect 11808 7834 11836 8842
rect 11716 7806 11836 7834
rect 11518 7576 11574 7585
rect 11518 7511 11574 7520
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11428 7200 11480 7206
rect 11426 7168 11428 7177
rect 11480 7168 11482 7177
rect 11426 7103 11482 7112
rect 11348 6038 11468 6066
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11348 5817 11376 5850
rect 11334 5808 11390 5817
rect 11334 5743 11390 5752
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11150 3224 11206 3233
rect 11150 3159 11206 3168
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10784 1148 10836 1154
rect 10784 1090 10836 1096
rect 10520 870 10640 898
rect 10520 800 10548 870
rect 9324 734 9444 762
rect 9416 406 9444 734
rect 9404 400 9456 406
rect 9404 342 9456 348
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10612 762 10640 870
rect 10796 800 10824 1090
rect 11072 800 11100 2790
rect 11164 2582 11192 3159
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11256 1154 11284 3470
rect 11348 2774 11376 5034
rect 11440 4214 11468 6038
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11440 3738 11468 4014
rect 11532 3738 11560 7346
rect 11610 7304 11666 7313
rect 11610 7239 11612 7248
rect 11664 7239 11666 7248
rect 11612 7210 11664 7216
rect 11610 7168 11666 7177
rect 11610 7103 11666 7112
rect 11624 6322 11652 7103
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11624 4214 11652 5578
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11716 3670 11744 7806
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 5914 11836 7686
rect 11992 7426 12020 8978
rect 12084 8090 12112 16374
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12268 14074 12296 15030
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12360 13818 12388 15438
rect 12636 14550 12664 21422
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12728 21010 12756 21082
rect 12716 21004 12768 21010
rect 12716 20946 12768 20952
rect 12808 20936 12860 20942
rect 12808 20878 12860 20884
rect 12820 19689 12848 20878
rect 12806 19680 12862 19689
rect 12806 19615 12862 19624
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12728 14940 12756 18566
rect 12820 16561 12848 19615
rect 12806 16552 12862 16561
rect 12806 16487 12862 16496
rect 12912 15094 12940 21830
rect 13004 20466 13032 34546
rect 13188 30569 13216 35430
rect 13268 34536 13320 34542
rect 13268 34478 13320 34484
rect 13174 30560 13230 30569
rect 13174 30495 13230 30504
rect 13082 26344 13138 26353
rect 13082 26279 13084 26288
rect 13136 26279 13138 26288
rect 13084 26250 13136 26256
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 13096 25265 13124 25638
rect 13082 25256 13138 25265
rect 13082 25191 13138 25200
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 13096 23322 13124 23666
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 13188 22710 13216 24346
rect 13176 22704 13228 22710
rect 13176 22646 13228 22652
rect 13174 22536 13230 22545
rect 13174 22471 13230 22480
rect 13082 22400 13138 22409
rect 13082 22335 13138 22344
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 12990 19680 13046 19689
rect 12990 19615 13046 19624
rect 13004 18154 13032 19615
rect 12992 18148 13044 18154
rect 12992 18090 13044 18096
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13004 16114 13032 16526
rect 13096 16182 13124 22335
rect 13188 21894 13216 22471
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 13174 21720 13230 21729
rect 13174 21655 13176 21664
rect 13228 21655 13230 21664
rect 13176 21626 13228 21632
rect 13174 21448 13230 21457
rect 13174 21383 13176 21392
rect 13228 21383 13230 21392
rect 13176 21354 13228 21360
rect 13174 21312 13230 21321
rect 13174 21247 13230 21256
rect 13188 20942 13216 21247
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13188 18630 13216 20742
rect 13280 19922 13308 34478
rect 13372 30433 13400 37198
rect 13464 36378 13492 37266
rect 13924 36922 13952 39200
rect 13912 36916 13964 36922
rect 13912 36858 13964 36864
rect 13728 36780 13780 36786
rect 13728 36722 13780 36728
rect 13452 36372 13504 36378
rect 13452 36314 13504 36320
rect 13740 34649 13768 36722
rect 14292 36378 14320 39200
rect 14660 39114 14688 39200
rect 14752 39114 14780 39222
rect 14660 39086 14780 39114
rect 15028 36802 15056 39222
rect 15106 39200 15162 40000
rect 15474 39200 15530 40000
rect 15934 39200 15990 40000
rect 16302 39200 16358 40000
rect 16670 39200 16726 40000
rect 17130 39200 17186 40000
rect 17498 39200 17554 40000
rect 17866 39200 17922 40000
rect 18326 39200 18382 40000
rect 18694 39200 18750 40000
rect 19154 39200 19210 40000
rect 19522 39200 19578 40000
rect 19890 39200 19946 40000
rect 20350 39200 20406 40000
rect 20718 39200 20774 40000
rect 21178 39200 21234 40000
rect 21546 39200 21602 40000
rect 21914 39200 21970 40000
rect 22374 39200 22430 40000
rect 22742 39200 22798 40000
rect 23202 39200 23258 40000
rect 23570 39200 23626 40000
rect 23938 39200 23994 40000
rect 24398 39200 24454 40000
rect 24766 39200 24822 40000
rect 25134 39200 25190 40000
rect 25594 39200 25650 40000
rect 25962 39200 26018 40000
rect 26422 39200 26478 40000
rect 26790 39200 26846 40000
rect 27158 39200 27214 40000
rect 27618 39200 27674 40000
rect 27986 39200 28042 40000
rect 28446 39200 28502 40000
rect 28814 39200 28870 40000
rect 29182 39200 29238 40000
rect 29642 39200 29698 40000
rect 30010 39200 30066 40000
rect 30116 39222 30328 39250
rect 15120 37074 15148 39200
rect 15384 37256 15436 37262
rect 15384 37198 15436 37204
rect 15200 37120 15252 37126
rect 15120 37068 15200 37074
rect 15120 37062 15252 37068
rect 15120 37046 15240 37062
rect 14464 36780 14516 36786
rect 15028 36774 15240 36802
rect 14464 36722 14516 36728
rect 14280 36372 14332 36378
rect 14280 36314 14332 36320
rect 14372 36168 14424 36174
rect 14372 36110 14424 36116
rect 14384 36009 14412 36110
rect 14370 36000 14426 36009
rect 14370 35935 14426 35944
rect 14476 35494 14504 36722
rect 15212 36718 15240 36774
rect 15200 36712 15252 36718
rect 15200 36654 15252 36660
rect 14464 35488 14516 35494
rect 14464 35430 14516 35436
rect 13726 34640 13782 34649
rect 13726 34575 13782 34584
rect 14476 34542 14504 35430
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 15016 34536 15068 34542
rect 15016 34478 15068 34484
rect 15028 31754 15056 34478
rect 15028 31726 15148 31754
rect 13358 30424 13414 30433
rect 13358 30359 13414 30368
rect 13360 26512 13412 26518
rect 13360 26454 13412 26460
rect 13372 23526 13400 26454
rect 13726 26344 13782 26353
rect 13726 26279 13782 26288
rect 13636 24336 13688 24342
rect 13634 24304 13636 24313
rect 13688 24304 13690 24313
rect 13634 24239 13690 24248
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13542 23624 13598 23633
rect 13542 23559 13598 23568
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13464 22817 13492 22918
rect 13450 22808 13506 22817
rect 13450 22743 13506 22752
rect 13464 22166 13492 22743
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 13450 21720 13506 21729
rect 13360 21684 13412 21690
rect 13450 21655 13506 21664
rect 13360 21626 13412 21632
rect 13372 21146 13400 21626
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13372 20806 13400 20946
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13358 19408 13414 19417
rect 13358 19343 13414 19352
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13188 18057 13216 18566
rect 13174 18048 13230 18057
rect 13174 17983 13230 17992
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13188 17270 13216 17818
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 13174 16688 13230 16697
rect 13174 16623 13176 16632
rect 13228 16623 13230 16632
rect 13176 16594 13228 16600
rect 13176 16448 13228 16454
rect 13174 16416 13176 16425
rect 13228 16416 13230 16425
rect 13174 16351 13230 16360
rect 13084 16176 13136 16182
rect 13084 16118 13136 16124
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 13004 15026 13032 16050
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12728 14912 12940 14940
rect 12624 14544 12676 14550
rect 12622 14512 12624 14521
rect 12716 14544 12768 14550
rect 12676 14512 12678 14521
rect 12716 14486 12768 14492
rect 12622 14447 12678 14456
rect 12728 14362 12756 14486
rect 12176 13790 12388 13818
rect 12636 14334 12756 14362
rect 12176 12594 12204 13790
rect 12254 13560 12310 13569
rect 12254 13495 12310 13504
rect 12268 13462 12296 13495
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12360 13161 12388 13330
rect 12346 13152 12402 13161
rect 12346 13087 12402 13096
rect 12176 12566 12388 12594
rect 12360 12458 12388 12566
rect 12360 12430 12480 12458
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12176 8634 12204 11698
rect 12452 10810 12480 12430
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11888 7404 11940 7410
rect 11992 7398 12112 7426
rect 11888 7346 11940 7352
rect 11900 7041 11928 7346
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11886 6760 11942 6769
rect 11886 6695 11942 6704
rect 11900 6458 11928 6695
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11794 5672 11850 5681
rect 11794 5607 11850 5616
rect 11808 5574 11836 5607
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11808 5370 11836 5510
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11348 2746 11468 2774
rect 11440 2514 11468 2746
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11612 1828 11664 1834
rect 11612 1770 11664 1776
rect 11244 1148 11296 1154
rect 11244 1090 11296 1096
rect 11440 870 11560 898
rect 11440 800 11468 870
rect 10612 734 10732 762
rect 10704 66 10732 734
rect 10692 60 10744 66
rect 10692 2 10744 8
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11532 626 11560 870
rect 11624 785 11652 1770
rect 11716 800 11744 3402
rect 11794 3360 11850 3369
rect 11794 3295 11850 3304
rect 11808 1426 11836 3295
rect 11900 3194 11928 5510
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11900 2514 11928 2790
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 11992 1766 12020 7278
rect 12084 6866 12112 7398
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 12084 5846 12112 6666
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 12176 5273 12204 8434
rect 12268 7342 12296 10746
rect 12438 10568 12494 10577
rect 12438 10503 12494 10512
rect 12452 10169 12480 10503
rect 12438 10160 12494 10169
rect 12438 10095 12494 10104
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12360 9602 12388 9998
rect 12360 9574 12480 9602
rect 12348 8424 12400 8430
rect 12346 8392 12348 8401
rect 12400 8392 12402 8401
rect 12346 8327 12402 8336
rect 12346 7984 12402 7993
rect 12346 7919 12402 7928
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12268 6066 12296 7142
rect 12360 6712 12388 7919
rect 12452 7002 12480 9574
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12440 6724 12492 6730
rect 12360 6684 12440 6712
rect 12360 6390 12388 6684
rect 12440 6666 12492 6672
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12268 6038 12388 6066
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12268 5817 12296 5850
rect 12254 5808 12310 5817
rect 12254 5743 12310 5752
rect 12360 5710 12388 6038
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12256 5296 12308 5302
rect 12162 5264 12218 5273
rect 12256 5238 12308 5244
rect 12162 5199 12218 5208
rect 12162 4856 12218 4865
rect 12162 4791 12218 4800
rect 12176 4010 12204 4791
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 12268 3194 12296 5238
rect 12438 4312 12494 4321
rect 12438 4247 12494 4256
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11796 1420 11848 1426
rect 11796 1362 11848 1368
rect 12084 800 12112 2246
rect 11610 776 11666 785
rect 11610 711 11666 720
rect 11532 598 11652 626
rect 11624 202 11652 598
rect 11612 196 11664 202
rect 11612 138 11664 144
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12268 202 12296 2994
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12360 800 12388 2926
rect 12452 2854 12480 4247
rect 12544 3618 12572 12378
rect 12636 11354 12664 14334
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12806 13696 12862 13705
rect 12728 13394 12756 13670
rect 12806 13631 12862 13640
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12728 12442 12756 13194
rect 12820 13161 12848 13631
rect 12806 13152 12862 13161
rect 12806 13087 12862 13096
rect 12912 13025 12940 14912
rect 13174 14648 13230 14657
rect 12992 14612 13044 14618
rect 13280 14618 13308 19110
rect 13372 18057 13400 19343
rect 13464 19281 13492 21655
rect 13556 20874 13584 23559
rect 13648 22642 13676 24142
rect 13740 22710 13768 26279
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 14108 24818 14136 25638
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 14188 24268 14240 24274
rect 14188 24210 14240 24216
rect 14096 24132 14148 24138
rect 14096 24074 14148 24080
rect 13912 23588 13964 23594
rect 13912 23530 13964 23536
rect 13728 22704 13780 22710
rect 13728 22646 13780 22652
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 13832 22094 13860 22646
rect 13924 22545 13952 23530
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 13910 22536 13966 22545
rect 13910 22471 13966 22480
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13740 22066 13860 22094
rect 13544 20868 13596 20874
rect 13544 20810 13596 20816
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13556 19961 13584 20334
rect 13542 19952 13598 19961
rect 13542 19887 13598 19896
rect 13544 19848 13596 19854
rect 13542 19816 13544 19825
rect 13596 19816 13598 19825
rect 13542 19751 13598 19760
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13556 19446 13584 19654
rect 13544 19440 13596 19446
rect 13648 19417 13676 20334
rect 13544 19382 13596 19388
rect 13634 19408 13690 19417
rect 13634 19343 13690 19352
rect 13544 19304 13596 19310
rect 13450 19272 13506 19281
rect 13544 19246 13596 19252
rect 13450 19207 13506 19216
rect 13556 19174 13584 19246
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13556 18698 13584 18838
rect 13544 18692 13596 18698
rect 13544 18634 13596 18640
rect 13358 18048 13414 18057
rect 13358 17983 13414 17992
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13372 17610 13400 17818
rect 13648 17746 13676 19178
rect 13740 18970 13768 22066
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13832 18034 13860 20402
rect 13740 18006 13860 18034
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13648 15706 13676 16730
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13740 15570 13768 18006
rect 13924 17678 13952 22374
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16454 13860 17070
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13450 15328 13506 15337
rect 13450 15263 13506 15272
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13174 14583 13176 14592
rect 12992 14554 13044 14560
rect 13228 14583 13230 14592
rect 13268 14612 13320 14618
rect 13176 14554 13228 14560
rect 13268 14554 13320 14560
rect 13004 13705 13032 14554
rect 13082 14512 13138 14521
rect 13082 14447 13138 14456
rect 12990 13696 13046 13705
rect 12990 13631 13046 13640
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12898 13016 12954 13025
rect 12820 12974 12898 13002
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12728 10470 12756 12242
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12622 9208 12678 9217
rect 12622 9143 12678 9152
rect 12636 9042 12664 9143
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12636 4826 12664 8978
rect 12728 8634 12756 10134
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12728 8362 12756 8570
rect 12820 8566 12848 12974
rect 12898 12951 12954 12960
rect 13004 12594 13032 13126
rect 12912 12566 13032 12594
rect 12912 11898 12940 12566
rect 12990 12472 13046 12481
rect 12990 12407 13046 12416
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 13004 11354 13032 12407
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12898 11248 12954 11257
rect 12898 11183 12900 11192
rect 12952 11183 12954 11192
rect 12900 11154 12952 11160
rect 13004 11098 13032 11290
rect 12912 11070 13032 11098
rect 12912 9353 12940 11070
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 13004 10198 13032 10950
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 12990 10024 13046 10033
rect 12990 9959 13046 9968
rect 13004 9926 13032 9959
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12898 9344 12954 9353
rect 12898 9279 12954 9288
rect 13004 9058 13032 9454
rect 13096 9178 13124 14447
rect 13372 14346 13400 15098
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13174 14240 13230 14249
rect 13174 14175 13230 14184
rect 13188 11082 13216 14175
rect 13372 13841 13400 14282
rect 13358 13832 13414 13841
rect 13358 13767 13414 13776
rect 13464 13190 13492 15263
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13556 13841 13584 14282
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13542 13832 13598 13841
rect 13542 13767 13598 13776
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13358 11928 13414 11937
rect 13358 11863 13360 11872
rect 13412 11863 13414 11872
rect 13360 11834 13412 11840
rect 13556 11744 13584 13670
rect 13372 11716 13584 11744
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13174 10976 13230 10985
rect 13174 10911 13230 10920
rect 13188 10169 13216 10911
rect 13280 10538 13308 11630
rect 13372 11150 13400 11716
rect 13648 11642 13676 14214
rect 13464 11626 13676 11642
rect 13452 11620 13676 11626
rect 13504 11614 13676 11620
rect 13452 11562 13504 11568
rect 13464 11370 13492 11562
rect 13464 11342 13584 11370
rect 13556 11150 13584 11342
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13174 10160 13230 10169
rect 13174 10095 13230 10104
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13188 9058 13216 10095
rect 13372 9568 13400 11086
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13464 10606 13492 10746
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13452 10600 13504 10606
rect 13556 10577 13584 10678
rect 13452 10542 13504 10548
rect 13542 10568 13598 10577
rect 13542 10503 13598 10512
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13004 9030 13216 9058
rect 13280 9540 13400 9568
rect 13004 8838 13032 9030
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12728 7478 12756 8298
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12728 5234 12756 7278
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12728 4554 12756 5170
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12820 4146 12848 8502
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 8090 13032 8230
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13280 8022 13308 9540
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 8974 13400 9386
rect 13556 9110 13584 10066
rect 13648 10044 13676 11222
rect 13740 10146 13768 15506
rect 13832 15502 13860 16390
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13910 14512 13966 14521
rect 13910 14447 13966 14456
rect 13924 14414 13952 14447
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 10248 13860 13806
rect 13924 11286 13952 14350
rect 14016 14346 14044 23462
rect 14108 23118 14136 24074
rect 14200 24070 14228 24210
rect 14188 24064 14240 24070
rect 14188 24006 14240 24012
rect 14278 23896 14334 23905
rect 14278 23831 14280 23840
rect 14332 23831 14334 23840
rect 14280 23802 14332 23808
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 14188 22976 14240 22982
rect 14188 22918 14240 22924
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 21593 14136 21966
rect 14094 21584 14150 21593
rect 14094 21519 14150 21528
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14108 19417 14136 19790
rect 14094 19408 14150 19417
rect 14094 19343 14150 19352
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14108 18873 14136 18906
rect 14094 18864 14150 18873
rect 14094 18799 14150 18808
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14108 17746 14136 18226
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 14108 17202 14136 17682
rect 14200 17270 14228 22918
rect 14292 22094 14320 23802
rect 14384 23526 14412 24550
rect 14372 23520 14424 23526
rect 14372 23462 14424 23468
rect 14384 23254 14412 23462
rect 14372 23248 14424 23254
rect 14372 23190 14424 23196
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14384 22710 14412 23054
rect 14372 22704 14424 22710
rect 14372 22646 14424 22652
rect 14292 22066 14412 22094
rect 14280 21548 14332 21554
rect 14280 21490 14332 21496
rect 14292 19145 14320 21490
rect 14384 21486 14412 22066
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14384 21185 14412 21286
rect 14370 21176 14426 21185
rect 14370 21111 14372 21120
rect 14424 21111 14426 21120
rect 14372 21082 14424 21088
rect 14384 21051 14412 21082
rect 14370 20632 14426 20641
rect 14370 20567 14426 20576
rect 14384 19922 14412 20567
rect 14372 19916 14424 19922
rect 14372 19858 14424 19864
rect 14278 19136 14334 19145
rect 14278 19071 14334 19080
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14292 17377 14320 18770
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14384 18426 14412 18702
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14476 17882 14504 25230
rect 14922 24984 14978 24993
rect 14922 24919 14978 24928
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 14740 23044 14792 23050
rect 14740 22986 14792 22992
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14660 22234 14688 22578
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14554 21992 14610 22001
rect 14554 21927 14610 21936
rect 14568 21622 14596 21927
rect 14556 21616 14608 21622
rect 14556 21558 14608 21564
rect 14646 21584 14702 21593
rect 14646 21519 14702 21528
rect 14660 21010 14688 21519
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14554 17504 14610 17513
rect 14554 17439 14610 17448
rect 14278 17368 14334 17377
rect 14278 17303 14334 17312
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14108 16182 14136 17138
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14384 16425 14412 16730
rect 14370 16416 14426 16425
rect 14370 16351 14426 16360
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14186 15736 14242 15745
rect 14186 15671 14242 15680
rect 14462 15736 14518 15745
rect 14462 15671 14464 15680
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14414 14136 14758
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14108 14006 14136 14350
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14016 13530 14044 13806
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14108 12850 14136 13262
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14094 12608 14150 12617
rect 14094 12543 14150 12552
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 13912 11280 13964 11286
rect 14016 11257 14044 11494
rect 13912 11222 13964 11228
rect 14002 11248 14058 11257
rect 14002 11183 14058 11192
rect 14016 11082 14044 11183
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 14002 10568 14058 10577
rect 14002 10503 14004 10512
rect 14056 10503 14058 10512
rect 14004 10474 14056 10480
rect 13832 10220 14044 10248
rect 13740 10118 13860 10146
rect 13648 10016 13768 10044
rect 13634 9888 13690 9897
rect 13634 9823 13690 9832
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8378 13400 8774
rect 13464 8566 13492 8978
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13372 8350 13492 8378
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13188 7857 13216 7890
rect 13174 7848 13230 7857
rect 13174 7783 13230 7792
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12912 6322 12940 6802
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12544 3590 12756 3618
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12452 1601 12480 2382
rect 12438 1592 12494 1601
rect 12438 1527 12494 1536
rect 12636 800 12664 3402
rect 12728 2922 12756 3590
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 13004 2446 13032 7142
rect 13096 6905 13124 7686
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 13082 6896 13138 6905
rect 13082 6831 13138 6840
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 6322 13124 6734
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13188 5778 13216 7414
rect 13280 7002 13308 7958
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13372 7478 13400 7890
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13280 5658 13308 6734
rect 13096 5630 13308 5658
rect 13096 5030 13124 5630
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13096 3126 13124 4966
rect 13188 4486 13216 5510
rect 13464 4758 13492 8350
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13556 6644 13584 8230
rect 13648 7410 13676 9823
rect 13740 8673 13768 10016
rect 13726 8664 13782 8673
rect 13726 8599 13782 8608
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13740 6866 13768 8599
rect 13832 7886 13860 10118
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13636 6656 13688 6662
rect 13556 6616 13636 6644
rect 13636 6598 13688 6604
rect 13542 6080 13598 6089
rect 13542 6015 13598 6024
rect 13556 5914 13584 6015
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13372 3738 13400 4150
rect 13556 4010 13584 4694
rect 13648 4690 13676 6598
rect 13726 6488 13782 6497
rect 13832 6474 13860 7278
rect 13782 6446 13860 6474
rect 13726 6423 13782 6432
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5846 13860 6054
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13726 5264 13782 5273
rect 13726 5199 13782 5208
rect 13740 5030 13768 5199
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13004 800 13032 2246
rect 13280 898 13308 2994
rect 13280 870 13400 898
rect 13280 800 13308 870
rect 12256 196 12308 202
rect 12256 138 12308 144
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13266 0 13322 800
rect 13372 338 13400 870
rect 13648 800 13676 3470
rect 13740 2961 13768 4966
rect 13818 4448 13874 4457
rect 13818 4383 13874 4392
rect 13832 3942 13860 4383
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13924 3738 13952 9522
rect 14016 9110 14044 10220
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 14016 8401 14044 9046
rect 14108 8673 14136 12543
rect 14200 9178 14228 15671
rect 14516 15671 14518 15680
rect 14464 15642 14516 15648
rect 14568 15144 14596 17439
rect 14476 15116 14596 15144
rect 14370 14104 14426 14113
rect 14370 14039 14426 14048
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14292 11529 14320 13126
rect 14278 11520 14334 11529
rect 14278 11455 14334 11464
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14292 10538 14320 10610
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14278 10432 14334 10441
rect 14278 10367 14334 10376
rect 14292 10062 14320 10367
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14292 9058 14320 9862
rect 14384 9178 14412 14039
rect 14476 13938 14504 15116
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14476 10169 14504 13738
rect 14568 10810 14596 14962
rect 14660 13802 14688 20334
rect 14752 19446 14780 22986
rect 14844 22778 14872 23122
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14844 22273 14872 22714
rect 14830 22264 14886 22273
rect 14830 22199 14886 22208
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 14844 20466 14872 21966
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14752 17882 14780 18566
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14752 15502 14780 16526
rect 14844 16114 14872 19790
rect 14936 16590 14964 24919
rect 15014 20632 15070 20641
rect 15014 20567 15070 20576
rect 15028 20466 15056 20567
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 15120 19922 15148 31726
rect 15198 25392 15254 25401
rect 15198 25327 15254 25336
rect 15212 24410 15240 25327
rect 15290 24848 15346 24857
rect 15290 24783 15346 24792
rect 15304 24585 15332 24783
rect 15290 24576 15346 24585
rect 15290 24511 15346 24520
rect 15200 24404 15252 24410
rect 15200 24346 15252 24352
rect 15292 23860 15344 23866
rect 15292 23802 15344 23808
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 15212 21962 15240 22102
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 15304 20874 15332 23802
rect 15396 22098 15424 37198
rect 15488 36378 15516 39200
rect 15948 37262 15976 39200
rect 15936 37256 15988 37262
rect 15936 37198 15988 37204
rect 16120 37188 16172 37194
rect 16120 37130 16172 37136
rect 15660 36780 15712 36786
rect 15660 36722 15712 36728
rect 15476 36372 15528 36378
rect 15476 36314 15528 36320
rect 15476 36168 15528 36174
rect 15476 36110 15528 36116
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15488 21554 15516 36110
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 15198 20632 15254 20641
rect 15198 20567 15254 20576
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 15212 19378 15240 20567
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14844 13954 14872 15642
rect 15028 15094 15056 19314
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15120 15881 15148 19246
rect 15198 18864 15254 18873
rect 15198 18799 15254 18808
rect 15106 15872 15162 15881
rect 15106 15807 15162 15816
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 14752 13926 14872 13954
rect 14924 13932 14976 13938
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14646 13560 14702 13569
rect 14646 13495 14702 13504
rect 14660 12646 14688 13495
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14752 12322 14780 13926
rect 15028 13920 15056 15030
rect 15108 14816 15160 14822
rect 15212 14804 15240 18799
rect 15304 18222 15332 19246
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15304 16998 15332 17070
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15160 14776 15240 14804
rect 15108 14758 15160 14764
rect 14976 13892 15056 13920
rect 14924 13874 14976 13880
rect 15120 13818 15148 14758
rect 15304 13841 15332 15098
rect 14936 13790 15148 13818
rect 15290 13832 15346 13841
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14844 12850 14872 13262
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14660 12294 14780 12322
rect 14660 11354 14688 12294
rect 14844 12238 14872 12786
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14740 11688 14792 11694
rect 14844 11676 14872 12174
rect 14792 11648 14872 11676
rect 14740 11630 14792 11636
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14830 11248 14886 11257
rect 14752 11150 14780 11222
rect 14830 11183 14886 11192
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14554 10568 14610 10577
rect 14554 10503 14610 10512
rect 14568 10266 14596 10503
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14462 10160 14518 10169
rect 14462 10095 14518 10104
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14462 9888 14518 9897
rect 14462 9823 14518 9832
rect 14476 9450 14504 9823
rect 14568 9722 14596 9998
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14660 9602 14688 11018
rect 14568 9574 14688 9602
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14200 9030 14320 9058
rect 14094 8664 14150 8673
rect 14094 8599 14150 8608
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14002 8392 14058 8401
rect 14002 8327 14058 8336
rect 14108 8265 14136 8502
rect 14094 8256 14150 8265
rect 14094 8191 14150 8200
rect 14096 7812 14148 7818
rect 14096 7754 14148 7760
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13820 2984 13872 2990
rect 13726 2952 13782 2961
rect 13820 2926 13872 2932
rect 13726 2887 13782 2896
rect 13832 1834 13860 2926
rect 14016 2446 14044 7686
rect 14108 7177 14136 7754
rect 14094 7168 14150 7177
rect 14094 7103 14150 7112
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 3942 14136 6598
rect 14200 6390 14228 9030
rect 14568 8922 14596 9574
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14292 8894 14596 8922
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14186 6216 14242 6225
rect 14186 6151 14188 6160
rect 14240 6151 14242 6160
rect 14188 6122 14240 6128
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 4622 14228 5102
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14188 4480 14240 4486
rect 14186 4448 14188 4457
rect 14240 4448 14242 4457
rect 14186 4383 14242 4392
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 14200 4049 14228 4150
rect 14292 4146 14320 8894
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14370 8392 14426 8401
rect 14370 8327 14426 8336
rect 14384 6662 14412 8327
rect 14462 7576 14518 7585
rect 14462 7511 14464 7520
rect 14516 7511 14518 7520
rect 14464 7482 14516 7488
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14476 6458 14504 7142
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14370 5672 14426 5681
rect 14370 5607 14372 5616
rect 14424 5607 14426 5616
rect 14372 5578 14424 5584
rect 14464 5568 14516 5574
rect 14384 5516 14464 5522
rect 14384 5510 14516 5516
rect 14384 5494 14504 5510
rect 14384 5166 14412 5494
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14186 4040 14242 4049
rect 14186 3975 14242 3984
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14384 3534 14412 3946
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14370 3224 14426 3233
rect 14568 3194 14596 8774
rect 14660 7478 14688 9386
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14660 6934 14688 7414
rect 14648 6928 14700 6934
rect 14648 6870 14700 6876
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14660 6186 14688 6258
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14660 3738 14688 5170
rect 14752 4826 14780 11086
rect 14844 10674 14872 11183
rect 14936 10810 14964 13790
rect 15290 13767 15346 13776
rect 15198 13288 15254 13297
rect 15108 13252 15160 13258
rect 15198 13223 15200 13232
rect 15108 13194 15160 13200
rect 15252 13223 15254 13232
rect 15200 13194 15252 13200
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 15028 12481 15056 12650
rect 15014 12472 15070 12481
rect 15120 12442 15148 13194
rect 15304 12968 15332 13767
rect 15212 12940 15332 12968
rect 15014 12407 15070 12416
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15108 12300 15160 12306
rect 15028 12260 15108 12288
rect 15028 11830 15056 12260
rect 15108 12242 15160 12248
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 15120 11098 15148 12038
rect 15212 11218 15240 12940
rect 15290 12880 15346 12889
rect 15290 12815 15292 12824
rect 15344 12815 15346 12824
rect 15292 12786 15344 12792
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15304 12102 15332 12378
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15304 11694 15332 11834
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15304 11354 15332 11630
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15120 11070 15332 11098
rect 15016 11008 15068 11014
rect 15014 10976 15016 10985
rect 15200 11008 15252 11014
rect 15068 10976 15070 10985
rect 15200 10950 15252 10956
rect 15014 10911 15070 10920
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14832 10532 14884 10538
rect 15028 10520 15056 10911
rect 15106 10840 15162 10849
rect 15106 10775 15162 10784
rect 14832 10474 14884 10480
rect 14936 10492 15056 10520
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14752 3670 14780 4626
rect 14844 3670 14872 10474
rect 14936 9926 14964 10492
rect 15014 10432 15070 10441
rect 15014 10367 15070 10376
rect 15028 10062 15056 10367
rect 15120 10266 15148 10775
rect 15212 10470 15240 10950
rect 15304 10810 15332 11070
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15290 10704 15346 10713
rect 15290 10639 15346 10648
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15304 10198 15332 10639
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 14922 9480 14978 9489
rect 14922 9415 14924 9424
rect 14976 9415 14978 9424
rect 14924 9386 14976 9392
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 14936 8974 14964 9046
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14936 8566 14964 8774
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 15028 8378 15056 9522
rect 15212 9518 15240 9862
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15120 8430 15148 9318
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 14936 8350 15056 8378
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 14936 5166 14964 8350
rect 15014 8256 15070 8265
rect 15014 8191 15070 8200
rect 15028 7886 15056 8191
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15014 7304 15070 7313
rect 15014 7239 15070 7248
rect 15028 5914 15056 7239
rect 15120 6798 15148 7822
rect 15212 7002 15240 8842
rect 15304 8401 15332 9522
rect 15290 8392 15346 8401
rect 15396 8362 15424 21422
rect 15476 20868 15528 20874
rect 15476 20810 15528 20816
rect 15488 16522 15516 20810
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 15474 16280 15530 16289
rect 15474 16215 15530 16224
rect 15488 16046 15516 16215
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15476 15428 15528 15434
rect 15580 15416 15608 22374
rect 15672 21078 15700 36722
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15764 24857 15792 24890
rect 15750 24848 15806 24857
rect 15750 24783 15806 24792
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15752 24064 15804 24070
rect 15752 24006 15804 24012
rect 15764 23866 15792 24006
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15856 22930 15884 24754
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15948 23118 15976 24550
rect 16132 23322 16160 37130
rect 16316 37126 16344 39200
rect 16684 37346 16712 39200
rect 16684 37318 16804 37346
rect 16672 37256 16724 37262
rect 16672 37198 16724 37204
rect 16580 37188 16632 37194
rect 16580 37130 16632 37136
rect 16304 37120 16356 37126
rect 16304 37062 16356 37068
rect 16304 26784 16356 26790
rect 16304 26726 16356 26732
rect 16316 24410 16344 26726
rect 16488 26580 16540 26586
rect 16488 26522 16540 26528
rect 16500 26314 16528 26522
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 16396 24744 16448 24750
rect 16396 24686 16448 24692
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16316 23798 16344 24346
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 16120 23316 16172 23322
rect 16120 23258 16172 23264
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15764 22902 15884 22930
rect 15764 22012 15792 22902
rect 15842 22808 15898 22817
rect 15842 22743 15844 22752
rect 15896 22743 15898 22752
rect 16028 22772 16080 22778
rect 15844 22714 15896 22720
rect 16028 22714 16080 22720
rect 16040 22438 16068 22714
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 15842 22264 15898 22273
rect 15842 22199 15898 22208
rect 15856 22094 15884 22199
rect 15856 22066 16068 22094
rect 15764 21984 15976 22012
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15660 21072 15712 21078
rect 15660 21014 15712 21020
rect 15658 19952 15714 19961
rect 15658 19887 15714 19896
rect 15672 19145 15700 19887
rect 15658 19136 15714 19145
rect 15658 19071 15714 19080
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15528 15388 15608 15416
rect 15476 15370 15528 15376
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15580 14414 15608 14894
rect 15672 14550 15700 17614
rect 15764 15434 15792 21830
rect 15842 21176 15898 21185
rect 15842 21111 15844 21120
rect 15896 21111 15898 21120
rect 15844 21082 15896 21088
rect 15948 21026 15976 21984
rect 15856 20998 15976 21026
rect 15856 17678 15884 20998
rect 16040 20534 16068 22066
rect 16028 20528 16080 20534
rect 16028 20470 16080 20476
rect 16132 20398 16160 23258
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16210 22808 16266 22817
rect 16210 22743 16266 22752
rect 16224 22409 16252 22743
rect 16210 22400 16266 22409
rect 16210 22335 16266 22344
rect 16316 22273 16344 22918
rect 16302 22264 16358 22273
rect 16302 22199 16358 22208
rect 16304 22092 16356 22098
rect 16304 22034 16356 22040
rect 16212 21412 16264 21418
rect 16212 21354 16264 21360
rect 16224 21010 16252 21354
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 16210 19952 16266 19961
rect 16210 19887 16212 19896
rect 16264 19887 16266 19896
rect 16212 19858 16264 19864
rect 16212 19780 16264 19786
rect 16212 19722 16264 19728
rect 16118 19680 16174 19689
rect 16118 19615 16174 19624
rect 16132 19378 16160 19615
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 15934 19272 15990 19281
rect 15934 19207 15990 19216
rect 15948 18834 15976 19207
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 16040 18426 16068 19314
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16026 18320 16082 18329
rect 16026 18255 16082 18264
rect 15844 17672 15896 17678
rect 16040 17649 16068 18255
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 15844 17614 15896 17620
rect 16026 17640 16082 17649
rect 16026 17575 16082 17584
rect 16026 16688 16082 16697
rect 16026 16623 16082 16632
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15856 16114 15884 16458
rect 15934 16144 15990 16153
rect 15844 16108 15896 16114
rect 15934 16079 15990 16088
rect 15844 16050 15896 16056
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15750 14104 15806 14113
rect 15750 14039 15806 14048
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15488 11830 15516 12786
rect 15672 12442 15700 13874
rect 15764 13870 15792 14039
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15856 13569 15884 14962
rect 15842 13560 15898 13569
rect 15842 13495 15898 13504
rect 15750 13288 15806 13297
rect 15750 13223 15806 13232
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15566 11792 15622 11801
rect 15290 8327 15346 8336
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15290 7712 15346 7721
rect 15290 7647 15346 7656
rect 15304 7206 15332 7647
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15396 7018 15424 7958
rect 15488 7886 15516 11766
rect 15566 11727 15568 11736
rect 15620 11727 15622 11736
rect 15672 11744 15700 12038
rect 15764 11898 15792 13223
rect 15948 13138 15976 16079
rect 15856 13110 15976 13138
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15752 11756 15804 11762
rect 15672 11716 15752 11744
rect 15568 11698 15620 11704
rect 15752 11698 15804 11704
rect 15750 11520 15806 11529
rect 15750 11455 15806 11464
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15580 10606 15608 11290
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15672 10996 15700 11086
rect 15764 11064 15792 11455
rect 15856 11218 15884 13110
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15948 11830 15976 12922
rect 15936 11824 15988 11830
rect 16040 11801 16068 16623
rect 16132 16454 16160 17682
rect 16224 17542 16252 19722
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16132 16289 16160 16390
rect 16118 16280 16174 16289
rect 16118 16215 16174 16224
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 15620 16160 16050
rect 16224 15745 16252 17478
rect 16316 16697 16344 22034
rect 16408 18970 16436 24686
rect 16500 23322 16528 26250
rect 16488 23316 16540 23322
rect 16488 23258 16540 23264
rect 16500 21010 16528 23258
rect 16592 21078 16620 37130
rect 16684 36922 16712 37198
rect 16672 36916 16724 36922
rect 16672 36858 16724 36864
rect 16776 36378 16804 37318
rect 17040 37256 17092 37262
rect 17040 37198 17092 37204
rect 17052 36553 17080 37198
rect 17144 36786 17172 39200
rect 17512 36802 17540 39200
rect 17776 37732 17828 37738
rect 17776 37674 17828 37680
rect 17132 36780 17184 36786
rect 17512 36774 17632 36802
rect 17132 36722 17184 36728
rect 17038 36544 17094 36553
rect 17038 36479 17094 36488
rect 16764 36372 16816 36378
rect 16764 36314 16816 36320
rect 16948 36168 17000 36174
rect 16948 36110 17000 36116
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16776 23866 16804 25094
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16868 23497 16896 24006
rect 16854 23488 16910 23497
rect 16854 23423 16910 23432
rect 16764 22092 16816 22098
rect 16764 22034 16816 22040
rect 16776 21876 16804 22034
rect 16856 22024 16908 22030
rect 16854 21992 16856 22001
rect 16908 21992 16910 22001
rect 16854 21927 16910 21936
rect 16776 21848 16896 21876
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 16592 20505 16620 20810
rect 16684 20777 16712 21422
rect 16776 21010 16804 21422
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16670 20768 16726 20777
rect 16670 20703 16726 20712
rect 16578 20496 16634 20505
rect 16578 20431 16634 20440
rect 16486 20360 16542 20369
rect 16486 20295 16542 20304
rect 16500 20262 16528 20295
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16670 20088 16726 20097
rect 16670 20023 16726 20032
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16500 19689 16528 19858
rect 16684 19718 16712 20023
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 16580 19712 16632 19718
rect 16486 19680 16542 19689
rect 16580 19654 16632 19660
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16486 19615 16542 19624
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16396 18964 16448 18970
rect 16396 18906 16448 18912
rect 16408 16998 16436 18906
rect 16500 18290 16528 19246
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16394 16824 16450 16833
rect 16394 16759 16450 16768
rect 16302 16688 16358 16697
rect 16408 16658 16436 16759
rect 16302 16623 16358 16632
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16500 16590 16528 18022
rect 16592 16640 16620 19654
rect 16672 18624 16724 18630
rect 16670 18592 16672 18601
rect 16724 18592 16726 18601
rect 16670 18527 16726 18536
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16684 18057 16712 18226
rect 16670 18048 16726 18057
rect 16670 17983 16726 17992
rect 16670 17232 16726 17241
rect 16776 17202 16804 19926
rect 16868 19786 16896 21848
rect 16960 21554 16988 36110
rect 17144 35834 17172 36722
rect 17500 36712 17552 36718
rect 17500 36654 17552 36660
rect 17132 35828 17184 35834
rect 17132 35770 17184 35776
rect 17408 27056 17460 27062
rect 17408 26998 17460 27004
rect 17316 24676 17368 24682
rect 17316 24618 17368 24624
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16670 17167 16672 17176
rect 16724 17167 16726 17176
rect 16764 17196 16816 17202
rect 16672 17138 16724 17144
rect 16764 17138 16816 17144
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16794 16712 16934
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16672 16652 16724 16658
rect 16592 16612 16672 16640
rect 16672 16594 16724 16600
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16670 16552 16726 16561
rect 16670 16487 16726 16496
rect 16394 16416 16450 16425
rect 16394 16351 16450 16360
rect 16210 15736 16266 15745
rect 16210 15671 16266 15680
rect 16132 15592 16252 15620
rect 16224 14929 16252 15592
rect 16210 14920 16266 14929
rect 16210 14855 16266 14864
rect 16118 14784 16174 14793
rect 16118 14719 16174 14728
rect 16132 12238 16160 14719
rect 16224 12986 16252 14855
rect 16304 14340 16356 14346
rect 16304 14282 16356 14288
rect 16316 13530 16344 14282
rect 16408 13841 16436 16351
rect 16684 16250 16712 16487
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16488 15904 16540 15910
rect 16486 15872 16488 15881
rect 16540 15872 16542 15881
rect 16486 15807 16542 15816
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16592 14958 16620 15302
rect 16684 15026 16712 15438
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 14278 16620 14758
rect 16684 14414 16712 14962
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16684 13938 16712 14350
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16394 13832 16450 13841
rect 16394 13767 16450 13776
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16210 12608 16266 12617
rect 16210 12543 16266 12552
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16120 12096 16172 12102
rect 16224 12084 16252 12543
rect 16316 12238 16344 13126
rect 16408 12730 16436 13767
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16408 12702 16528 12730
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16408 12442 16436 12582
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16500 12374 16528 12702
rect 16592 12646 16620 12922
rect 16684 12646 16712 13262
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16172 12056 16252 12084
rect 16120 12038 16172 12044
rect 15936 11766 15988 11772
rect 16026 11792 16082 11801
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15948 11098 15976 11766
rect 16026 11727 16082 11736
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16040 11218 16068 11630
rect 16132 11540 16160 12038
rect 16316 11898 16344 12174
rect 16684 12170 16712 12242
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16132 11512 16344 11540
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 16132 11150 16160 11290
rect 16120 11144 16172 11150
rect 15948 11070 16068 11098
rect 16120 11086 16172 11092
rect 15764 11036 15884 11064
rect 15672 10968 15792 10996
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 10130 15608 10406
rect 15672 10130 15700 10746
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15764 10010 15792 10968
rect 15580 9982 15792 10010
rect 15580 8498 15608 9982
rect 15856 9654 15884 11036
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15948 10033 15976 10406
rect 15934 10024 15990 10033
rect 15934 9959 15990 9968
rect 15844 9648 15896 9654
rect 15750 9616 15806 9625
rect 15844 9590 15896 9596
rect 15750 9551 15752 9560
rect 15804 9551 15806 9560
rect 15752 9522 15804 9528
rect 15658 9480 15714 9489
rect 15658 9415 15714 9424
rect 15752 9444 15804 9450
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15568 8288 15620 8294
rect 15566 8256 15568 8265
rect 15620 8256 15622 8265
rect 15566 8191 15622 8200
rect 15672 7886 15700 9415
rect 15752 9386 15804 9392
rect 15764 8906 15792 9386
rect 15752 8900 15804 8906
rect 15752 8842 15804 8848
rect 15764 8498 15792 8842
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15764 8022 15792 8434
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15568 7744 15620 7750
rect 15856 7698 15884 9590
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 15568 7686 15620 7692
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15304 6990 15424 7018
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15304 6610 15332 6990
rect 15382 6896 15438 6905
rect 15382 6831 15438 6840
rect 15212 6582 15332 6610
rect 15108 6384 15160 6390
rect 15106 6352 15108 6361
rect 15160 6352 15162 6361
rect 15106 6287 15162 6296
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 14936 4826 14964 5102
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 15028 3602 15056 5102
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15120 4162 15148 4966
rect 15212 4622 15240 6582
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15304 5778 15332 6394
rect 15396 6254 15424 6831
rect 15384 6248 15436 6254
rect 15382 6216 15384 6225
rect 15436 6216 15438 6225
rect 15382 6151 15438 6160
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15120 4134 15240 4162
rect 15212 3777 15240 4134
rect 15304 3942 15332 5714
rect 15384 4072 15436 4078
rect 15382 4040 15384 4049
rect 15436 4040 15438 4049
rect 15382 3975 15438 3984
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15198 3768 15254 3777
rect 15198 3703 15254 3712
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15106 3360 15162 3369
rect 15106 3295 15162 3304
rect 14370 3159 14372 3168
rect 14424 3159 14426 3168
rect 14556 3188 14608 3194
rect 14372 3130 14424 3136
rect 14556 3130 14608 3136
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 13912 2304 13964 2310
rect 13912 2246 13964 2252
rect 13820 1828 13872 1834
rect 13820 1770 13872 1776
rect 13924 800 13952 2246
rect 14292 898 14320 2994
rect 14660 2774 14688 2994
rect 14568 2746 14688 2774
rect 14292 870 14412 898
rect 14292 800 14320 870
rect 13360 332 13412 338
rect 13360 274 13412 280
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14384 134 14412 870
rect 14568 800 14596 2746
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14844 800 14872 2246
rect 15120 814 15148 3295
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15108 808 15160 814
rect 14372 128 14424 134
rect 14372 70 14424 76
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15212 800 15240 2246
rect 15396 1358 15424 3975
rect 15488 2378 15516 7686
rect 15580 2446 15608 7686
rect 15672 7670 15884 7698
rect 15672 6458 15700 7670
rect 15948 7562 15976 9046
rect 16040 8430 16068 11070
rect 16118 10024 16174 10033
rect 16118 9959 16174 9968
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16132 7857 16160 9959
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8566 16252 8774
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16316 7970 16344 11512
rect 16408 10985 16436 12038
rect 16500 11354 16528 12038
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16776 11257 16804 14350
rect 16762 11248 16818 11257
rect 16762 11183 16818 11192
rect 16670 11112 16726 11121
rect 16670 11047 16726 11056
rect 16684 11014 16712 11047
rect 16672 11008 16724 11014
rect 16394 10976 16450 10985
rect 16672 10950 16724 10956
rect 16394 10911 16450 10920
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16224 7942 16344 7970
rect 16118 7848 16174 7857
rect 16028 7812 16080 7818
rect 16118 7783 16174 7792
rect 16028 7754 16080 7760
rect 15856 7534 15976 7562
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15658 6352 15714 6361
rect 15658 6287 15714 6296
rect 15672 5710 15700 6287
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15672 5370 15700 5646
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15672 2258 15700 3470
rect 15764 2922 15792 7142
rect 15856 4146 15884 7534
rect 15936 7472 15988 7478
rect 15936 7414 15988 7420
rect 15948 6186 15976 7414
rect 16040 7342 16068 7754
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16040 6338 16068 7278
rect 16132 6458 16160 7783
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16040 6310 16160 6338
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15842 4040 15898 4049
rect 15842 3975 15898 3984
rect 15856 3641 15884 3975
rect 15842 3632 15898 3641
rect 15842 3567 15898 3576
rect 15948 3505 15976 5510
rect 15934 3496 15990 3505
rect 15934 3431 15990 3440
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 16040 2774 16068 5714
rect 16132 5370 16160 6310
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16224 4758 16252 7942
rect 16304 7880 16356 7886
rect 16302 7848 16304 7857
rect 16356 7848 16358 7857
rect 16302 7783 16358 7792
rect 16302 7168 16358 7177
rect 16302 7103 16358 7112
rect 16316 6866 16344 7103
rect 16408 6984 16436 9522
rect 16500 9450 16528 10474
rect 16592 9602 16620 10610
rect 16762 10568 16818 10577
rect 16762 10503 16818 10512
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 10305 16712 10406
rect 16670 10296 16726 10305
rect 16670 10231 16726 10240
rect 16776 10198 16804 10503
rect 16868 10305 16896 18158
rect 16960 18086 16988 21286
rect 17052 19666 17080 24550
rect 17224 24404 17276 24410
rect 17224 24346 17276 24352
rect 17236 24070 17264 24346
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17132 23860 17184 23866
rect 17132 23802 17184 23808
rect 17144 20874 17172 23802
rect 17236 22710 17264 24006
rect 17328 23050 17356 24618
rect 17420 24410 17448 26998
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 17408 23792 17460 23798
rect 17408 23734 17460 23740
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17224 22704 17276 22710
rect 17224 22646 17276 22652
rect 17132 20868 17184 20874
rect 17132 20810 17184 20816
rect 17236 20398 17264 22646
rect 17420 22098 17448 23734
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17408 21888 17460 21894
rect 17406 21856 17408 21865
rect 17460 21856 17462 21865
rect 17406 21791 17462 21800
rect 17316 21616 17368 21622
rect 17316 21558 17368 21564
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17144 19825 17172 20198
rect 17130 19816 17186 19825
rect 17130 19751 17186 19760
rect 17236 19689 17264 20198
rect 17222 19680 17278 19689
rect 17052 19638 17172 19666
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16960 17241 16988 17818
rect 16946 17232 17002 17241
rect 16946 17167 17002 17176
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 16960 12714 16988 16186
rect 17052 14090 17080 18838
rect 17144 18698 17172 19638
rect 17222 19615 17278 19624
rect 17222 19272 17278 19281
rect 17222 19207 17278 19216
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17130 18456 17186 18465
rect 17130 18391 17186 18400
rect 17144 18290 17172 18391
rect 17236 18329 17264 19207
rect 17328 18426 17356 21558
rect 17420 19990 17448 21791
rect 17512 21078 17540 36654
rect 17604 36378 17632 36774
rect 17788 36553 17816 37674
rect 17774 36544 17830 36553
rect 17774 36479 17830 36488
rect 17592 36372 17644 36378
rect 17880 36360 17908 39200
rect 18052 37868 18104 37874
rect 18052 37810 18104 37816
rect 17960 36372 18012 36378
rect 17880 36332 17960 36360
rect 17592 36314 17644 36320
rect 17960 36314 18012 36320
rect 17592 36168 17644 36174
rect 17592 36110 17644 36116
rect 17604 23322 17632 36110
rect 18064 31754 18092 37810
rect 18340 37330 18368 39200
rect 18328 37324 18380 37330
rect 18328 37266 18380 37272
rect 18604 37188 18656 37194
rect 18604 37130 18656 37136
rect 18236 36780 18288 36786
rect 18236 36722 18288 36728
rect 17972 31726 18092 31754
rect 17684 24880 17736 24886
rect 17684 24822 17736 24828
rect 17696 23662 17724 24822
rect 17776 24404 17828 24410
rect 17776 24346 17828 24352
rect 17684 23656 17736 23662
rect 17684 23598 17736 23604
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 17696 23202 17724 23598
rect 17788 23526 17816 24346
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17866 23488 17922 23497
rect 17866 23423 17922 23432
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 17604 23174 17724 23202
rect 17500 21072 17552 21078
rect 17500 21014 17552 21020
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17408 19984 17460 19990
rect 17408 19926 17460 19932
rect 17512 19786 17540 20334
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17512 19334 17540 19722
rect 17420 19306 17540 19334
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17222 18320 17278 18329
rect 17132 18284 17184 18290
rect 17420 18290 17448 19306
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17222 18255 17278 18264
rect 17408 18284 17460 18290
rect 17132 18226 17184 18232
rect 17236 18222 17264 18255
rect 17408 18226 17460 18232
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17130 17912 17186 17921
rect 17130 17847 17132 17856
rect 17184 17847 17186 17856
rect 17132 17818 17184 17824
rect 17236 17746 17264 18158
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17328 17678 17356 18158
rect 17512 18057 17540 18702
rect 17498 18048 17554 18057
rect 17498 17983 17554 17992
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17420 17678 17448 17818
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17408 17672 17460 17678
rect 17500 17672 17552 17678
rect 17408 17614 17460 17620
rect 17498 17640 17500 17649
rect 17552 17640 17554 17649
rect 17224 17604 17276 17610
rect 17498 17575 17554 17584
rect 17224 17546 17276 17552
rect 17236 17202 17264 17546
rect 17316 17536 17368 17542
rect 17500 17536 17552 17542
rect 17368 17496 17448 17524
rect 17316 17478 17368 17484
rect 17420 17377 17448 17496
rect 17500 17478 17552 17484
rect 17406 17368 17462 17377
rect 17512 17338 17540 17478
rect 17406 17303 17462 17312
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17604 16776 17632 23174
rect 17684 23044 17736 23050
rect 17684 22986 17736 22992
rect 17696 18766 17724 22986
rect 17788 22080 17816 23258
rect 17880 22642 17908 23423
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 17788 22052 17908 22080
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17788 18578 17816 21898
rect 17880 19990 17908 22052
rect 17972 21554 18000 31726
rect 18052 24880 18104 24886
rect 18052 24822 18104 24828
rect 18064 23905 18092 24822
rect 18050 23896 18106 23905
rect 18050 23831 18106 23840
rect 18052 23248 18104 23254
rect 18050 23216 18052 23225
rect 18104 23216 18106 23225
rect 18050 23151 18106 23160
rect 18248 22642 18276 36722
rect 18328 36168 18380 36174
rect 18328 36110 18380 36116
rect 18340 34649 18368 36110
rect 18420 35080 18472 35086
rect 18420 35022 18472 35028
rect 18326 34640 18382 34649
rect 18326 34575 18382 34584
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18156 22409 18184 22510
rect 18142 22400 18198 22409
rect 18142 22335 18198 22344
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17972 20330 18000 21490
rect 18052 21072 18104 21078
rect 18050 21040 18052 21049
rect 18104 21040 18106 21049
rect 18050 20975 18106 20984
rect 18156 20913 18184 21966
rect 18340 21962 18368 23462
rect 18432 22098 18460 35022
rect 18510 26072 18566 26081
rect 18510 26007 18566 26016
rect 18524 23497 18552 26007
rect 18510 23488 18566 23497
rect 18510 23423 18566 23432
rect 18616 23322 18644 37130
rect 18708 36922 18736 39200
rect 19064 37324 19116 37330
rect 19064 37266 19116 37272
rect 18696 36916 18748 36922
rect 18696 36858 18748 36864
rect 19076 35834 19104 37266
rect 19168 35894 19196 39200
rect 19536 37108 19564 39200
rect 19904 37210 19932 39200
rect 20260 37936 20312 37942
rect 20260 37878 20312 37884
rect 20076 37324 20128 37330
rect 20076 37266 20128 37272
rect 19904 37182 20024 37210
rect 19444 37080 19564 37108
rect 19444 36786 19472 37080
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 19340 36032 19392 36038
rect 19340 35974 19392 35980
rect 19352 35894 19380 35974
rect 19168 35866 19380 35894
rect 19444 35834 19472 36722
rect 19892 36712 19944 36718
rect 19892 36654 19944 36660
rect 19904 36145 19932 36654
rect 19996 36378 20024 37182
rect 19984 36372 20036 36378
rect 19984 36314 20036 36320
rect 19890 36136 19946 36145
rect 19890 36071 19946 36080
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 20088 35894 20116 37266
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19996 35866 20116 35894
rect 19064 35828 19116 35834
rect 19064 35770 19116 35776
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 19430 35320 19486 35329
rect 19430 35255 19486 35264
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 18880 25424 18932 25430
rect 18880 25366 18932 25372
rect 18892 25226 18920 25366
rect 18880 25220 18932 25226
rect 18880 25162 18932 25168
rect 18696 24948 18748 24954
rect 18696 24890 18748 24896
rect 18788 24948 18840 24954
rect 18788 24890 18840 24896
rect 18708 23866 18736 24890
rect 18800 24410 18828 24890
rect 19246 24848 19302 24857
rect 19246 24783 19302 24792
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 19156 24404 19208 24410
rect 19156 24346 19208 24352
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18694 23488 18750 23497
rect 18694 23423 18750 23432
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18510 23216 18566 23225
rect 18510 23151 18566 23160
rect 18524 22817 18552 23151
rect 18510 22808 18566 22817
rect 18510 22743 18566 22752
rect 18420 22092 18472 22098
rect 18420 22034 18472 22040
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18236 21344 18288 21350
rect 18340 21321 18368 21898
rect 18420 21344 18472 21350
rect 18236 21286 18288 21292
rect 18326 21312 18382 21321
rect 18142 20904 18198 20913
rect 18142 20839 18198 20848
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 18064 20210 18092 20538
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 17972 20182 18092 20210
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 17868 18828 17920 18834
rect 17868 18770 17920 18776
rect 17696 18550 17816 18578
rect 17696 16794 17724 18550
rect 17774 18456 17830 18465
rect 17774 18391 17830 18400
rect 17328 16748 17632 16776
rect 17684 16788 17736 16794
rect 17224 15632 17276 15638
rect 17224 15574 17276 15580
rect 17236 15366 17264 15574
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17052 14062 17172 14090
rect 17040 14000 17092 14006
rect 17040 13942 17092 13948
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16946 12200 17002 12209
rect 16946 12135 16948 12144
rect 17000 12135 17002 12144
rect 16948 12106 17000 12112
rect 17052 11914 17080 13942
rect 16960 11886 17080 11914
rect 16854 10296 16910 10305
rect 16854 10231 16910 10240
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16764 9988 16816 9994
rect 16764 9930 16816 9936
rect 16684 9761 16712 9930
rect 16776 9897 16804 9930
rect 16762 9888 16818 9897
rect 16762 9823 16818 9832
rect 16670 9752 16726 9761
rect 16960 9722 16988 11886
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17052 11393 17080 11698
rect 17038 11384 17094 11393
rect 17038 11319 17094 11328
rect 17144 11218 17172 14062
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17236 12753 17264 13126
rect 17222 12744 17278 12753
rect 17222 12679 17278 12688
rect 17328 12374 17356 16748
rect 17684 16730 17736 16736
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17408 15360 17460 15366
rect 17406 15328 17408 15337
rect 17460 15328 17462 15337
rect 17406 15263 17462 15272
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17420 13462 17448 14486
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17420 12850 17448 13126
rect 17498 12880 17554 12889
rect 17408 12844 17460 12850
rect 17498 12815 17500 12824
rect 17408 12786 17460 12792
rect 17552 12815 17554 12824
rect 17500 12786 17552 12792
rect 17604 12434 17632 16594
rect 17788 16182 17816 18391
rect 17880 18222 17908 18770
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17880 17746 17908 18158
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17972 17626 18000 20182
rect 18156 20058 18184 20402
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18248 19922 18276 21286
rect 18420 21286 18472 21292
rect 18326 21247 18382 21256
rect 18432 20856 18460 21286
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18340 20828 18460 20856
rect 18340 20534 18368 20828
rect 18418 20768 18474 20777
rect 18418 20703 18474 20712
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18432 20210 18460 20703
rect 18524 20534 18552 20946
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18708 20346 18736 23423
rect 18800 20482 18828 24142
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18892 21010 18920 23802
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 19076 22098 19104 23666
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 19168 20942 19196 24346
rect 19260 23186 19288 24783
rect 19352 24138 19380 26318
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19352 23633 19380 23666
rect 19338 23624 19394 23633
rect 19338 23559 19394 23568
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 19248 22976 19300 22982
rect 19246 22944 19248 22953
rect 19300 22944 19302 22953
rect 19246 22879 19302 22888
rect 19352 22545 19380 22986
rect 19338 22536 19394 22545
rect 19338 22471 19394 22480
rect 19444 22098 19472 35255
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19996 24410 20024 35866
rect 20168 35012 20220 35018
rect 20168 34954 20220 34960
rect 20076 32496 20128 32502
rect 20076 32438 20128 32444
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19890 22672 19946 22681
rect 19890 22607 19946 22616
rect 19904 22574 19932 22607
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19248 21956 19300 21962
rect 19248 21898 19300 21904
rect 19260 21865 19288 21898
rect 19246 21856 19302 21865
rect 19246 21791 19302 21800
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 19076 20754 19104 20810
rect 19076 20726 19196 20754
rect 18970 20632 19026 20641
rect 18970 20567 18972 20576
rect 19024 20567 19026 20576
rect 18972 20538 19024 20544
rect 18800 20454 19104 20482
rect 18708 20318 18828 20346
rect 18696 20256 18748 20262
rect 18432 20182 18552 20210
rect 18696 20198 18748 20204
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18142 19816 18198 19825
rect 18142 19751 18198 19760
rect 18156 19718 18184 19751
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18340 19378 18368 19654
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18142 19272 18198 19281
rect 18142 19207 18198 19216
rect 18236 19236 18288 19242
rect 18156 18902 18184 19207
rect 18236 19178 18288 19184
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 18064 18698 18092 18770
rect 18248 18748 18276 19178
rect 18156 18720 18276 18748
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 18064 18601 18092 18634
rect 18050 18592 18106 18601
rect 18050 18527 18106 18536
rect 18156 18442 18184 18720
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18064 18414 18184 18442
rect 18064 17785 18092 18414
rect 18156 18408 18184 18414
rect 18236 18420 18288 18426
rect 18156 18380 18236 18408
rect 18236 18362 18288 18368
rect 18144 18080 18196 18086
rect 18142 18048 18144 18057
rect 18340 18057 18368 18566
rect 18196 18048 18198 18057
rect 18142 17983 18198 17992
rect 18326 18048 18382 18057
rect 18326 17983 18382 17992
rect 18142 17912 18198 17921
rect 18432 17882 18460 19994
rect 18524 19378 18552 20182
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18524 18154 18552 18566
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18142 17847 18198 17856
rect 18420 17876 18472 17882
rect 18050 17776 18106 17785
rect 18050 17711 18106 17720
rect 17880 17598 18000 17626
rect 17880 17542 17908 17598
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 17880 16522 17908 17478
rect 17972 17270 18000 17478
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17776 16176 17828 16182
rect 17776 16118 17828 16124
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17682 15736 17738 15745
rect 17682 15671 17738 15680
rect 17420 12406 17632 12434
rect 17316 12368 17368 12374
rect 17314 12336 17316 12345
rect 17368 12336 17370 12345
rect 17314 12271 17370 12280
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17328 12102 17356 12174
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17420 11914 17448 12406
rect 17590 12336 17646 12345
rect 17590 12271 17646 12280
rect 17604 12238 17632 12271
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17512 12073 17540 12174
rect 17592 12096 17644 12102
rect 17498 12064 17554 12073
rect 17592 12038 17644 12044
rect 17498 11999 17554 12008
rect 17236 11886 17448 11914
rect 17500 11892 17552 11898
rect 17236 11234 17264 11886
rect 17500 11834 17552 11840
rect 17406 11792 17462 11801
rect 17406 11727 17462 11736
rect 17132 11212 17184 11218
rect 17236 11206 17356 11234
rect 17132 11154 17184 11160
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 16670 9687 16726 9696
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16946 9616 17002 9625
rect 16592 9574 16804 9602
rect 16580 9512 16632 9518
rect 16672 9512 16724 9518
rect 16632 9472 16672 9500
rect 16580 9454 16632 9460
rect 16672 9454 16724 9460
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16672 9376 16724 9382
rect 16776 9330 16804 9574
rect 16946 9551 17002 9560
rect 17052 9568 17080 11018
rect 17222 10840 17278 10849
rect 17222 10775 17278 10784
rect 17236 10606 17264 10775
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17222 10024 17278 10033
rect 17222 9959 17224 9968
rect 17276 9959 17278 9968
rect 17224 9930 17276 9936
rect 16960 9500 16988 9551
rect 17052 9540 17172 9568
rect 16724 9324 16804 9330
rect 16672 9318 16804 9324
rect 16684 9302 16804 9318
rect 16868 9472 16988 9500
rect 17038 9480 17094 9489
rect 16486 9208 16542 9217
rect 16762 9208 16818 9217
rect 16486 9143 16488 9152
rect 16540 9143 16542 9152
rect 16580 9172 16632 9178
rect 16488 9114 16540 9120
rect 16868 9178 16896 9472
rect 17038 9415 17040 9424
rect 17092 9415 17094 9424
rect 17040 9386 17092 9392
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16762 9143 16818 9152
rect 16856 9172 16908 9178
rect 16580 9114 16632 9120
rect 16592 9058 16620 9114
rect 16776 9110 16804 9143
rect 16856 9114 16908 9120
rect 16500 9030 16620 9058
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16500 7410 16528 9030
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16408 6956 16528 6984
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16394 6080 16450 6089
rect 16394 6015 16450 6024
rect 16408 5914 16436 6015
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16212 4752 16264 4758
rect 16212 4694 16264 4700
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 15948 2746 16068 2774
rect 15948 2446 15976 2746
rect 15936 2440 15988 2446
rect 15842 2408 15898 2417
rect 15936 2382 15988 2388
rect 15842 2343 15898 2352
rect 15856 2310 15884 2343
rect 15488 2230 15700 2258
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 15488 800 15516 2230
rect 15948 1170 15976 2246
rect 15856 1142 15976 1170
rect 15856 800 15884 1142
rect 16132 898 16160 2994
rect 16132 870 16252 898
rect 16316 882 16344 5170
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16408 3126 16436 4558
rect 16500 4298 16528 6956
rect 16592 5914 16620 8366
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16684 6746 16712 8230
rect 16776 6882 16804 8910
rect 16960 8616 16988 9318
rect 17038 9208 17094 9217
rect 17038 9143 17094 9152
rect 17052 8906 17080 9143
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 16868 8588 16988 8616
rect 16868 8294 16896 8588
rect 16946 8528 17002 8537
rect 16946 8463 17002 8472
rect 16960 8362 16988 8463
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16856 8288 16908 8294
rect 17144 8242 17172 9540
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17236 9178 17264 9454
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 16856 8230 16908 8236
rect 17052 8214 17172 8242
rect 16948 7880 17000 7886
rect 16946 7848 16948 7857
rect 17000 7848 17002 7857
rect 16946 7783 17002 7792
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16776 6854 16896 6882
rect 16684 6718 16804 6746
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16684 5302 16712 6598
rect 16776 5953 16804 6718
rect 16762 5944 16818 5953
rect 16762 5879 16818 5888
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 16684 4826 16712 5238
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16500 4270 16620 4298
rect 16592 4146 16620 4270
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16396 3120 16448 3126
rect 16396 3062 16448 3068
rect 16132 800 16160 870
rect 15108 750 15160 756
rect 15198 0 15254 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16224 270 16252 870
rect 16304 876 16356 882
rect 16304 818 16356 824
rect 16500 800 16528 3470
rect 16580 3392 16632 3398
rect 16578 3360 16580 3369
rect 16632 3360 16634 3369
rect 16578 3295 16634 3304
rect 16776 2938 16804 5646
rect 16868 5370 16896 6854
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16854 5128 16910 5137
rect 16854 5063 16910 5072
rect 16684 2910 16804 2938
rect 16684 2854 16712 2910
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16776 800 16804 2790
rect 16212 264 16264 270
rect 16212 206 16264 212
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 16868 746 16896 5063
rect 16960 5012 16988 7414
rect 17052 5710 17080 8214
rect 17130 6896 17186 6905
rect 17130 6831 17186 6840
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 17040 5024 17092 5030
rect 16960 4984 17040 5012
rect 17040 4966 17092 4972
rect 17052 3233 17080 4966
rect 17038 3224 17094 3233
rect 17038 3159 17094 3168
rect 17144 3058 17172 6831
rect 17236 6769 17264 8910
rect 17328 7313 17356 11206
rect 17420 8673 17448 11727
rect 17512 11694 17540 11834
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 8974 17540 11494
rect 17604 10266 17632 12038
rect 17696 10690 17724 15671
rect 17788 11626 17816 15846
rect 17972 15502 18000 16050
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17880 14249 17908 15302
rect 18064 15026 18092 17478
rect 18156 16658 18184 17847
rect 18420 17818 18472 17824
rect 18510 17776 18566 17785
rect 18510 17711 18566 17720
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18340 17066 18368 17614
rect 18524 17610 18552 17711
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18616 17490 18644 19790
rect 18708 17746 18736 20198
rect 18800 19242 18828 20318
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18892 18873 18920 19110
rect 18878 18864 18934 18873
rect 18878 18799 18934 18808
rect 18788 18692 18840 18698
rect 18788 18634 18840 18640
rect 18800 18290 18828 18634
rect 18878 18456 18934 18465
rect 18878 18391 18880 18400
rect 18932 18391 18934 18400
rect 18880 18362 18932 18368
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18800 17610 18828 18226
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18788 17604 18840 17610
rect 18524 17462 18644 17490
rect 18708 17564 18788 17592
rect 18524 17202 18552 17462
rect 18602 17368 18658 17377
rect 18602 17303 18604 17312
rect 18656 17303 18658 17312
rect 18604 17274 18656 17280
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 18512 16992 18564 16998
rect 18564 16969 18644 16980
rect 18564 16960 18658 16969
rect 18564 16952 18602 16960
rect 18512 16934 18564 16940
rect 18602 16895 18658 16904
rect 18418 16824 18474 16833
rect 18236 16788 18288 16794
rect 18418 16759 18474 16768
rect 18236 16730 18288 16736
rect 18144 16652 18196 16658
rect 18144 16594 18196 16600
rect 18248 16425 18276 16730
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18234 16416 18290 16425
rect 18234 16351 18290 16360
rect 18234 16280 18290 16289
rect 18234 16215 18290 16224
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 17866 14240 17922 14249
rect 18050 14240 18106 14249
rect 17866 14175 17922 14184
rect 17972 14198 18050 14226
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17880 12617 17908 13330
rect 17972 12968 18000 14198
rect 18050 14175 18106 14184
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18064 13938 18092 14010
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 18156 13734 18184 15642
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18142 13424 18198 13433
rect 18142 13359 18198 13368
rect 18156 13190 18184 13359
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 17972 12940 18184 12968
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17866 12608 17922 12617
rect 17866 12543 17922 12552
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17866 11384 17922 11393
rect 17972 11370 18000 12786
rect 18050 12472 18106 12481
rect 18050 12407 18106 12416
rect 18064 12374 18092 12407
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 17972 11342 18092 11370
rect 17866 11319 17868 11328
rect 17920 11319 17922 11328
rect 17868 11290 17920 11296
rect 18064 11234 18092 11342
rect 17880 11206 18092 11234
rect 17696 10662 17816 10690
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17696 10062 17724 10542
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17788 9722 17816 10662
rect 17880 10198 17908 11206
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17590 9480 17646 9489
rect 17590 9415 17592 9424
rect 17644 9415 17646 9424
rect 17592 9386 17644 9392
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17406 8664 17462 8673
rect 17406 8599 17462 8608
rect 17406 8120 17462 8129
rect 17406 8055 17408 8064
rect 17460 8055 17462 8064
rect 17408 8026 17460 8032
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17314 7304 17370 7313
rect 17314 7239 17370 7248
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17222 6760 17278 6769
rect 17222 6695 17278 6704
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17052 800 17080 2926
rect 17236 2446 17264 6598
rect 17328 4826 17356 6938
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17328 4457 17356 4762
rect 17314 4448 17370 4457
rect 17314 4383 17370 4392
rect 17314 4176 17370 4185
rect 17420 4146 17448 7754
rect 17314 4111 17370 4120
rect 17408 4140 17460 4146
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17328 2106 17356 4111
rect 17408 4082 17460 4088
rect 17512 2514 17540 8774
rect 17604 8362 17632 9114
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17604 7478 17632 8298
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17604 5817 17632 6054
rect 17590 5808 17646 5817
rect 17590 5743 17646 5752
rect 17592 5704 17644 5710
rect 17590 5672 17592 5681
rect 17644 5672 17646 5681
rect 17590 5607 17646 5616
rect 17696 4321 17724 9590
rect 17880 9586 17908 9998
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17972 9382 18000 10202
rect 18064 9738 18092 11018
rect 18156 10674 18184 12940
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 18142 10296 18198 10305
rect 18142 10231 18144 10240
rect 18196 10231 18198 10240
rect 18144 10202 18196 10208
rect 18064 9710 18184 9738
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17960 9376 18012 9382
rect 17866 9344 17922 9353
rect 17960 9318 18012 9324
rect 17866 9279 17922 9288
rect 17880 8634 17908 9279
rect 18064 9217 18092 9454
rect 18050 9208 18106 9217
rect 18050 9143 18106 9152
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17682 4312 17738 4321
rect 17682 4247 17738 4256
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17604 2854 17632 4014
rect 17788 3194 17816 8434
rect 17880 6458 17908 8570
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17972 7274 18000 8230
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17880 5370 17908 6190
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17972 5030 18000 6870
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17592 2848 17644 2854
rect 17592 2790 17644 2796
rect 17774 2680 17830 2689
rect 17774 2615 17830 2624
rect 17788 2582 17816 2615
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17316 2100 17368 2106
rect 17316 2042 17368 2048
rect 17314 1592 17370 1601
rect 17314 1527 17370 1536
rect 17328 1290 17356 1527
rect 17316 1284 17368 1290
rect 17316 1226 17368 1232
rect 17420 800 17448 2314
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17788 1170 17816 2246
rect 17880 1737 17908 3334
rect 17972 3194 18000 3402
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18064 2922 18092 8842
rect 18156 7954 18184 9710
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18144 7812 18196 7818
rect 18144 7754 18196 7760
rect 18156 5370 18184 7754
rect 18248 6730 18276 16215
rect 18340 15366 18368 16526
rect 18432 15910 18460 16759
rect 18708 16640 18736 17564
rect 18788 17546 18840 17552
rect 18786 17368 18842 17377
rect 18786 17303 18842 17312
rect 18800 17270 18828 17303
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18800 16794 18828 17070
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18708 16612 18828 16640
rect 18694 16552 18750 16561
rect 18694 16487 18750 16496
rect 18708 16454 18736 16487
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18616 16046 18644 16390
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18340 13870 18368 15302
rect 18432 14822 18460 15846
rect 18602 15192 18658 15201
rect 18602 15127 18604 15136
rect 18656 15127 18658 15136
rect 18696 15156 18748 15162
rect 18604 15098 18656 15104
rect 18696 15098 18748 15104
rect 18602 14920 18658 14929
rect 18602 14855 18658 14864
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18616 14532 18644 14855
rect 18708 14657 18736 15098
rect 18694 14648 18750 14657
rect 18694 14583 18750 14592
rect 18616 14504 18736 14532
rect 18708 14414 18736 14504
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 13988 18460 14214
rect 18512 14000 18564 14006
rect 18432 13960 18512 13988
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18432 13512 18460 13960
rect 18512 13942 18564 13948
rect 18604 13932 18656 13938
rect 18708 13920 18736 14350
rect 18656 13892 18736 13920
rect 18604 13874 18656 13880
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18616 13546 18644 13738
rect 18340 13484 18460 13512
rect 18524 13518 18644 13546
rect 18340 13326 18368 13484
rect 18524 13444 18552 13518
rect 18432 13416 18552 13444
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18340 12714 18368 12922
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18432 12617 18460 13416
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18602 13288 18658 13297
rect 18418 12608 18474 12617
rect 18418 12543 18474 12552
rect 18326 12472 18382 12481
rect 18326 12407 18382 12416
rect 18340 12238 18368 12407
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18340 11937 18368 12174
rect 18326 11928 18382 11937
rect 18326 11863 18382 11872
rect 18432 11676 18460 12543
rect 18524 11778 18552 13262
rect 18602 13223 18658 13232
rect 18616 12646 18644 13223
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18616 12073 18644 12582
rect 18708 12442 18736 12922
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18602 12064 18658 12073
rect 18602 11999 18658 12008
rect 18602 11928 18658 11937
rect 18602 11863 18604 11872
rect 18656 11863 18658 11872
rect 18604 11834 18656 11840
rect 18524 11750 18644 11778
rect 18432 11648 18552 11676
rect 18418 11248 18474 11257
rect 18418 11183 18474 11192
rect 18432 11150 18460 11183
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18328 11008 18380 11014
rect 18524 10996 18552 11648
rect 18328 10950 18380 10956
rect 18432 10968 18552 10996
rect 18340 9654 18368 10950
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18340 8945 18368 9454
rect 18326 8936 18382 8945
rect 18326 8871 18382 8880
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 18340 5914 18368 8871
rect 18432 8022 18460 10968
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18524 10266 18552 10474
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18512 9988 18564 9994
rect 18512 9930 18564 9936
rect 18524 9761 18552 9930
rect 18616 9908 18644 11750
rect 18800 11642 18828 16612
rect 18892 16289 18920 17682
rect 18984 17649 19012 19994
rect 18970 17640 19026 17649
rect 18970 17575 19026 17584
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 16998 19012 17478
rect 19076 17082 19104 20454
rect 19168 20058 19196 20726
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19260 19530 19288 21286
rect 19352 20874 19380 22034
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19892 21616 19944 21622
rect 19892 21558 19944 21564
rect 19798 21312 19854 21321
rect 19798 21247 19854 21256
rect 19812 21078 19840 21247
rect 19800 21072 19852 21078
rect 19800 21014 19852 21020
rect 19904 20942 19932 21558
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19996 20874 20024 24210
rect 20088 23866 20116 32438
rect 20076 23860 20128 23866
rect 20076 23802 20128 23808
rect 20088 22094 20116 23802
rect 20180 22642 20208 34954
rect 20272 24857 20300 37878
rect 20364 36922 20392 39200
rect 20732 37262 20760 39200
rect 20904 37936 20956 37942
rect 20904 37878 20956 37884
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 20352 36916 20404 36922
rect 20352 36858 20404 36864
rect 20628 36780 20680 36786
rect 20628 36722 20680 36728
rect 20536 36168 20588 36174
rect 20536 36110 20588 36116
rect 20444 36100 20496 36106
rect 20444 36042 20496 36048
rect 20350 28928 20406 28937
rect 20350 28863 20406 28872
rect 20258 24848 20314 24857
rect 20258 24783 20314 24792
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 20272 23526 20300 24074
rect 20260 23520 20312 23526
rect 20260 23462 20312 23468
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 20088 22066 20208 22094
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 19168 19502 19288 19530
rect 19168 19310 19196 19502
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19168 19174 19196 19246
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19154 19000 19210 19009
rect 19154 18935 19210 18944
rect 19168 18154 19196 18935
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19260 17882 19288 19382
rect 19156 17876 19208 17882
rect 19156 17818 19208 17824
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19168 17542 19196 17818
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19076 17054 19196 17082
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18878 16280 18934 16289
rect 18878 16215 18934 16224
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18892 16017 18920 16050
rect 18878 16008 18934 16017
rect 18878 15943 18934 15952
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18892 13802 18920 14962
rect 18984 14890 19012 16934
rect 19168 16833 19196 17054
rect 19154 16824 19210 16833
rect 19154 16759 19210 16768
rect 19156 16720 19208 16726
rect 19062 16688 19118 16697
rect 19156 16662 19208 16668
rect 19062 16623 19118 16632
rect 19076 16046 19104 16623
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 19076 15881 19104 15982
rect 19168 15978 19196 16662
rect 19260 16182 19288 17818
rect 19352 16998 19380 20810
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19522 20496 19578 20505
rect 19522 20431 19578 20440
rect 19536 20398 19564 20431
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19430 20088 19486 20097
rect 19430 20023 19486 20032
rect 19444 19514 19472 20023
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19996 19446 20024 20810
rect 20180 19854 20208 22066
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19444 17626 19472 19314
rect 19628 19310 19656 19382
rect 19892 19372 19944 19378
rect 20272 19334 20300 21966
rect 19892 19314 19944 19320
rect 19616 19304 19668 19310
rect 19522 19272 19578 19281
rect 19616 19246 19668 19252
rect 19522 19207 19524 19216
rect 19576 19207 19578 19216
rect 19800 19236 19852 19242
rect 19524 19178 19576 19184
rect 19800 19178 19852 19184
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19706 19136 19762 19145
rect 19524 18896 19576 18902
rect 19628 18884 19656 19110
rect 19706 19071 19762 19080
rect 19576 18856 19656 18884
rect 19524 18838 19576 18844
rect 19616 18760 19668 18766
rect 19720 18748 19748 19071
rect 19812 18902 19840 19178
rect 19800 18896 19852 18902
rect 19800 18838 19852 18844
rect 19668 18720 19748 18748
rect 19798 18728 19854 18737
rect 19616 18702 19668 18708
rect 19798 18663 19800 18672
rect 19852 18663 19854 18672
rect 19800 18634 19852 18640
rect 19904 18612 19932 19314
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 20180 19306 20300 19334
rect 19904 18584 19950 18612
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19922 18408 19950 18584
rect 19904 18380 19950 18408
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19536 18086 19564 18158
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19536 17954 19564 18022
rect 19536 17926 19656 17954
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19536 17746 19564 17818
rect 19524 17740 19576 17746
rect 19524 17682 19576 17688
rect 19628 17649 19656 17926
rect 19720 17785 19748 18158
rect 19800 17808 19852 17814
rect 19706 17776 19762 17785
rect 19800 17750 19852 17756
rect 19706 17711 19762 17720
rect 19812 17678 19840 17750
rect 19800 17672 19852 17678
rect 19614 17640 19670 17649
rect 19444 17598 19564 17626
rect 19536 17524 19564 17598
rect 19800 17614 19852 17620
rect 19614 17575 19670 17584
rect 19444 17496 19564 17524
rect 19904 17524 19932 18380
rect 19996 18154 20024 19246
rect 20076 18896 20128 18902
rect 20076 18838 20128 18844
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19982 17776 20038 17785
rect 19982 17711 20038 17720
rect 19996 17678 20024 17711
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19904 17496 19950 17524
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16794 19380 16934
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19062 15872 19118 15881
rect 19062 15807 19118 15816
rect 19352 15722 19380 16458
rect 19444 15978 19472 17496
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19922 17320 19950 17496
rect 19982 17504 20038 17513
rect 19982 17439 20038 17448
rect 19628 17292 19950 17320
rect 19628 17134 19656 17292
rect 19996 17270 20024 17439
rect 19984 17264 20036 17270
rect 19706 17232 19762 17241
rect 19984 17206 20036 17212
rect 19706 17167 19762 17176
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19628 16658 19656 17070
rect 19720 16794 19748 17167
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19812 16697 19840 17070
rect 19798 16688 19854 16697
rect 19616 16652 19668 16658
rect 19798 16623 19854 16632
rect 19616 16594 19668 16600
rect 19996 16590 20024 17206
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 20088 16425 20116 18838
rect 20180 18714 20208 19306
rect 20260 19236 20312 19242
rect 20260 19178 20312 19184
rect 20272 18970 20300 19178
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20364 18902 20392 28863
rect 20456 23186 20484 36042
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20548 22098 20576 36110
rect 20536 22092 20588 22098
rect 20536 22034 20588 22040
rect 20640 21554 20668 36722
rect 20732 36378 20760 37198
rect 20720 36372 20772 36378
rect 20720 36314 20772 36320
rect 20810 27432 20866 27441
rect 20810 27367 20866 27376
rect 20718 25936 20774 25945
rect 20718 25871 20774 25880
rect 20732 25265 20760 25871
rect 20718 25256 20774 25265
rect 20718 25191 20774 25200
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 21010 20484 21286
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20536 20800 20588 20806
rect 20442 20768 20498 20777
rect 20536 20742 20588 20748
rect 20442 20703 20498 20712
rect 20456 20602 20484 20703
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20456 20058 20484 20538
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20456 19446 20484 19994
rect 20548 19530 20576 20742
rect 20732 20097 20760 23462
rect 20824 20602 20852 27367
rect 20916 20806 20944 37878
rect 21086 37496 21142 37505
rect 21086 37431 21142 37440
rect 21100 37398 21128 37431
rect 21088 37392 21140 37398
rect 21088 37334 21140 37340
rect 21192 36922 21220 39200
rect 21456 37664 21508 37670
rect 21456 37606 21508 37612
rect 21180 36916 21232 36922
rect 21180 36858 21232 36864
rect 20996 34672 21048 34678
rect 20996 34614 21048 34620
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20718 20088 20774 20097
rect 20718 20023 20774 20032
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20640 19689 20668 19790
rect 20626 19680 20682 19689
rect 20626 19615 20682 19624
rect 20548 19502 20668 19530
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20534 19272 20590 19281
rect 20534 19207 20590 19216
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20352 18896 20404 18902
rect 20456 18873 20484 19110
rect 20352 18838 20404 18844
rect 20442 18864 20498 18873
rect 20442 18799 20498 18808
rect 20456 18766 20484 18799
rect 20444 18760 20496 18766
rect 20180 18686 20300 18714
rect 20444 18702 20496 18708
rect 20272 17954 20300 18686
rect 20350 18320 20406 18329
rect 20350 18255 20406 18264
rect 20180 17926 20300 17954
rect 20180 16946 20208 17926
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20272 17241 20300 17478
rect 20258 17232 20314 17241
rect 20258 17167 20314 17176
rect 20364 17134 20392 18255
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20456 18057 20484 18158
rect 20548 18154 20576 19207
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 20442 18048 20498 18057
rect 20442 17983 20498 17992
rect 20442 17912 20498 17921
rect 20442 17847 20444 17856
rect 20496 17847 20498 17856
rect 20444 17818 20496 17824
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20444 17264 20496 17270
rect 20444 17206 20496 17212
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20180 16918 20392 16946
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20180 16658 20208 16730
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20260 16584 20312 16590
rect 20180 16532 20260 16538
rect 20180 16526 20312 16532
rect 20180 16510 20300 16526
rect 20074 16416 20130 16425
rect 19574 16348 19882 16368
rect 20074 16351 20130 16360
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19982 16280 20038 16289
rect 19904 16224 19982 16232
rect 19904 16215 20038 16224
rect 19904 16204 20024 16215
rect 19904 16114 19932 16204
rect 20076 16176 20128 16182
rect 20076 16118 20128 16124
rect 19892 16108 19944 16114
rect 19720 16068 19892 16096
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19614 15872 19670 15881
rect 19614 15807 19670 15816
rect 19076 15694 19380 15722
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 19076 13818 19104 15694
rect 19248 15632 19300 15638
rect 19246 15600 19248 15609
rect 19300 15600 19302 15609
rect 19156 15564 19208 15570
rect 19628 15570 19656 15807
rect 19246 15535 19302 15544
rect 19616 15564 19668 15570
rect 19156 15506 19208 15512
rect 19616 15506 19668 15512
rect 19168 14657 19196 15506
rect 19524 15496 19576 15502
rect 19720 15450 19748 16068
rect 19892 16050 19944 16056
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19996 15881 20024 16050
rect 19982 15872 20038 15881
rect 19982 15807 20038 15816
rect 20088 15722 20116 16118
rect 19576 15444 19748 15450
rect 19524 15438 19748 15444
rect 19536 15422 19748 15438
rect 19996 15694 20116 15722
rect 19996 15434 20024 15694
rect 20074 15600 20130 15609
rect 20180 15570 20208 16510
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20074 15535 20130 15544
rect 20168 15564 20220 15570
rect 20088 15502 20116 15535
rect 20168 15506 20220 15512
rect 20076 15496 20128 15502
rect 20272 15473 20300 16390
rect 20076 15438 20128 15444
rect 20258 15464 20314 15473
rect 19984 15428 20036 15434
rect 20258 15399 20314 15408
rect 19984 15370 20036 15376
rect 19430 15328 19486 15337
rect 19430 15263 19486 15272
rect 19444 15144 19472 15263
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19996 15201 20024 15370
rect 20168 15360 20220 15366
rect 20166 15328 20168 15337
rect 20220 15328 20222 15337
rect 20166 15263 20222 15272
rect 19982 15192 20038 15201
rect 19444 15116 19564 15144
rect 20364 15144 20392 16918
rect 20456 15314 20484 17206
rect 20548 17134 20576 17478
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20640 16522 20668 19502
rect 20718 19136 20774 19145
rect 20718 19071 20774 19080
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20534 16416 20590 16425
rect 20534 16351 20590 16360
rect 20548 16114 20576 16351
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20534 16008 20590 16017
rect 20534 15943 20590 15952
rect 20548 15910 20576 15943
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20548 15706 20576 15846
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20534 15600 20590 15609
rect 20640 15586 20668 16458
rect 20732 15978 20760 19071
rect 20824 18766 20852 20538
rect 20916 20466 20944 20742
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20916 19174 20944 20198
rect 21008 19922 21036 34614
rect 21178 23488 21234 23497
rect 21178 23423 21234 23432
rect 21192 22710 21220 23423
rect 21364 23248 21416 23254
rect 21364 23190 21416 23196
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21180 22704 21232 22710
rect 21180 22646 21232 22652
rect 21284 22506 21312 23054
rect 21088 22500 21140 22506
rect 21088 22442 21140 22448
rect 21272 22500 21324 22506
rect 21272 22442 21324 22448
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 21100 19446 21128 22442
rect 21376 22409 21404 23190
rect 21362 22400 21418 22409
rect 21362 22335 21418 22344
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21088 19440 21140 19446
rect 21088 19382 21140 19388
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 20812 18420 20864 18426
rect 21008 18408 21036 18566
rect 20864 18380 21036 18408
rect 20812 18362 20864 18368
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 20902 17912 20958 17921
rect 20902 17847 20904 17856
rect 20956 17847 20958 17856
rect 20904 17818 20956 17824
rect 21008 17542 21036 18226
rect 21100 17746 21128 19382
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 21192 17626 21220 19654
rect 21284 19553 21312 19790
rect 21270 19544 21326 19553
rect 21270 19479 21326 19488
rect 21376 19446 21404 21082
rect 21468 20806 21496 37606
rect 21560 36378 21588 39200
rect 21824 38072 21876 38078
rect 21824 38014 21876 38020
rect 21548 36372 21600 36378
rect 21548 36314 21600 36320
rect 21836 35894 21864 38014
rect 21928 37176 21956 39200
rect 22100 37188 22152 37194
rect 21928 37148 22100 37176
rect 22100 37130 22152 37136
rect 21836 35866 21956 35894
rect 21548 33108 21600 33114
rect 21548 33050 21600 33056
rect 21560 23254 21588 33050
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21548 23248 21600 23254
rect 21548 23190 21600 23196
rect 21640 23248 21692 23254
rect 21640 23190 21692 23196
rect 21652 21185 21680 23190
rect 21744 21350 21772 24142
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21638 21176 21694 21185
rect 21638 21111 21694 21120
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21364 19440 21416 19446
rect 21100 17598 21220 17626
rect 21284 19388 21364 19394
rect 21284 19382 21416 19388
rect 21284 19366 21404 19382
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 20810 17368 20866 17377
rect 20810 17303 20866 17312
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20824 15745 20852 17303
rect 21008 16998 21036 17478
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20916 16250 20944 16730
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20810 15736 20866 15745
rect 20810 15671 20866 15680
rect 20916 15638 20944 16186
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 20904 15632 20956 15638
rect 20590 15558 20668 15586
rect 20534 15535 20590 15544
rect 20640 15434 20668 15558
rect 20718 15600 20774 15609
rect 20904 15574 20956 15580
rect 20718 15535 20720 15544
rect 20772 15535 20774 15544
rect 20720 15506 20772 15512
rect 21008 15450 21036 15982
rect 20628 15428 20680 15434
rect 20628 15370 20680 15376
rect 20732 15422 21036 15450
rect 20456 15286 20668 15314
rect 19982 15127 20038 15136
rect 19432 14884 19484 14890
rect 19260 14844 19432 14872
rect 19154 14648 19210 14657
rect 19154 14583 19210 14592
rect 19260 14498 19288 14844
rect 19432 14826 19484 14832
rect 19536 14793 19564 15116
rect 20272 15116 20392 15144
rect 20536 15156 20588 15162
rect 19892 15088 19944 15094
rect 19892 15030 19944 15036
rect 19616 14952 19668 14958
rect 19616 14894 19668 14900
rect 19522 14784 19578 14793
rect 19522 14719 19578 14728
rect 19628 14618 19656 14894
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19168 14470 19288 14498
rect 19168 14113 19196 14470
rect 19720 14414 19748 14758
rect 19904 14600 19932 15030
rect 19984 15020 20036 15026
rect 20168 15020 20220 15026
rect 20036 14980 20116 15008
rect 19984 14962 20036 14968
rect 19984 14612 20036 14618
rect 19904 14572 19984 14600
rect 19248 14408 19300 14414
rect 19432 14408 19484 14414
rect 19300 14368 19380 14396
rect 19248 14350 19300 14356
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19154 14104 19210 14113
rect 19260 14074 19288 14214
rect 19154 14039 19210 14048
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 18880 13796 18932 13802
rect 18880 13738 18932 13744
rect 18984 13790 19104 13818
rect 18892 13394 18920 13738
rect 18880 13388 18932 13394
rect 18880 13330 18932 13336
rect 18880 13252 18932 13258
rect 18880 13194 18932 13200
rect 18892 13161 18920 13194
rect 18878 13152 18934 13161
rect 18878 13087 18934 13096
rect 18984 12730 19012 13790
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19076 12850 19104 13670
rect 19168 12986 19196 13670
rect 19246 13560 19302 13569
rect 19246 13495 19302 13504
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19260 12918 19288 13495
rect 19352 12986 19380 14368
rect 19432 14350 19484 14356
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19444 14249 19472 14350
rect 19904 14260 19932 14572
rect 19984 14554 20036 14560
rect 20088 14550 20116 14980
rect 20168 14962 20220 14968
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 20180 14278 20208 14962
rect 20168 14272 20220 14278
rect 19430 14240 19486 14249
rect 19904 14232 19950 14260
rect 19430 14175 19486 14184
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19922 14056 19950 14232
rect 20074 14240 20130 14249
rect 20168 14214 20220 14220
rect 20074 14175 20130 14184
rect 19812 14028 19950 14056
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19706 13832 19762 13841
rect 19444 13530 19472 13806
rect 19524 13796 19576 13802
rect 19706 13767 19708 13776
rect 19524 13738 19576 13744
rect 19760 13767 19762 13776
rect 19708 13738 19760 13744
rect 19536 13705 19564 13738
rect 19522 13696 19578 13705
rect 19522 13631 19578 13640
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19340 12776 19392 12782
rect 18984 12702 19104 12730
rect 19340 12718 19392 12724
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18984 12084 19012 12582
rect 19076 12442 19104 12702
rect 19064 12436 19116 12442
rect 19352 12424 19380 12718
rect 19444 12646 19472 13466
rect 19524 13456 19576 13462
rect 19576 13404 19748 13410
rect 19524 13398 19748 13404
rect 19536 13394 19748 13398
rect 19536 13388 19760 13394
rect 19536 13382 19708 13388
rect 19708 13330 19760 13336
rect 19812 13172 19840 14028
rect 20088 13938 20116 14175
rect 20180 13938 20208 14214
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20272 13870 20300 15116
rect 20536 15098 20588 15104
rect 20350 15056 20406 15065
rect 20350 14991 20406 15000
rect 20364 14550 20392 14991
rect 20444 14884 20496 14890
rect 20444 14826 20496 14832
rect 20456 14618 20484 14826
rect 20548 14793 20576 15098
rect 20534 14784 20590 14793
rect 20534 14719 20590 14728
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20352 14068 20404 14074
rect 20640 14056 20668 15286
rect 20352 14010 20404 14016
rect 20456 14028 20668 14056
rect 20260 13864 20312 13870
rect 19982 13832 20038 13841
rect 19982 13767 20038 13776
rect 20166 13832 20222 13841
rect 20260 13806 20312 13812
rect 20166 13767 20168 13776
rect 19812 13144 19950 13172
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19922 12968 19950 13144
rect 19904 12940 19950 12968
rect 19708 12912 19760 12918
rect 19706 12880 19708 12889
rect 19760 12880 19762 12889
rect 19706 12815 19762 12824
rect 19904 12764 19932 12940
rect 19996 12918 20024 13767
rect 20220 13767 20222 13776
rect 20168 13738 20220 13744
rect 20364 13682 20392 14010
rect 20180 13654 20392 13682
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19904 12736 20024 12764
rect 19432 12640 19484 12646
rect 19616 12640 19668 12646
rect 19432 12582 19484 12588
rect 19614 12608 19616 12617
rect 19668 12608 19670 12617
rect 19614 12543 19670 12552
rect 19064 12378 19116 12384
rect 19168 12396 19380 12424
rect 19432 12436 19484 12442
rect 19168 12322 19196 12396
rect 19432 12378 19484 12384
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 18708 11614 18828 11642
rect 18892 12056 19012 12084
rect 19076 12294 19196 12322
rect 19340 12300 19392 12306
rect 18708 11082 18736 11614
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18800 11014 18828 11494
rect 18892 11150 18920 12056
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18708 10062 18736 10610
rect 18984 10606 19012 11698
rect 19076 10985 19104 12294
rect 19340 12242 19392 12248
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19168 11694 19196 12174
rect 19352 12170 19380 12242
rect 19444 12238 19472 12378
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19062 10976 19118 10985
rect 19062 10911 19118 10920
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18880 10532 18932 10538
rect 18880 10474 18932 10480
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18696 10056 18748 10062
rect 18800 10033 18828 10406
rect 18696 9998 18748 10004
rect 18786 10024 18842 10033
rect 18786 9959 18842 9968
rect 18616 9880 18736 9908
rect 18510 9752 18566 9761
rect 18510 9687 18566 9696
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 18524 9178 18552 9590
rect 18602 9480 18658 9489
rect 18602 9415 18658 9424
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18512 8900 18564 8906
rect 18512 8842 18564 8848
rect 18524 8498 18552 8842
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18432 5794 18460 7414
rect 18248 5766 18460 5794
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18248 4826 18276 5766
rect 18524 5574 18552 8434
rect 18616 8294 18644 9415
rect 18708 9110 18736 9880
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18694 8528 18750 8537
rect 18694 8463 18696 8472
rect 18748 8463 18750 8472
rect 18696 8434 18748 8440
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18602 8120 18658 8129
rect 18602 8055 18604 8064
rect 18656 8055 18658 8064
rect 18604 8026 18656 8032
rect 18616 7478 18644 8026
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18616 6474 18644 6734
rect 18616 6446 18736 6474
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18326 5400 18382 5409
rect 18326 5335 18382 5344
rect 18420 5364 18472 5370
rect 18340 5302 18368 5335
rect 18420 5306 18472 5312
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 17866 1728 17922 1737
rect 17866 1663 17922 1672
rect 17868 1556 17920 1562
rect 17868 1498 17920 1504
rect 17696 1142 17816 1170
rect 17696 800 17724 1142
rect 16856 740 16908 746
rect 16856 682 16908 688
rect 17038 0 17094 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 17880 406 17908 1498
rect 18156 1154 18184 3470
rect 18248 2689 18276 4082
rect 18234 2680 18290 2689
rect 18234 2615 18290 2624
rect 17960 1148 18012 1154
rect 17960 1090 18012 1096
rect 18144 1148 18196 1154
rect 18144 1090 18196 1096
rect 17972 950 18000 1090
rect 18156 1034 18184 1090
rect 18064 1006 18184 1034
rect 17960 944 18012 950
rect 17960 886 18012 892
rect 18064 800 18092 1006
rect 18340 800 18368 4082
rect 18432 1766 18460 5306
rect 18512 4548 18564 4554
rect 18512 4490 18564 4496
rect 18524 4146 18552 4490
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18616 3398 18644 6258
rect 18708 3641 18736 6446
rect 18800 5914 18828 9454
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18892 3738 18920 10474
rect 18972 10192 19024 10198
rect 18972 10134 19024 10140
rect 18984 8809 19012 10134
rect 19064 9716 19116 9722
rect 19168 9704 19196 11018
rect 19260 10849 19288 12106
rect 19352 11830 19380 12106
rect 19536 12084 19564 12378
rect 19706 12336 19762 12345
rect 19706 12271 19708 12280
rect 19760 12271 19762 12280
rect 19708 12242 19760 12248
rect 19444 12073 19564 12084
rect 19430 12064 19564 12073
rect 19486 12056 19564 12064
rect 19430 11999 19486 12008
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19340 11824 19392 11830
rect 19708 11824 19760 11830
rect 19340 11766 19392 11772
rect 19430 11792 19486 11801
rect 19430 11727 19486 11736
rect 19614 11792 19670 11801
rect 19708 11766 19760 11772
rect 19614 11727 19670 11736
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19246 10840 19302 10849
rect 19246 10775 19302 10784
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19260 10062 19288 10678
rect 19352 10282 19380 11290
rect 19444 10810 19472 11727
rect 19628 11558 19656 11727
rect 19720 11694 19748 11766
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19720 11354 19748 11494
rect 19904 11393 19932 11698
rect 19890 11384 19946 11393
rect 19708 11348 19760 11354
rect 19890 11319 19946 11328
rect 19708 11290 19760 11296
rect 19996 11234 20024 12736
rect 20088 11558 20116 13126
rect 20180 11762 20208 13654
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 12646 20300 13262
rect 20456 12866 20484 14028
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20364 12838 20484 12866
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20364 12374 20392 12838
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 12646 20484 12718
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20352 12368 20404 12374
rect 20352 12310 20404 12316
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20272 11665 20300 11834
rect 20258 11656 20314 11665
rect 20258 11591 20314 11600
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20074 11384 20130 11393
rect 20074 11319 20076 11328
rect 20128 11319 20130 11328
rect 20076 11290 20128 11296
rect 19996 11206 20116 11234
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19982 10840 20038 10849
rect 19432 10804 19484 10810
rect 19982 10775 19984 10784
rect 19432 10746 19484 10752
rect 20036 10775 20038 10784
rect 19984 10746 20036 10752
rect 19890 10704 19946 10713
rect 20088 10690 20116 11206
rect 20258 11112 20314 11121
rect 20168 11076 20220 11082
rect 20258 11047 20260 11056
rect 20168 11018 20220 11024
rect 20312 11047 20314 11056
rect 20260 11018 20312 11024
rect 19890 10639 19946 10648
rect 19996 10662 20116 10690
rect 19904 10538 19932 10639
rect 19892 10532 19944 10538
rect 19892 10474 19944 10480
rect 19352 10254 19472 10282
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19168 9676 19288 9704
rect 19064 9658 19116 9664
rect 19076 9602 19104 9658
rect 19076 9574 19196 9602
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 19076 9081 19104 9454
rect 19168 9217 19196 9574
rect 19260 9518 19288 9676
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19154 9208 19210 9217
rect 19154 9143 19210 9152
rect 19062 9072 19118 9081
rect 19062 9007 19118 9016
rect 18970 8800 19026 8809
rect 18970 8735 19026 8744
rect 19154 8664 19210 8673
rect 19154 8599 19156 8608
rect 19208 8599 19210 8608
rect 19156 8570 19208 8576
rect 19260 8566 19288 9454
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 18970 8120 19026 8129
rect 18970 8055 19026 8064
rect 19156 8084 19208 8090
rect 18984 7721 19012 8055
rect 19156 8026 19208 8032
rect 18970 7712 19026 7721
rect 18970 7647 19026 7656
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18972 5840 19024 5846
rect 18972 5782 19024 5788
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18694 3632 18750 3641
rect 18694 3567 18750 3576
rect 18984 3534 19012 5782
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18524 2009 18552 2382
rect 18510 2000 18566 2009
rect 18510 1935 18566 1944
rect 18420 1760 18472 1766
rect 18420 1702 18472 1708
rect 18708 800 18736 2790
rect 18984 800 19012 3470
rect 19076 3058 19104 6734
rect 19168 6254 19196 8026
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 19260 6730 19288 7414
rect 19248 6724 19300 6730
rect 19248 6666 19300 6672
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19260 5914 19288 6666
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19352 5794 19380 10134
rect 19444 9926 19472 10254
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19430 9752 19486 9761
rect 19574 9744 19882 9764
rect 19996 9704 20024 10662
rect 20074 10160 20130 10169
rect 20074 10095 20130 10104
rect 19486 9696 19564 9704
rect 19430 9687 19564 9696
rect 19444 9676 19564 9687
rect 19536 9489 19564 9676
rect 19812 9676 20024 9704
rect 19522 9480 19578 9489
rect 19522 9415 19578 9424
rect 19812 8820 19840 9676
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 19904 9081 19932 9386
rect 20088 9178 20116 10095
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19984 9104 20036 9110
rect 19890 9072 19946 9081
rect 19984 9046 20036 9052
rect 19890 9007 19946 9016
rect 19812 8792 19950 8820
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19922 8616 19950 8792
rect 19996 8673 20024 9046
rect 20076 8900 20128 8906
rect 20180 8888 20208 11018
rect 20364 10674 20392 12310
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20456 12102 20484 12174
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20548 11694 20576 13874
rect 20628 13456 20680 13462
rect 20628 13398 20680 13404
rect 20640 13326 20668 13398
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20732 13190 20760 15422
rect 20994 15328 21050 15337
rect 20994 15263 21050 15272
rect 20810 15192 20866 15201
rect 20810 15127 20812 15136
rect 20864 15127 20866 15136
rect 20812 15098 20864 15104
rect 21008 15026 21036 15263
rect 21100 15042 21128 17598
rect 21284 17202 21312 19366
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21376 18426 21404 19110
rect 21468 18902 21496 20742
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 21560 18970 21588 19722
rect 21652 19718 21680 20334
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 21456 18896 21508 18902
rect 21456 18838 21508 18844
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21454 18456 21510 18465
rect 21364 18420 21416 18426
rect 21454 18391 21456 18400
rect 21364 18362 21416 18368
rect 21508 18391 21510 18400
rect 21456 18362 21508 18368
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 21376 17678 21404 18158
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21376 17542 21404 17614
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21180 17060 21232 17066
rect 21180 17002 21232 17008
rect 21192 16590 21220 17002
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21284 16454 21312 16594
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 21192 15162 21220 15846
rect 21284 15570 21312 16390
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21270 15464 21326 15473
rect 21270 15399 21272 15408
rect 21324 15399 21326 15408
rect 21272 15370 21324 15376
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 20996 15020 21048 15026
rect 21100 15014 21220 15042
rect 20996 14962 21048 14968
rect 20812 14952 20864 14958
rect 21008 14929 21036 14962
rect 20812 14894 20864 14900
rect 20994 14920 21050 14929
rect 20824 14657 20852 14894
rect 20994 14855 21050 14864
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 20810 14648 20866 14657
rect 20810 14583 20866 14592
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20824 14113 20852 14350
rect 20810 14104 20866 14113
rect 20810 14039 20866 14048
rect 20824 13705 20852 14039
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20810 13696 20866 13705
rect 20810 13631 20866 13640
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12986 20760 13126
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20628 12912 20680 12918
rect 20628 12854 20680 12860
rect 20640 12481 20668 12854
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20626 12472 20682 12481
rect 20626 12407 20682 12416
rect 20626 12200 20682 12209
rect 20626 12135 20682 12144
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 20640 11234 20668 12135
rect 20732 11898 20760 12582
rect 20916 12434 20944 13874
rect 20824 12406 20944 12434
rect 20824 12073 20852 12406
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 20810 12064 20866 12073
rect 20810 11999 20866 12008
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20548 11206 20668 11234
rect 20732 11218 20760 11698
rect 20810 11656 20866 11665
rect 20810 11591 20812 11600
rect 20864 11591 20866 11600
rect 20812 11562 20864 11568
rect 20720 11212 20772 11218
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20272 8906 20300 10542
rect 20456 10520 20484 11018
rect 20548 10985 20576 11206
rect 20720 11154 20772 11160
rect 20628 11144 20680 11150
rect 20916 11098 20944 12310
rect 21008 12209 21036 14758
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 21100 14113 21128 14282
rect 21086 14104 21142 14113
rect 21086 14039 21142 14048
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 21100 13394 21128 13942
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 21192 12918 21220 15014
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21284 14464 21312 14962
rect 21376 14890 21404 17478
rect 21560 16658 21588 18702
rect 21640 18692 21692 18698
rect 21640 18634 21692 18640
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21456 16176 21508 16182
rect 21456 16118 21508 16124
rect 21364 14884 21416 14890
rect 21364 14826 21416 14832
rect 21468 14498 21496 16118
rect 21548 16108 21600 16114
rect 21548 16050 21600 16056
rect 21560 15706 21588 16050
rect 21652 15745 21680 18634
rect 21744 18358 21772 21286
rect 21928 20330 21956 35866
rect 22112 35834 22140 37130
rect 22388 36922 22416 39200
rect 22560 37732 22612 37738
rect 22560 37674 22612 37680
rect 22572 37398 22600 37674
rect 22468 37392 22520 37398
rect 22468 37334 22520 37340
rect 22560 37392 22612 37398
rect 22560 37334 22612 37340
rect 22376 36916 22428 36922
rect 22376 36858 22428 36864
rect 22192 36168 22244 36174
rect 22192 36110 22244 36116
rect 22100 35828 22152 35834
rect 22100 35770 22152 35776
rect 22204 35222 22232 36110
rect 22376 35284 22428 35290
rect 22376 35226 22428 35232
rect 22192 35216 22244 35222
rect 22192 35158 22244 35164
rect 22098 26480 22154 26489
rect 22098 26415 22154 26424
rect 22112 24410 22140 26415
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 22112 23798 22140 24346
rect 22100 23792 22152 23798
rect 22100 23734 22152 23740
rect 22190 23080 22246 23089
rect 22190 23015 22246 23024
rect 22284 23044 22336 23050
rect 22204 22710 22232 23015
rect 22284 22986 22336 22992
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 22006 22264 22062 22273
rect 22204 22234 22232 22646
rect 22006 22199 22062 22208
rect 22192 22228 22244 22234
rect 22020 22114 22048 22199
rect 22192 22170 22244 22176
rect 22020 22086 22140 22114
rect 21916 20324 21968 20330
rect 21916 20266 21968 20272
rect 22006 19544 22062 19553
rect 22006 19479 22062 19488
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 21836 18737 21864 19246
rect 21822 18728 21878 18737
rect 21822 18663 21878 18672
rect 21732 18352 21784 18358
rect 21732 18294 21784 18300
rect 21744 17921 21772 18294
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21730 17912 21786 17921
rect 21730 17847 21786 17856
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21744 17202 21772 17546
rect 21732 17196 21784 17202
rect 21732 17138 21784 17144
rect 21638 15736 21694 15745
rect 21548 15700 21600 15706
rect 21638 15671 21694 15680
rect 21548 15642 21600 15648
rect 21640 15632 21692 15638
rect 21546 15600 21602 15609
rect 21640 15574 21692 15580
rect 21546 15535 21602 15544
rect 21560 15502 21588 15535
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21468 14470 21588 14498
rect 21284 14436 21404 14464
rect 21270 14376 21326 14385
rect 21270 14311 21272 14320
rect 21324 14311 21326 14320
rect 21272 14282 21324 14288
rect 21376 14226 21404 14436
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21284 14198 21404 14226
rect 21284 13530 21312 14198
rect 21468 13977 21496 14350
rect 21454 13968 21510 13977
rect 21454 13903 21510 13912
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21180 12912 21232 12918
rect 21180 12854 21232 12860
rect 21088 12708 21140 12714
rect 21088 12650 21140 12656
rect 20994 12200 21050 12209
rect 20994 12135 21050 12144
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 21008 11626 21036 11698
rect 20996 11620 21048 11626
rect 20996 11562 21048 11568
rect 21100 11354 21128 12650
rect 21178 12608 21234 12617
rect 21178 12543 21234 12552
rect 21192 12434 21220 12543
rect 21192 12406 21312 12434
rect 21180 12164 21232 12170
rect 21180 12106 21232 12112
rect 21192 12073 21220 12106
rect 21178 12064 21234 12073
rect 21178 11999 21234 12008
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 20628 11086 20680 11092
rect 20640 11014 20668 11086
rect 20732 11070 20944 11098
rect 20994 11112 21050 11121
rect 20628 11008 20680 11014
rect 20534 10976 20590 10985
rect 20628 10950 20680 10956
rect 20534 10911 20590 10920
rect 20536 10532 20588 10538
rect 20456 10492 20536 10520
rect 20536 10474 20588 10480
rect 20536 10192 20588 10198
rect 20534 10160 20536 10169
rect 20588 10160 20590 10169
rect 20534 10095 20590 10104
rect 20352 10056 20404 10062
rect 20404 10016 20484 10044
rect 20352 9998 20404 10004
rect 20352 9648 20404 9654
rect 20352 9590 20404 9596
rect 20364 8906 20392 9590
rect 20128 8860 20208 8888
rect 20260 8900 20312 8906
rect 20076 8842 20128 8848
rect 20260 8842 20312 8848
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 20272 8786 20300 8842
rect 20088 8758 20300 8786
rect 19904 8588 19950 8616
rect 19982 8664 20038 8673
rect 19982 8599 20038 8608
rect 19904 8362 19932 8588
rect 20088 8566 20116 8758
rect 20364 8650 20392 8842
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 20272 8622 20392 8650
rect 20076 8560 20128 8566
rect 20076 8502 20128 8508
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19536 8265 19564 8298
rect 19522 8256 19578 8265
rect 19522 8191 19578 8200
rect 19800 7880 19852 7886
rect 19798 7848 19800 7857
rect 19852 7848 19854 7857
rect 19798 7783 19854 7792
rect 20088 7750 20116 8502
rect 20076 7744 20128 7750
rect 19982 7712 20038 7721
rect 19574 7644 19882 7664
rect 20076 7686 20128 7692
rect 19982 7647 20038 7656
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19430 7440 19486 7449
rect 19430 7375 19432 7384
rect 19484 7375 19486 7384
rect 19432 7346 19484 7352
rect 19996 7206 20024 7647
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19720 6769 19748 6802
rect 19706 6760 19762 6769
rect 19524 6724 19576 6730
rect 19260 5766 19380 5794
rect 19444 6684 19524 6712
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19168 2774 19196 4014
rect 19260 3942 19288 5766
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19352 4010 19380 5578
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19338 3496 19394 3505
rect 19444 3466 19472 6684
rect 19706 6695 19762 6704
rect 19524 6666 19576 6672
rect 20074 6624 20130 6633
rect 19574 6556 19882 6576
rect 20074 6559 20130 6568
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19982 6488 20038 6497
rect 19982 6423 20038 6432
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 19720 5681 19748 6326
rect 19706 5672 19762 5681
rect 19706 5607 19762 5616
rect 19812 5556 19840 6326
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19904 5914 19932 6258
rect 19996 6186 20024 6423
rect 20088 6361 20116 6559
rect 20074 6352 20130 6361
rect 20074 6287 20130 6296
rect 20076 6248 20128 6254
rect 20076 6190 20128 6196
rect 19984 6180 20036 6186
rect 19984 6122 20036 6128
rect 19892 5908 19944 5914
rect 19892 5850 19944 5856
rect 19812 5528 20024 5556
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19536 4690 19564 5238
rect 19996 4826 20024 5528
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19996 3602 20024 4422
rect 20088 3602 20116 6190
rect 20180 3738 20208 8570
rect 20272 8430 20300 8622
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 20272 7410 20300 8366
rect 20352 8356 20404 8362
rect 20352 8298 20404 8304
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 5080 20300 6598
rect 20364 6458 20392 8298
rect 20456 7002 20484 10016
rect 20628 9988 20680 9994
rect 20548 9948 20628 9976
rect 20548 9897 20576 9948
rect 20628 9930 20680 9936
rect 20534 9888 20590 9897
rect 20534 9823 20590 9832
rect 20732 9654 20760 11070
rect 20994 11047 21050 11056
rect 21088 11076 21140 11082
rect 20810 10976 20866 10985
rect 20810 10911 20866 10920
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20824 9466 20852 10911
rect 21008 10470 21036 11047
rect 21088 11018 21140 11024
rect 20996 10464 21048 10470
rect 20902 10432 20958 10441
rect 20996 10406 21048 10412
rect 20902 10367 20958 10376
rect 20916 9897 20944 10367
rect 20902 9888 20958 9897
rect 20902 9823 20958 9832
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20548 9438 20852 9466
rect 20548 9178 20576 9438
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20640 8401 20668 9318
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 20626 8392 20682 8401
rect 20536 8356 20588 8362
rect 20824 8362 20852 9046
rect 20626 8327 20682 8336
rect 20812 8356 20864 8362
rect 20536 8298 20588 8304
rect 20812 8298 20864 8304
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20350 6352 20406 6361
rect 20350 6287 20406 6296
rect 20364 5778 20392 6287
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20272 5052 20484 5080
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20260 4004 20312 4010
rect 20260 3946 20312 3952
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 19338 3431 19340 3440
rect 19392 3431 19394 3440
rect 19432 3460 19484 3466
rect 19340 3402 19392 3408
rect 19432 3402 19484 3408
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19168 2746 19288 2774
rect 19260 800 19288 2746
rect 19904 2650 19932 2858
rect 19892 2644 19944 2650
rect 19892 2586 19944 2592
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19444 1170 19472 2246
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 2020 20024 2994
rect 19904 1992 20024 2020
rect 19444 1142 19656 1170
rect 19628 800 19656 1142
rect 19904 800 19932 1992
rect 20272 1562 20300 3946
rect 20364 3534 20392 4558
rect 20456 4049 20484 5052
rect 20442 4040 20498 4049
rect 20442 3975 20498 3984
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20456 3670 20484 3878
rect 20444 3664 20496 3670
rect 20444 3606 20496 3612
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20364 2774 20392 3470
rect 20548 3194 20576 8298
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20640 6905 20668 7142
rect 20732 6934 20760 7278
rect 20720 6928 20772 6934
rect 20626 6896 20682 6905
rect 20720 6870 20772 6876
rect 20626 6831 20682 6840
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20640 6458 20668 6734
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20640 3058 20668 5306
rect 20732 4457 20760 6054
rect 20718 4448 20774 4457
rect 20718 4383 20774 4392
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20732 3126 20760 3606
rect 20720 3120 20772 3126
rect 20720 3062 20772 3068
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20364 2746 20576 2774
rect 20548 2394 20576 2746
rect 20824 2446 20852 7686
rect 20916 3194 20944 9522
rect 21008 9042 21036 10406
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 21008 3738 21036 8298
rect 21100 7993 21128 11018
rect 21178 10296 21234 10305
rect 21178 10231 21234 10240
rect 21192 9994 21220 10231
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 21178 9888 21234 9897
rect 21178 9823 21234 9832
rect 21086 7984 21142 7993
rect 21086 7919 21142 7928
rect 21192 7868 21220 9823
rect 21284 8498 21312 12406
rect 21376 11150 21404 13330
rect 21454 13288 21510 13297
rect 21454 13223 21456 13232
rect 21508 13223 21510 13232
rect 21456 13194 21508 13200
rect 21454 12064 21510 12073
rect 21454 11999 21510 12008
rect 21364 11144 21416 11150
rect 21468 11121 21496 11999
rect 21560 11830 21588 14470
rect 21548 11824 21600 11830
rect 21548 11766 21600 11772
rect 21364 11086 21416 11092
rect 21454 11112 21510 11121
rect 21454 11047 21510 11056
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21376 8945 21404 10542
rect 21560 10266 21588 11018
rect 21652 10810 21680 15574
rect 21744 14618 21772 17138
rect 21822 16688 21878 16697
rect 21822 16623 21878 16632
rect 21836 16250 21864 16623
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21928 15026 21956 18022
rect 22020 16697 22048 19479
rect 22112 16833 22140 22086
rect 22296 22094 22324 22986
rect 22388 22778 22416 35226
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 22296 22066 22416 22094
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22296 21350 22324 21558
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22192 20800 22244 20806
rect 22190 20768 22192 20777
rect 22244 20768 22246 20777
rect 22190 20703 22246 20712
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22204 17882 22232 19994
rect 22296 18358 22324 21286
rect 22388 18850 22416 22066
rect 22480 20806 22508 37334
rect 22652 36780 22704 36786
rect 22652 36722 22704 36728
rect 22664 35766 22692 36722
rect 22756 36378 22784 39200
rect 23216 37262 23244 39200
rect 23204 37256 23256 37262
rect 23204 37198 23256 37204
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 23204 36780 23256 36786
rect 23204 36722 23256 36728
rect 22744 36372 22796 36378
rect 22744 36314 22796 36320
rect 22652 35760 22704 35766
rect 22652 35702 22704 35708
rect 23216 35494 23244 36722
rect 23400 36378 23428 37198
rect 23584 36922 23612 39200
rect 23848 37800 23900 37806
rect 23848 37742 23900 37748
rect 23572 36916 23624 36922
rect 23572 36858 23624 36864
rect 23664 36780 23716 36786
rect 23664 36722 23716 36728
rect 23388 36372 23440 36378
rect 23388 36314 23440 36320
rect 23296 36168 23348 36174
rect 23296 36110 23348 36116
rect 23388 36168 23440 36174
rect 23388 36110 23440 36116
rect 23204 35488 23256 35494
rect 23204 35430 23256 35436
rect 22836 34604 22888 34610
rect 22836 34546 22888 34552
rect 22744 34536 22796 34542
rect 22744 34478 22796 34484
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22572 18970 22600 22578
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22664 20806 22692 20946
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22650 20632 22706 20641
rect 22650 20567 22652 20576
rect 22704 20567 22706 20576
rect 22652 20538 22704 20544
rect 22756 19378 22784 34478
rect 22848 19922 22876 34546
rect 23216 33862 23244 35430
rect 23308 34950 23336 36110
rect 23400 34950 23428 36110
rect 23676 35494 23704 36722
rect 23664 35488 23716 35494
rect 23664 35430 23716 35436
rect 23296 34944 23348 34950
rect 23296 34886 23348 34892
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23204 33856 23256 33862
rect 23204 33798 23256 33804
rect 23308 29481 23336 34886
rect 23400 34542 23428 34886
rect 23676 34678 23704 35430
rect 23664 34672 23716 34678
rect 23664 34614 23716 34620
rect 23388 34536 23440 34542
rect 23388 34478 23440 34484
rect 23860 31754 23888 37742
rect 23952 36378 23980 39200
rect 24308 37664 24360 37670
rect 24308 37606 24360 37612
rect 23940 36372 23992 36378
rect 23940 36314 23992 36320
rect 24216 35148 24268 35154
rect 24216 35090 24268 35096
rect 23676 31726 23888 31754
rect 23294 29472 23350 29481
rect 23294 29407 23350 29416
rect 23202 26072 23258 26081
rect 23202 26007 23258 26016
rect 23020 25220 23072 25226
rect 23020 25162 23072 25168
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 22940 21622 22968 24754
rect 22928 21616 22980 21622
rect 22928 21558 22980 21564
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22744 19372 22796 19378
rect 22744 19314 22796 19320
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22388 18822 22508 18850
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22284 18352 22336 18358
rect 22284 18294 22336 18300
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22098 16824 22154 16833
rect 22098 16759 22154 16768
rect 22006 16688 22062 16697
rect 22006 16623 22062 16632
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22008 16516 22060 16522
rect 22008 16458 22060 16464
rect 22020 15434 22048 16458
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 22020 15201 22048 15370
rect 22006 15192 22062 15201
rect 22006 15127 22062 15136
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21822 14784 21878 14793
rect 21822 14719 21878 14728
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21744 13433 21772 14350
rect 21836 13870 21864 14719
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 21916 13728 21968 13734
rect 21916 13670 21968 13676
rect 21822 13560 21878 13569
rect 21822 13495 21878 13504
rect 21730 13424 21786 13433
rect 21730 13359 21786 13368
rect 21732 13252 21784 13258
rect 21732 13194 21784 13200
rect 21744 12753 21772 13194
rect 21836 13025 21864 13495
rect 21928 13462 21956 13670
rect 21916 13456 21968 13462
rect 21916 13398 21968 13404
rect 21916 13252 21968 13258
rect 21916 13194 21968 13200
rect 21928 13161 21956 13194
rect 21914 13152 21970 13161
rect 21914 13087 21970 13096
rect 21822 13016 21878 13025
rect 21822 12951 21878 12960
rect 21730 12744 21786 12753
rect 21730 12679 21786 12688
rect 22020 12594 22048 14554
rect 22112 14278 22140 16594
rect 22204 15026 22232 16934
rect 22296 15638 22324 17274
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22388 15570 22416 18702
rect 22480 17649 22508 18822
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22664 17814 22692 18634
rect 22652 17808 22704 17814
rect 22652 17750 22704 17756
rect 22466 17640 22522 17649
rect 22466 17575 22522 17584
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22466 17096 22522 17105
rect 22466 17031 22522 17040
rect 22480 16833 22508 17031
rect 22466 16824 22522 16833
rect 22466 16759 22522 16768
rect 22480 16726 22508 16759
rect 22468 16720 22520 16726
rect 22468 16662 22520 16668
rect 22572 16658 22600 17138
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22466 16552 22522 16561
rect 22466 16487 22522 16496
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 22480 15450 22508 16487
rect 22560 15972 22612 15978
rect 22560 15914 22612 15920
rect 22296 15422 22508 15450
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 22100 13796 22152 13802
rect 22204 13784 22232 14486
rect 22152 13756 22232 13784
rect 22100 13738 22152 13744
rect 22098 13560 22154 13569
rect 22098 13495 22100 13504
rect 22152 13495 22154 13504
rect 22100 13466 22152 13472
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 21928 12566 22048 12594
rect 21732 12368 21784 12374
rect 21732 12310 21784 12316
rect 21744 12238 21772 12310
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21822 12200 21878 12209
rect 21822 12135 21878 12144
rect 21836 11898 21864 12135
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 21732 11620 21784 11626
rect 21732 11562 21784 11568
rect 21640 10804 21692 10810
rect 21640 10746 21692 10752
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21362 8936 21418 8945
rect 21362 8871 21418 8880
rect 21468 8809 21496 9318
rect 21454 8800 21510 8809
rect 21454 8735 21510 8744
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 21100 7840 21220 7868
rect 21100 6202 21128 7840
rect 21284 7818 21312 8298
rect 21454 8256 21510 8265
rect 21454 8191 21510 8200
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21364 7812 21416 7818
rect 21364 7754 21416 7760
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21192 7324 21220 7482
rect 21284 7449 21312 7754
rect 21270 7440 21326 7449
rect 21270 7375 21326 7384
rect 21192 7296 21312 7324
rect 21284 6746 21312 7296
rect 21376 6866 21404 7754
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21284 6718 21404 6746
rect 21100 6174 21220 6202
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21100 5273 21128 6054
rect 21192 5914 21220 6174
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 21086 5264 21142 5273
rect 21086 5199 21142 5208
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 20364 2366 20576 2394
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20260 1556 20312 1562
rect 20260 1498 20312 1504
rect 20364 1442 20392 2366
rect 20536 2304 20588 2310
rect 20536 2246 20588 2252
rect 20272 1414 20392 1442
rect 20444 1420 20496 1426
rect 20168 1284 20220 1290
rect 20168 1226 20220 1232
rect 20180 1057 20208 1226
rect 20166 1048 20222 1057
rect 20166 983 20222 992
rect 20272 800 20300 1414
rect 20444 1362 20496 1368
rect 20456 1290 20484 1362
rect 20444 1284 20496 1290
rect 20444 1226 20496 1232
rect 20548 800 20576 2246
rect 20720 2100 20772 2106
rect 20720 2042 20772 2048
rect 20732 1601 20760 2042
rect 20718 1592 20774 1601
rect 20718 1527 20774 1536
rect 20916 800 20944 2994
rect 21100 2378 21128 3878
rect 21284 3534 21312 4626
rect 21376 3738 21404 6718
rect 21468 6254 21496 8191
rect 21560 7478 21588 10202
rect 21744 9926 21772 11562
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21652 8634 21680 8910
rect 21744 8634 21772 9522
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21652 7546 21680 7686
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21548 7472 21600 7478
rect 21548 7414 21600 7420
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21468 4282 21496 4422
rect 21456 4276 21508 4282
rect 21456 4218 21508 4224
rect 21560 4185 21588 4422
rect 21546 4176 21602 4185
rect 21652 4146 21680 6190
rect 21546 4111 21602 4120
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 21272 3528 21324 3534
rect 21272 3470 21324 3476
rect 21284 2774 21312 3470
rect 21192 2746 21312 2774
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 21192 800 21220 2746
rect 21744 2446 21772 6598
rect 21836 3194 21864 11698
rect 21928 11694 21956 12566
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 21916 11688 21968 11694
rect 21916 11630 21968 11636
rect 22020 10810 22048 11766
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22020 10606 22048 10746
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 21916 10464 21968 10470
rect 21914 10432 21916 10441
rect 21968 10432 21970 10441
rect 21914 10367 21970 10376
rect 22112 10282 22140 11766
rect 22204 10742 22232 12786
rect 22192 10736 22244 10742
rect 22192 10678 22244 10684
rect 21928 10254 22140 10282
rect 21928 9722 21956 10254
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21928 7993 21956 8230
rect 22020 8090 22048 9862
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22112 9450 22140 9658
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 22098 9208 22154 9217
rect 22098 9143 22100 9152
rect 22152 9143 22154 9152
rect 22100 9114 22152 9120
rect 22204 9081 22232 9862
rect 22190 9072 22246 9081
rect 22190 9007 22246 9016
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 21914 7984 21970 7993
rect 21914 7919 21970 7928
rect 21928 7886 21956 7919
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 22020 7410 22048 7822
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22112 7410 22140 7686
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22296 6905 22324 15422
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22388 14482 22416 15098
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22388 13734 22416 14418
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22388 9450 22416 13466
rect 22480 12238 22508 14282
rect 22572 13530 22600 15914
rect 22664 13938 22692 16934
rect 22756 16046 22784 18702
rect 22926 18456 22982 18465
rect 22926 18391 22928 18400
rect 22980 18391 22982 18400
rect 22928 18362 22980 18368
rect 23032 18290 23060 25162
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 23020 18284 23072 18290
rect 23020 18226 23072 18232
rect 23124 18170 23152 21558
rect 23216 21078 23244 26007
rect 23480 21480 23532 21486
rect 23478 21448 23480 21457
rect 23532 21448 23534 21457
rect 23478 21383 23534 21392
rect 23676 21350 23704 31726
rect 23848 25288 23900 25294
rect 23848 25230 23900 25236
rect 23756 21684 23808 21690
rect 23756 21626 23808 21632
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23204 21072 23256 21078
rect 23204 21014 23256 21020
rect 23204 20868 23256 20874
rect 23204 20810 23256 20816
rect 23216 19310 23244 20810
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 23204 19304 23256 19310
rect 23204 19246 23256 19252
rect 23216 18329 23244 19246
rect 23202 18320 23258 18329
rect 23308 18306 23336 20742
rect 23492 20618 23520 21286
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23400 20590 23520 20618
rect 23400 19854 23428 20590
rect 23676 20097 23704 20742
rect 23662 20088 23718 20097
rect 23662 20023 23718 20032
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23492 19689 23520 19722
rect 23478 19680 23534 19689
rect 23478 19615 23534 19624
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23386 18320 23442 18329
rect 23308 18278 23386 18306
rect 23202 18255 23258 18264
rect 23386 18255 23442 18264
rect 23296 18216 23348 18222
rect 23124 18142 23244 18170
rect 23296 18158 23348 18164
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 22940 17105 22968 17682
rect 23020 17604 23072 17610
rect 23020 17546 23072 17552
rect 22926 17096 22982 17105
rect 22926 17031 22982 17040
rect 23032 16998 23060 17546
rect 23216 17542 23244 18142
rect 23308 17785 23336 18158
rect 23492 18034 23520 18906
rect 23584 18426 23612 19382
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23400 18006 23520 18034
rect 23294 17776 23350 17785
rect 23294 17711 23350 17720
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23110 17232 23166 17241
rect 23110 17167 23166 17176
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 22940 16658 22968 16934
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 22836 16176 22888 16182
rect 22836 16118 22888 16124
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22756 15144 22784 15438
rect 22848 15337 22876 16118
rect 22928 15632 22980 15638
rect 22928 15574 22980 15580
rect 22834 15328 22890 15337
rect 22834 15263 22890 15272
rect 22756 15116 22876 15144
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 22756 14793 22784 14962
rect 22848 14958 22876 15116
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22836 14816 22888 14822
rect 22742 14784 22798 14793
rect 22836 14758 22888 14764
rect 22742 14719 22798 14728
rect 22756 14362 22784 14719
rect 22848 14550 22876 14758
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 22756 14334 22876 14362
rect 22742 14104 22798 14113
rect 22742 14039 22798 14048
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22650 13560 22706 13569
rect 22560 13524 22612 13530
rect 22650 13495 22706 13504
rect 22560 13466 22612 13472
rect 22558 13424 22614 13433
rect 22558 13359 22614 13368
rect 22572 13258 22600 13359
rect 22560 13252 22612 13258
rect 22560 13194 22612 13200
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22572 11506 22600 12854
rect 22664 11898 22692 13495
rect 22756 13433 22784 14039
rect 22742 13424 22798 13433
rect 22742 13359 22798 13368
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22848 11626 22876 14334
rect 22940 12782 22968 15574
rect 23032 12850 23060 16934
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 23124 12434 23152 17167
rect 23204 17128 23256 17134
rect 23204 17070 23256 17076
rect 23216 16946 23244 17070
rect 23400 17066 23428 18006
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23388 17060 23440 17066
rect 23388 17002 23440 17008
rect 23216 16918 23428 16946
rect 23294 16824 23350 16833
rect 23204 16788 23256 16794
rect 23294 16759 23350 16768
rect 23204 16730 23256 16736
rect 23216 16182 23244 16730
rect 23308 16590 23336 16759
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23308 16182 23336 16390
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23296 16176 23348 16182
rect 23296 16118 23348 16124
rect 23296 15428 23348 15434
rect 23216 15388 23296 15416
rect 23216 15094 23244 15388
rect 23296 15370 23348 15376
rect 23204 15088 23256 15094
rect 23204 15030 23256 15036
rect 23294 15056 23350 15065
rect 23216 14385 23244 15030
rect 23294 14991 23350 15000
rect 23308 14958 23336 14991
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23202 14376 23258 14385
rect 23202 14311 23258 14320
rect 23216 13326 23244 14311
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23032 12406 23152 12434
rect 22836 11620 22888 11626
rect 22836 11562 22888 11568
rect 22480 11478 22600 11506
rect 22480 11014 22508 11478
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22572 11121 22600 11290
rect 22836 11144 22888 11150
rect 22558 11112 22614 11121
rect 22836 11086 22888 11092
rect 22558 11047 22614 11056
rect 22744 11076 22796 11082
rect 22744 11018 22796 11024
rect 22468 11008 22520 11014
rect 22468 10950 22520 10956
rect 22480 10062 22508 10950
rect 22756 10742 22784 11018
rect 22744 10736 22796 10742
rect 22744 10678 22796 10684
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22376 9444 22428 9450
rect 22376 9386 22428 9392
rect 22468 9444 22520 9450
rect 22468 9386 22520 9392
rect 22388 8498 22416 9386
rect 22480 9110 22508 9386
rect 22664 9382 22692 10066
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22572 9217 22600 9318
rect 22558 9208 22614 9217
rect 22558 9143 22614 9152
rect 22468 9104 22520 9110
rect 22468 9046 22520 9052
rect 22558 9072 22614 9081
rect 22558 9007 22560 9016
rect 22612 9007 22614 9016
rect 22560 8978 22612 8984
rect 22572 8566 22600 8978
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22374 8120 22430 8129
rect 22374 8055 22430 8064
rect 22388 7954 22416 8055
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22664 7460 22692 9318
rect 22756 8634 22784 9522
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 22572 7432 22692 7460
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 21914 6896 21970 6905
rect 21914 6831 21970 6840
rect 22282 6896 22338 6905
rect 22282 6831 22338 6840
rect 21928 6390 21956 6831
rect 21916 6384 21968 6390
rect 21916 6326 21968 6332
rect 22190 5672 22246 5681
rect 22190 5607 22192 5616
rect 22244 5607 22246 5616
rect 22192 5578 22244 5584
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21732 2440 21784 2446
rect 21732 2382 21784 2388
rect 21456 2304 21508 2310
rect 21456 2246 21508 2252
rect 21468 800 21496 2246
rect 21836 800 21864 2994
rect 21928 2825 21956 5102
rect 21914 2816 21970 2825
rect 21914 2751 21970 2760
rect 22020 1630 22048 5510
rect 22388 5273 22416 7278
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 22374 5264 22430 5273
rect 22192 5228 22244 5234
rect 22374 5199 22430 5208
rect 22192 5170 22244 5176
rect 22100 4752 22152 4758
rect 22100 4694 22152 4700
rect 22112 4593 22140 4694
rect 22098 4584 22154 4593
rect 22098 4519 22154 4528
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 22008 1624 22060 1630
rect 22008 1566 22060 1572
rect 22112 800 22140 3470
rect 22204 3058 22232 5170
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22190 1320 22246 1329
rect 22190 1255 22192 1264
rect 22244 1255 22246 1264
rect 22192 1226 22244 1232
rect 22296 1086 22324 4966
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22388 3126 22416 4082
rect 22376 3120 22428 3126
rect 22376 3062 22428 3068
rect 22480 2774 22508 5510
rect 22572 2922 22600 7432
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22664 3670 22692 6938
rect 22756 4457 22784 8298
rect 22742 4448 22798 4457
rect 22742 4383 22798 4392
rect 22744 4208 22796 4214
rect 22744 4150 22796 4156
rect 22652 3664 22704 3670
rect 22652 3606 22704 3612
rect 22756 3534 22784 4150
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22848 3194 22876 11086
rect 22928 11076 22980 11082
rect 22928 11018 22980 11024
rect 22940 6769 22968 11018
rect 23032 6866 23060 12406
rect 23308 12322 23336 14758
rect 23400 14550 23428 16918
rect 23492 16250 23520 17138
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23478 16008 23534 16017
rect 23478 15943 23534 15952
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 23386 14104 23442 14113
rect 23386 14039 23388 14048
rect 23440 14039 23442 14048
rect 23388 14010 23440 14016
rect 23492 13954 23520 15943
rect 23584 14958 23612 17478
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23584 14249 23612 14418
rect 23570 14240 23626 14249
rect 23570 14175 23626 14184
rect 23676 13977 23704 19314
rect 23768 15978 23796 21626
rect 23860 21162 23888 25230
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 23860 21134 23980 21162
rect 23846 19408 23902 19417
rect 23846 19343 23902 19352
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 23860 15502 23888 19343
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23662 13968 23718 13977
rect 23492 13926 23526 13954
rect 23498 13852 23526 13926
rect 23662 13903 23718 13912
rect 23492 13824 23526 13852
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23124 12294 23336 12322
rect 23124 7426 23152 12294
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23216 11354 23244 12174
rect 23400 12102 23428 13738
rect 23492 12986 23520 13824
rect 23572 13796 23624 13802
rect 23572 13738 23624 13744
rect 23584 13297 23612 13738
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23676 13433 23704 13670
rect 23662 13424 23718 13433
rect 23662 13359 23718 13368
rect 23570 13288 23626 13297
rect 23570 13223 23626 13232
rect 23768 13172 23796 14010
rect 23860 13682 23888 14758
rect 23952 14006 23980 21134
rect 24032 21072 24084 21078
rect 24032 21014 24084 21020
rect 24044 18290 24072 21014
rect 24136 20466 24164 21286
rect 24228 20602 24256 35090
rect 24216 20596 24268 20602
rect 24216 20538 24268 20544
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24214 20224 24270 20233
rect 24214 20159 24270 20168
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24032 18148 24084 18154
rect 24032 18090 24084 18096
rect 24044 17338 24072 18090
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24032 16992 24084 16998
rect 24030 16960 24032 16969
rect 24084 16960 24086 16969
rect 24030 16895 24086 16904
rect 24030 16144 24086 16153
rect 24030 16079 24086 16088
rect 24044 16046 24072 16079
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 24030 14920 24086 14929
rect 24030 14855 24032 14864
rect 24084 14855 24086 14864
rect 24032 14826 24084 14832
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 23860 13654 23980 13682
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23860 13433 23888 13466
rect 23846 13424 23902 13433
rect 23846 13359 23902 13368
rect 23584 13144 23796 13172
rect 23584 13025 23612 13144
rect 23570 13016 23626 13025
rect 23480 12980 23532 12986
rect 23754 13016 23810 13025
rect 23570 12951 23626 12960
rect 23664 12980 23716 12986
rect 23480 12922 23532 12928
rect 23754 12951 23810 12960
rect 23664 12922 23716 12928
rect 23676 12850 23704 12922
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23478 12744 23534 12753
rect 23478 12679 23480 12688
rect 23532 12679 23534 12688
rect 23480 12650 23532 12656
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23308 11286 23336 12038
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23296 11280 23348 11286
rect 23296 11222 23348 11228
rect 23296 10736 23348 10742
rect 23296 10678 23348 10684
rect 23204 10532 23256 10538
rect 23204 10474 23256 10480
rect 23216 7750 23244 10474
rect 23308 10266 23336 10678
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 23124 7398 23244 7426
rect 23110 7304 23166 7313
rect 23110 7239 23166 7248
rect 23020 6860 23072 6866
rect 23020 6802 23072 6808
rect 22926 6760 22982 6769
rect 22926 6695 22982 6704
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 22940 5817 22968 6054
rect 23124 5914 23152 7239
rect 23216 6662 23244 7398
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 23308 6322 23336 10202
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23400 8294 23428 9454
rect 23492 8362 23520 11834
rect 23664 11620 23716 11626
rect 23664 11562 23716 11568
rect 23572 11552 23624 11558
rect 23570 11520 23572 11529
rect 23624 11520 23626 11529
rect 23570 11455 23626 11464
rect 23676 11354 23704 11562
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23768 11218 23796 12951
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23676 10810 23704 11086
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 23664 9104 23716 9110
rect 23664 9046 23716 9052
rect 23676 8906 23704 9046
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 23860 8838 23888 12786
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23768 8566 23796 8774
rect 23846 8664 23902 8673
rect 23846 8599 23902 8608
rect 23756 8560 23808 8566
rect 23756 8502 23808 8508
rect 23860 8362 23888 8599
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23848 8356 23900 8362
rect 23848 8298 23900 8304
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 22926 5808 22982 5817
rect 22926 5743 22982 5752
rect 23204 5772 23256 5778
rect 23204 5714 23256 5720
rect 23020 5636 23072 5642
rect 23020 5578 23072 5584
rect 22926 5128 22982 5137
rect 22926 5063 22928 5072
rect 22980 5063 22982 5072
rect 22928 5034 22980 5040
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 22480 2746 22600 2774
rect 22468 2304 22520 2310
rect 22468 2246 22520 2252
rect 22284 1080 22336 1086
rect 22284 1022 22336 1028
rect 22480 800 22508 2246
rect 22572 1018 22600 2746
rect 22560 1012 22612 1018
rect 22560 954 22612 960
rect 22756 800 22784 2994
rect 22940 1970 22968 3878
rect 23032 3058 23060 5578
rect 23112 4480 23164 4486
rect 23112 4422 23164 4428
rect 23124 4185 23152 4422
rect 23110 4176 23166 4185
rect 23110 4111 23166 4120
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 22928 1964 22980 1970
rect 22928 1906 22980 1912
rect 23124 800 23152 3130
rect 17868 400 17920 406
rect 17868 342 17920 348
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23216 338 23244 5714
rect 23308 3516 23336 5850
rect 23400 5098 23428 7822
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23768 7410 23796 7686
rect 23860 7585 23888 8298
rect 23846 7576 23902 7585
rect 23846 7511 23902 7520
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23952 6798 23980 13654
rect 24044 11880 24072 14350
rect 24136 12442 24164 17070
rect 24228 15638 24256 20159
rect 24320 18970 24348 37606
rect 24412 37262 24440 39200
rect 24780 37482 24808 39200
rect 24952 38004 25004 38010
rect 24952 37946 25004 37952
rect 24780 37454 24900 37482
rect 24768 37324 24820 37330
rect 24768 37266 24820 37272
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 24412 35834 24440 37198
rect 24400 35828 24452 35834
rect 24400 35770 24452 35776
rect 24674 30424 24730 30433
rect 24674 30359 24730 30368
rect 24582 25392 24638 25401
rect 24582 25327 24638 25336
rect 24398 23760 24454 23769
rect 24398 23695 24454 23704
rect 24308 18964 24360 18970
rect 24308 18906 24360 18912
rect 24306 17912 24362 17921
rect 24306 17847 24362 17856
rect 24320 15978 24348 17847
rect 24412 16250 24440 23695
rect 24492 20800 24544 20806
rect 24492 20742 24544 20748
rect 24504 20534 24532 20742
rect 24492 20528 24544 20534
rect 24490 20496 24492 20505
rect 24544 20496 24546 20505
rect 24490 20431 24546 20440
rect 24504 20405 24532 20431
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24308 15972 24360 15978
rect 24308 15914 24360 15920
rect 24398 15736 24454 15745
rect 24398 15671 24454 15680
rect 24216 15632 24268 15638
rect 24216 15574 24268 15580
rect 24412 15502 24440 15671
rect 24504 15609 24532 18566
rect 24596 16425 24624 25327
rect 24688 16726 24716 30359
rect 24780 20874 24808 37266
rect 24872 36922 24900 37454
rect 24860 36916 24912 36922
rect 24860 36858 24912 36864
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 24780 19145 24808 19654
rect 24766 19136 24822 19145
rect 24766 19071 24822 19080
rect 24768 18760 24820 18766
rect 24872 18737 24900 20198
rect 24964 19854 24992 37946
rect 25148 36378 25176 39200
rect 25320 37732 25372 37738
rect 25320 37674 25372 37680
rect 25228 36780 25280 36786
rect 25228 36722 25280 36728
rect 25136 36372 25188 36378
rect 25136 36314 25188 36320
rect 25044 36168 25096 36174
rect 25044 36110 25096 36116
rect 25056 34950 25084 36110
rect 25240 35494 25268 36722
rect 25228 35488 25280 35494
rect 25228 35430 25280 35436
rect 25044 34944 25096 34950
rect 25044 34886 25096 34892
rect 25056 28937 25084 34886
rect 25240 34610 25268 35430
rect 25228 34604 25280 34610
rect 25228 34546 25280 34552
rect 25042 28928 25098 28937
rect 25042 28863 25098 28872
rect 25228 26920 25280 26926
rect 25228 26862 25280 26868
rect 25136 25764 25188 25770
rect 25136 25706 25188 25712
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 25056 19553 25084 19722
rect 25042 19544 25098 19553
rect 25042 19479 25098 19488
rect 24950 19000 25006 19009
rect 24950 18935 24952 18944
rect 25004 18935 25006 18944
rect 24952 18906 25004 18912
rect 24950 18864 25006 18873
rect 24950 18799 25006 18808
rect 24768 18702 24820 18708
rect 24858 18728 24914 18737
rect 24780 18426 24808 18702
rect 24858 18663 24914 18672
rect 24964 18426 24992 18799
rect 24768 18420 24820 18426
rect 24768 18362 24820 18368
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24780 17513 24808 18226
rect 25148 18034 25176 25706
rect 24872 18006 25176 18034
rect 24766 17504 24822 17513
rect 24766 17439 24822 17448
rect 24780 17134 24808 17439
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24582 16416 24638 16425
rect 24582 16351 24638 16360
rect 24596 15638 24624 16351
rect 24872 15978 24900 18006
rect 25240 17954 25268 26862
rect 25332 21146 25360 37674
rect 25608 37262 25636 39200
rect 25596 37256 25648 37262
rect 25596 37198 25648 37204
rect 25608 36378 25636 37198
rect 25976 36922 26004 39200
rect 25964 36916 26016 36922
rect 25964 36858 26016 36864
rect 26056 36780 26108 36786
rect 26056 36722 26108 36728
rect 25596 36372 25648 36378
rect 25596 36314 25648 36320
rect 25596 35556 25648 35562
rect 25596 35498 25648 35504
rect 25502 23216 25558 23225
rect 25502 23151 25558 23160
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25332 20534 25360 21082
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 25516 19394 25544 23151
rect 25608 20058 25636 35498
rect 26068 35494 26096 36722
rect 26436 36378 26464 39200
rect 26804 37262 26832 39200
rect 26884 37324 26936 37330
rect 26884 37266 26936 37272
rect 26792 37256 26844 37262
rect 26792 37198 26844 37204
rect 26424 36372 26476 36378
rect 26424 36314 26476 36320
rect 26516 36168 26568 36174
rect 26516 36110 26568 36116
rect 26332 35624 26384 35630
rect 26332 35566 26384 35572
rect 26056 35488 26108 35494
rect 26056 35430 26108 35436
rect 26068 35018 26096 35430
rect 26344 35290 26372 35566
rect 26528 35290 26556 36110
rect 26332 35284 26384 35290
rect 26332 35226 26384 35232
rect 26516 35284 26568 35290
rect 26516 35226 26568 35232
rect 26240 35216 26292 35222
rect 26240 35158 26292 35164
rect 26056 35012 26108 35018
rect 26056 34954 26108 34960
rect 25780 34740 25832 34746
rect 25780 34682 25832 34688
rect 25688 20868 25740 20874
rect 25688 20810 25740 20816
rect 25596 20052 25648 20058
rect 25596 19994 25648 20000
rect 25516 19366 25636 19394
rect 25504 19304 25556 19310
rect 25502 19272 25504 19281
rect 25556 19272 25558 19281
rect 25502 19207 25558 19216
rect 25502 18320 25558 18329
rect 25320 18284 25372 18290
rect 25502 18255 25558 18264
rect 25320 18226 25372 18232
rect 25332 18086 25360 18226
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25056 17926 25268 17954
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24964 16114 24992 17478
rect 25056 16658 25084 17926
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 25056 16250 25084 16594
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24860 15972 24912 15978
rect 24860 15914 24912 15920
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 24584 15632 24636 15638
rect 24490 15600 24546 15609
rect 24584 15574 24636 15580
rect 24490 15535 24546 15544
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24214 15192 24270 15201
rect 24214 15127 24270 15136
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24124 11892 24176 11898
rect 24044 11852 24124 11880
rect 24124 11834 24176 11840
rect 24228 11150 24256 15127
rect 24400 14952 24452 14958
rect 24400 14894 24452 14900
rect 24308 13932 24360 13938
rect 24308 13874 24360 13880
rect 24320 13190 24348 13874
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24320 12714 24348 13126
rect 24308 12708 24360 12714
rect 24308 12650 24360 12656
rect 24412 12594 24440 14894
rect 24504 13326 24532 15535
rect 24688 15162 24716 15846
rect 24964 15706 24992 16050
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 24676 14884 24728 14890
rect 24952 14884 25004 14890
rect 24728 14844 24808 14872
rect 24676 14826 24728 14832
rect 24584 14816 24636 14822
rect 24584 14758 24636 14764
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24492 12912 24544 12918
rect 24492 12854 24544 12860
rect 24320 12566 24440 12594
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 24136 10470 24164 11018
rect 24320 11014 24348 12566
rect 24504 12170 24532 12854
rect 24400 12164 24452 12170
rect 24400 12106 24452 12112
rect 24492 12164 24544 12170
rect 24492 12106 24544 12112
rect 24412 11529 24440 12106
rect 24492 11756 24544 11762
rect 24492 11698 24544 11704
rect 24504 11558 24532 11698
rect 24492 11552 24544 11558
rect 24398 11520 24454 11529
rect 24492 11494 24544 11500
rect 24398 11455 24454 11464
rect 24398 11384 24454 11393
rect 24398 11319 24400 11328
rect 24452 11319 24454 11328
rect 24400 11290 24452 11296
rect 24504 11234 24532 11494
rect 24412 11206 24532 11234
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24124 10464 24176 10470
rect 24124 10406 24176 10412
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 23940 6792 23992 6798
rect 23846 6760 23902 6769
rect 23940 6734 23992 6740
rect 23846 6695 23902 6704
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23388 5092 23440 5098
rect 23388 5034 23440 5040
rect 23388 3528 23440 3534
rect 23308 3488 23388 3516
rect 23308 3194 23336 3488
rect 23388 3470 23440 3476
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23492 2446 23520 6598
rect 23572 6384 23624 6390
rect 23570 6352 23572 6361
rect 23624 6352 23626 6361
rect 23570 6287 23626 6296
rect 23664 5568 23716 5574
rect 23664 5510 23716 5516
rect 23676 5370 23704 5510
rect 23664 5364 23716 5370
rect 23664 5306 23716 5312
rect 23662 4992 23718 5001
rect 23662 4927 23718 4936
rect 23676 4826 23704 4927
rect 23664 4820 23716 4826
rect 23664 4762 23716 4768
rect 23570 4720 23626 4729
rect 23570 4655 23572 4664
rect 23624 4655 23626 4664
rect 23572 4626 23624 4632
rect 23572 3596 23624 3602
rect 23572 3538 23624 3544
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23388 2304 23440 2310
rect 23388 2246 23440 2252
rect 23400 800 23428 2246
rect 23584 950 23612 3538
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 23572 944 23624 950
rect 23572 886 23624 892
rect 23676 800 23704 2994
rect 23768 2446 23796 6598
rect 23860 3194 23888 6695
rect 24044 6390 24072 9862
rect 24136 9042 24164 10406
rect 24308 9920 24360 9926
rect 24308 9862 24360 9868
rect 24216 9648 24268 9654
rect 24214 9616 24216 9625
rect 24268 9616 24270 9625
rect 24214 9551 24270 9560
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 24216 8832 24268 8838
rect 24216 8774 24268 8780
rect 24124 7336 24176 7342
rect 24124 7278 24176 7284
rect 24032 6384 24084 6390
rect 24032 6326 24084 6332
rect 23940 5160 23992 5166
rect 23940 5102 23992 5108
rect 23952 4026 23980 5102
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 24044 4185 24072 4966
rect 24136 4554 24164 7278
rect 24124 4548 24176 4554
rect 24124 4490 24176 4496
rect 24030 4176 24086 4185
rect 24030 4111 24086 4120
rect 23952 3998 24072 4026
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23952 1698 23980 3878
rect 24044 3534 24072 3998
rect 24124 4004 24176 4010
rect 24124 3946 24176 3952
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 23940 1692 23992 1698
rect 23940 1634 23992 1640
rect 24044 800 24072 3470
rect 24136 1222 24164 3946
rect 24228 3194 24256 8774
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24320 2446 24348 9862
rect 24412 8786 24440 11206
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24504 8945 24532 9114
rect 24490 8936 24546 8945
rect 24490 8871 24546 8880
rect 24412 8758 24532 8786
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24308 2440 24360 2446
rect 24308 2382 24360 2388
rect 24308 2304 24360 2310
rect 24308 2246 24360 2252
rect 24124 1216 24176 1222
rect 24124 1158 24176 1164
rect 24320 800 24348 2246
rect 24412 1193 24440 7686
rect 24504 6866 24532 8758
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24596 6798 24624 14758
rect 24674 14512 24730 14521
rect 24674 14447 24730 14456
rect 24688 14414 24716 14447
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24688 14074 24716 14350
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24780 13394 24808 14844
rect 24952 14826 25004 14832
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24780 11336 24808 12922
rect 24872 12646 24900 14350
rect 24964 14346 24992 14826
rect 24952 14340 25004 14346
rect 24952 14282 25004 14288
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 25056 12322 25084 14962
rect 24964 12294 25084 12322
rect 24780 11308 24900 11336
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24688 10606 24716 10950
rect 24780 10810 24808 11154
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24676 10600 24728 10606
rect 24674 10568 24676 10577
rect 24728 10568 24730 10577
rect 24674 10503 24730 10512
rect 24872 10266 24900 11308
rect 24964 10441 24992 12294
rect 24950 10432 25006 10441
rect 24950 10367 25006 10376
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 24872 9994 24900 10202
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24858 9480 24914 9489
rect 24858 9415 24914 9424
rect 24872 8809 24900 9415
rect 25042 9344 25098 9353
rect 25042 9279 25098 9288
rect 25056 8838 25084 9279
rect 25044 8832 25096 8838
rect 24858 8800 24914 8809
rect 24858 8735 24914 8744
rect 25042 8800 25044 8809
rect 25096 8800 25098 8809
rect 25042 8735 25098 8744
rect 25042 8256 25098 8265
rect 25042 8191 25098 8200
rect 25056 8090 25084 8191
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 25148 7954 25176 17682
rect 25412 16992 25464 16998
rect 25412 16934 25464 16940
rect 25228 16516 25280 16522
rect 25228 16458 25280 16464
rect 25240 15201 25268 16458
rect 25318 16280 25374 16289
rect 25318 16215 25320 16224
rect 25372 16215 25374 16224
rect 25320 16186 25372 16192
rect 25318 15464 25374 15473
rect 25318 15399 25374 15408
rect 25226 15192 25282 15201
rect 25226 15127 25282 15136
rect 25332 14006 25360 15399
rect 25320 14000 25372 14006
rect 25320 13942 25372 13948
rect 25228 13728 25280 13734
rect 25228 13670 25280 13676
rect 25240 12782 25268 13670
rect 25332 13530 25360 13942
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25318 13288 25374 13297
rect 25318 13223 25374 13232
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 25240 11937 25268 12242
rect 25226 11928 25282 11937
rect 25332 11898 25360 13223
rect 25226 11863 25282 11872
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25240 10713 25268 11494
rect 25226 10704 25282 10713
rect 25226 10639 25282 10648
rect 25240 10441 25268 10639
rect 25226 10432 25282 10441
rect 25226 10367 25282 10376
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25240 9353 25268 9658
rect 25226 9344 25282 9353
rect 25226 9279 25282 9288
rect 25424 8022 25452 16934
rect 25516 16726 25544 18255
rect 25504 16720 25556 16726
rect 25504 16662 25556 16668
rect 25502 15192 25558 15201
rect 25608 15162 25636 19366
rect 25700 17882 25728 20810
rect 25792 20602 25820 34682
rect 26252 34542 26280 35158
rect 26528 35086 26556 35226
rect 26516 35080 26568 35086
rect 26516 35022 26568 35028
rect 26240 34536 26292 34542
rect 26240 34478 26292 34484
rect 26608 27328 26660 27334
rect 26608 27270 26660 27276
rect 26332 24948 26384 24954
rect 26332 24890 26384 24896
rect 26240 22500 26292 22506
rect 26240 22442 26292 22448
rect 26148 22160 26200 22166
rect 26148 22102 26200 22108
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25688 15428 25740 15434
rect 25688 15370 25740 15376
rect 25502 15127 25558 15136
rect 25596 15156 25648 15162
rect 25516 15094 25544 15127
rect 25596 15098 25648 15104
rect 25504 15088 25556 15094
rect 25504 15030 25556 15036
rect 25516 13530 25544 15030
rect 25700 14006 25728 15370
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 25516 13410 25544 13466
rect 25516 13382 25636 13410
rect 25608 12434 25636 13382
rect 25516 12406 25636 12434
rect 25686 12472 25742 12481
rect 25686 12407 25688 12416
rect 25516 10742 25544 12406
rect 25740 12407 25742 12416
rect 25688 12378 25740 12384
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25700 10985 25728 11018
rect 25686 10976 25742 10985
rect 25686 10911 25742 10920
rect 25504 10736 25556 10742
rect 25504 10678 25556 10684
rect 25596 10600 25648 10606
rect 25596 10542 25648 10548
rect 25504 10192 25556 10198
rect 25504 10134 25556 10140
rect 25516 9994 25544 10134
rect 25608 10062 25636 10542
rect 25792 10282 25820 20402
rect 25870 19408 25926 19417
rect 25870 19343 25926 19352
rect 25884 16794 25912 19343
rect 25872 16788 25924 16794
rect 25872 16730 25924 16736
rect 25872 15632 25924 15638
rect 25872 15574 25924 15580
rect 25884 12889 25912 15574
rect 25976 13734 26004 20878
rect 26054 19408 26110 19417
rect 26054 19343 26110 19352
rect 26068 17882 26096 19343
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 26068 17066 26096 17818
rect 26056 17060 26108 17066
rect 26056 17002 26108 17008
rect 26160 15881 26188 22102
rect 26146 15872 26202 15881
rect 26146 15807 26202 15816
rect 26160 15706 26188 15807
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26056 15632 26108 15638
rect 26056 15574 26108 15580
rect 26068 15337 26096 15574
rect 26054 15328 26110 15337
rect 26054 15263 26110 15272
rect 26068 14618 26096 15263
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 26160 13938 26188 15642
rect 26148 13932 26200 13938
rect 26148 13874 26200 13880
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 26068 13297 26096 13330
rect 26054 13288 26110 13297
rect 26054 13223 26110 13232
rect 26148 13252 26200 13258
rect 26148 13194 26200 13200
rect 25962 13152 26018 13161
rect 25962 13087 26018 13096
rect 25976 12986 26004 13087
rect 26160 12986 26188 13194
rect 25964 12980 26016 12986
rect 25964 12922 26016 12928
rect 26148 12980 26200 12986
rect 26148 12922 26200 12928
rect 25870 12880 25926 12889
rect 25870 12815 25926 12824
rect 26160 12442 26188 12922
rect 26148 12436 26200 12442
rect 26148 12378 26200 12384
rect 26252 12345 26280 22442
rect 26344 18222 26372 24890
rect 26620 21146 26648 27270
rect 26790 24712 26846 24721
rect 26790 24647 26846 24656
rect 26608 21140 26660 21146
rect 26608 21082 26660 21088
rect 26620 19334 26648 21082
rect 26528 19306 26648 19334
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26332 18216 26384 18222
rect 26332 18158 26384 18164
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26330 16280 26386 16289
rect 26330 16215 26386 16224
rect 26344 16182 26372 16215
rect 26332 16176 26384 16182
rect 26332 16118 26384 16124
rect 26344 16017 26372 16118
rect 26330 16008 26386 16017
rect 26330 15943 26386 15952
rect 26330 15736 26386 15745
rect 26330 15671 26332 15680
rect 26384 15671 26386 15680
rect 26332 15642 26384 15648
rect 26436 15570 26464 16390
rect 26332 15564 26384 15570
rect 26332 15506 26384 15512
rect 26424 15564 26476 15570
rect 26424 15506 26476 15512
rect 26344 15162 26372 15506
rect 26436 15162 26464 15506
rect 26332 15156 26384 15162
rect 26332 15098 26384 15104
rect 26424 15156 26476 15162
rect 26424 15098 26476 15104
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 26344 13326 26372 14214
rect 26332 13320 26384 13326
rect 26332 13262 26384 13268
rect 26238 12336 26294 12345
rect 26238 12271 26294 12280
rect 26238 11248 26294 11257
rect 26238 11183 26294 11192
rect 26252 11082 26280 11183
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 25700 10254 25820 10282
rect 25700 10169 25728 10254
rect 25780 10192 25832 10198
rect 25686 10160 25742 10169
rect 25780 10134 25832 10140
rect 25686 10095 25742 10104
rect 25596 10056 25648 10062
rect 25596 9998 25648 10004
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 25502 9888 25558 9897
rect 25502 9823 25558 9832
rect 25516 8634 25544 9823
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25594 8120 25650 8129
rect 25594 8055 25596 8064
rect 25648 8055 25650 8064
rect 25596 8026 25648 8032
rect 25412 8016 25464 8022
rect 25412 7958 25464 7964
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24492 6180 24544 6186
rect 24492 6122 24544 6128
rect 24504 1834 24532 6122
rect 24584 6112 24636 6118
rect 24584 6054 24636 6060
rect 24596 5710 24624 6054
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24584 3936 24636 3942
rect 24584 3878 24636 3884
rect 24596 3505 24624 3878
rect 24582 3496 24638 3505
rect 24582 3431 24638 3440
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24596 2990 24624 3334
rect 24688 2990 24716 4966
rect 24584 2984 24636 2990
rect 24584 2926 24636 2932
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 24492 1828 24544 1834
rect 24492 1770 24544 1776
rect 24398 1184 24454 1193
rect 24398 1119 24454 1128
rect 24688 800 24716 2926
rect 24780 882 24808 7142
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 24872 3398 24900 5510
rect 24952 4480 25004 4486
rect 24952 4422 25004 4428
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 24964 4185 24992 4422
rect 24950 4176 25006 4185
rect 24950 4111 25006 4120
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24768 876 24820 882
rect 24768 818 24820 824
rect 24964 800 24992 3470
rect 25056 3126 25084 4422
rect 25148 4214 25176 6598
rect 25136 4208 25188 4214
rect 25136 4150 25188 4156
rect 25136 3936 25188 3942
rect 25134 3904 25136 3913
rect 25188 3904 25190 3913
rect 25134 3839 25190 3848
rect 25240 3534 25268 6598
rect 25412 6112 25464 6118
rect 25412 6054 25464 6060
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25044 3120 25096 3126
rect 25044 3062 25096 3068
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25148 1902 25176 2246
rect 25136 1896 25188 1902
rect 25136 1838 25188 1844
rect 25240 800 25268 2790
rect 23204 332 23256 338
rect 23204 274 23256 280
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 24030 0 24086 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25332 66 25360 3878
rect 25424 1154 25452 6054
rect 25596 5024 25648 5030
rect 25596 4966 25648 4972
rect 25608 2530 25636 4966
rect 25700 3602 25728 6054
rect 25688 3596 25740 3602
rect 25688 3538 25740 3544
rect 25688 3392 25740 3398
rect 25688 3334 25740 3340
rect 25516 2502 25636 2530
rect 25412 1148 25464 1154
rect 25412 1090 25464 1096
rect 25516 202 25544 2502
rect 25596 2440 25648 2446
rect 25596 2382 25648 2388
rect 25608 800 25636 2382
rect 25700 2038 25728 3334
rect 25792 3058 25820 10134
rect 26252 10033 26280 11018
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26238 10024 26294 10033
rect 26238 9959 26294 9968
rect 25964 9648 26016 9654
rect 25962 9616 25964 9625
rect 26016 9616 26018 9625
rect 25962 9551 26018 9560
rect 25976 9178 26004 9551
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 26344 8498 26372 10406
rect 26436 9178 26464 14962
rect 26528 12918 26556 19306
rect 26608 18624 26660 18630
rect 26606 18592 26608 18601
rect 26660 18592 26662 18601
rect 26606 18527 26662 18536
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26516 12912 26568 12918
rect 26516 12854 26568 12860
rect 26620 12764 26648 15846
rect 26712 15026 26740 19314
rect 26804 16250 26832 24647
rect 26896 20874 26924 37266
rect 27172 36922 27200 39200
rect 27436 37868 27488 37874
rect 27436 37810 27488 37816
rect 27448 37466 27476 37810
rect 27436 37460 27488 37466
rect 27436 37402 27488 37408
rect 27528 37256 27580 37262
rect 27528 37198 27580 37204
rect 27540 36922 27568 37198
rect 27160 36916 27212 36922
rect 27160 36858 27212 36864
rect 27528 36916 27580 36922
rect 27528 36858 27580 36864
rect 27068 36780 27120 36786
rect 27068 36722 27120 36728
rect 27080 35494 27108 36722
rect 27632 36378 27660 39200
rect 27712 37868 27764 37874
rect 27712 37810 27764 37816
rect 27620 36372 27672 36378
rect 27620 36314 27672 36320
rect 27620 36168 27672 36174
rect 27620 36110 27672 36116
rect 27632 35562 27660 36110
rect 27620 35556 27672 35562
rect 27620 35498 27672 35504
rect 27068 35488 27120 35494
rect 27068 35430 27120 35436
rect 26976 24744 27028 24750
rect 26976 24686 27028 24692
rect 26884 20868 26936 20874
rect 26884 20810 26936 20816
rect 26884 19780 26936 19786
rect 26884 19722 26936 19728
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26804 15706 26832 16186
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 26700 15020 26752 15026
rect 26700 14962 26752 14968
rect 26792 14340 26844 14346
rect 26792 14282 26844 14288
rect 26700 13252 26752 13258
rect 26700 13194 26752 13200
rect 26528 12736 26648 12764
rect 26424 9172 26476 9178
rect 26424 9114 26476 9120
rect 26332 8492 26384 8498
rect 26332 8434 26384 8440
rect 25964 8424 26016 8430
rect 25962 8392 25964 8401
rect 26016 8392 26018 8401
rect 25962 8327 26018 8336
rect 26146 7168 26202 7177
rect 26146 7103 26202 7112
rect 26160 5574 26188 7103
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 26148 5568 26200 5574
rect 26148 5510 26200 5516
rect 26252 3516 26280 6054
rect 26332 5024 26384 5030
rect 26332 4966 26384 4972
rect 26160 3488 26280 3516
rect 26160 3126 26188 3488
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 25872 3120 25924 3126
rect 25872 3062 25924 3068
rect 26148 3120 26200 3126
rect 26148 3062 26200 3068
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 25792 2446 25820 2790
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 25688 2032 25740 2038
rect 25688 1974 25740 1980
rect 25884 800 25912 3062
rect 25962 2544 26018 2553
rect 25962 2479 25964 2488
rect 26016 2479 26018 2488
rect 25964 2450 26016 2456
rect 26252 800 26280 3334
rect 25504 196 25556 202
rect 25504 138 25556 144
rect 25320 60 25372 66
rect 25320 2 25372 8
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26238 0 26294 800
rect 26344 270 26372 4966
rect 26424 4480 26476 4486
rect 26424 4422 26476 4428
rect 26436 2854 26464 4422
rect 26424 2848 26476 2854
rect 26424 2790 26476 2796
rect 26528 2496 26556 12736
rect 26712 12102 26740 13194
rect 26700 12096 26752 12102
rect 26700 12038 26752 12044
rect 26712 10810 26740 12038
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 26804 10690 26832 14282
rect 26620 10662 26832 10690
rect 26620 5302 26648 10662
rect 26792 9988 26844 9994
rect 26792 9930 26844 9936
rect 26700 9580 26752 9586
rect 26700 9522 26752 9528
rect 26608 5296 26660 5302
rect 26608 5238 26660 5244
rect 26608 4480 26660 4486
rect 26608 4422 26660 4428
rect 26436 2468 26556 2496
rect 26436 1873 26464 2468
rect 26516 2372 26568 2378
rect 26516 2314 26568 2320
rect 26422 1864 26478 1873
rect 26422 1799 26478 1808
rect 26528 800 26556 2314
rect 26332 264 26384 270
rect 26332 206 26384 212
rect 26514 0 26570 800
rect 26620 134 26648 4422
rect 26712 3058 26740 9522
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 26804 2990 26832 9930
rect 26896 8362 26924 19722
rect 26988 19417 27016 24686
rect 27080 23322 27108 35430
rect 27632 35329 27660 35498
rect 27618 35320 27674 35329
rect 27618 35255 27674 35264
rect 27252 34536 27304 34542
rect 27252 34478 27304 34484
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 27068 23316 27120 23322
rect 27068 23258 27120 23264
rect 27172 19990 27200 24074
rect 27264 20466 27292 34478
rect 27526 25664 27582 25673
rect 27526 25599 27582 25608
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 27160 19984 27212 19990
rect 27160 19926 27212 19932
rect 27160 19712 27212 19718
rect 27160 19654 27212 19660
rect 26974 19408 27030 19417
rect 26974 19343 27030 19352
rect 26976 18692 27028 18698
rect 26976 18634 27028 18640
rect 26988 16998 27016 18634
rect 27068 18080 27120 18086
rect 27068 18022 27120 18028
rect 27080 17678 27108 18022
rect 27068 17672 27120 17678
rect 27068 17614 27120 17620
rect 26976 16992 27028 16998
rect 26976 16934 27028 16940
rect 26988 16232 27016 16934
rect 27066 16824 27122 16833
rect 27066 16759 27122 16768
rect 27080 16726 27108 16759
rect 27068 16720 27120 16726
rect 27068 16662 27120 16668
rect 26988 16204 27108 16232
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 26988 15706 27016 16050
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 26974 14784 27030 14793
rect 26974 14719 27030 14728
rect 26988 14618 27016 14719
rect 26976 14612 27028 14618
rect 26976 14554 27028 14560
rect 27080 14550 27108 16204
rect 27068 14544 27120 14550
rect 27068 14486 27120 14492
rect 26976 13864 27028 13870
rect 26976 13806 27028 13812
rect 26988 12442 27016 13806
rect 27080 12646 27108 14486
rect 27068 12640 27120 12646
rect 27068 12582 27120 12588
rect 26976 12436 27028 12442
rect 26976 12378 27028 12384
rect 26976 11552 27028 11558
rect 26976 11494 27028 11500
rect 26988 10674 27016 11494
rect 26976 10668 27028 10674
rect 26976 10610 27028 10616
rect 26988 9466 27016 10610
rect 27172 10169 27200 19654
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27250 19272 27306 19281
rect 27250 19207 27306 19216
rect 27264 18970 27292 19207
rect 27252 18964 27304 18970
rect 27252 18906 27304 18912
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 27264 18086 27292 18226
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 27252 17672 27304 17678
rect 27252 17614 27304 17620
rect 27264 15094 27292 17614
rect 27252 15088 27304 15094
rect 27252 15030 27304 15036
rect 27252 12640 27304 12646
rect 27252 12582 27304 12588
rect 27264 11354 27292 12582
rect 27252 11348 27304 11354
rect 27252 11290 27304 11296
rect 27158 10160 27214 10169
rect 27158 10095 27214 10104
rect 27252 10124 27304 10130
rect 27252 10066 27304 10072
rect 27264 9722 27292 10066
rect 27252 9716 27304 9722
rect 27252 9658 27304 9664
rect 27356 9518 27384 19314
rect 27448 18426 27476 20198
rect 27436 18420 27488 18426
rect 27436 18362 27488 18368
rect 27540 17241 27568 25599
rect 27724 21690 27752 37810
rect 28000 37262 28028 39200
rect 28172 37936 28224 37942
rect 28172 37878 28224 37884
rect 28184 37466 28212 37878
rect 28172 37460 28224 37466
rect 28172 37402 28224 37408
rect 27988 37256 28040 37262
rect 27988 37198 28040 37204
rect 28460 36922 28488 39200
rect 28448 36916 28500 36922
rect 28448 36858 28500 36864
rect 28540 36780 28592 36786
rect 28540 36722 28592 36728
rect 28552 36378 28580 36722
rect 28540 36372 28592 36378
rect 28540 36314 28592 36320
rect 28552 33114 28580 36314
rect 28828 35834 28856 39200
rect 29196 37262 29224 39200
rect 29184 37256 29236 37262
rect 29184 37198 29236 37204
rect 29656 36922 29684 39200
rect 30024 39114 30052 39200
rect 30116 39114 30144 39222
rect 30024 39086 30144 39114
rect 30012 38072 30064 38078
rect 30012 38014 30064 38020
rect 29828 37800 29880 37806
rect 29828 37742 29880 37748
rect 29736 37392 29788 37398
rect 29736 37334 29788 37340
rect 29644 36916 29696 36922
rect 29644 36858 29696 36864
rect 29552 36780 29604 36786
rect 29552 36722 29604 36728
rect 28816 35828 28868 35834
rect 28816 35770 28868 35776
rect 28724 35760 28776 35766
rect 28724 35702 28776 35708
rect 28540 33108 28592 33114
rect 28540 33050 28592 33056
rect 28080 29640 28132 29646
rect 28080 29582 28132 29588
rect 27894 25936 27950 25945
rect 27894 25871 27950 25880
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27724 20534 27752 21626
rect 27804 21412 27856 21418
rect 27804 21354 27856 21360
rect 27712 20528 27764 20534
rect 27712 20470 27764 20476
rect 27618 19816 27674 19825
rect 27618 19751 27620 19760
rect 27672 19751 27674 19760
rect 27620 19722 27672 19728
rect 27620 19236 27672 19242
rect 27620 19178 27672 19184
rect 27632 18970 27660 19178
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 27526 17232 27582 17241
rect 27526 17167 27582 17176
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27632 16250 27660 16730
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27436 15632 27488 15638
rect 27436 15574 27488 15580
rect 27448 15366 27476 15574
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 27448 14657 27476 14758
rect 27434 14648 27490 14657
rect 27434 14583 27436 14592
rect 27488 14583 27490 14592
rect 27436 14554 27488 14560
rect 27448 14249 27476 14554
rect 27540 14385 27568 15302
rect 27632 14618 27660 16186
rect 27710 15056 27766 15065
rect 27710 14991 27712 15000
rect 27764 14991 27766 15000
rect 27712 14962 27764 14968
rect 27816 14906 27844 21354
rect 27908 17882 27936 25871
rect 28092 21146 28120 29582
rect 28262 25800 28318 25809
rect 28262 25735 28318 25744
rect 28080 21140 28132 21146
rect 28080 21082 28132 21088
rect 28172 20052 28224 20058
rect 28172 19994 28224 20000
rect 28184 19174 28212 19994
rect 28172 19168 28224 19174
rect 28172 19110 28224 19116
rect 28080 18420 28132 18426
rect 28080 18362 28132 18368
rect 27896 17876 27948 17882
rect 27896 17818 27948 17824
rect 27908 17202 27936 17818
rect 27986 17232 28042 17241
rect 27896 17196 27948 17202
rect 27986 17167 28042 17176
rect 27896 17138 27948 17144
rect 27724 14878 27844 14906
rect 27620 14612 27672 14618
rect 27620 14554 27672 14560
rect 27526 14376 27582 14385
rect 27526 14311 27582 14320
rect 27434 14240 27490 14249
rect 27434 14175 27490 14184
rect 27540 14006 27568 14311
rect 27528 14000 27580 14006
rect 27528 13942 27580 13948
rect 27632 13530 27660 14554
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27528 13184 27580 13190
rect 27528 13126 27580 13132
rect 27436 12096 27488 12102
rect 27434 12064 27436 12073
rect 27488 12064 27490 12073
rect 27434 11999 27490 12008
rect 27540 11898 27568 13126
rect 27620 12912 27672 12918
rect 27620 12854 27672 12860
rect 27528 11892 27580 11898
rect 27528 11834 27580 11840
rect 27632 11830 27660 12854
rect 27620 11824 27672 11830
rect 27620 11766 27672 11772
rect 27724 10849 27752 14878
rect 27804 14816 27856 14822
rect 27804 14758 27856 14764
rect 27816 12918 27844 14758
rect 27896 14272 27948 14278
rect 27896 14214 27948 14220
rect 27908 13394 27936 14214
rect 27896 13388 27948 13394
rect 27896 13330 27948 13336
rect 27894 13288 27950 13297
rect 27894 13223 27950 13232
rect 27804 12912 27856 12918
rect 27804 12854 27856 12860
rect 27804 12232 27856 12238
rect 27804 12174 27856 12180
rect 27816 11898 27844 12174
rect 27804 11892 27856 11898
rect 27804 11834 27856 11840
rect 27710 10840 27766 10849
rect 27710 10775 27766 10784
rect 27908 10062 27936 13223
rect 28000 12306 28028 17167
rect 27988 12300 28040 12306
rect 27988 12242 28040 12248
rect 27986 11792 28042 11801
rect 27986 11727 27988 11736
rect 28040 11727 28042 11736
rect 27988 11698 28040 11704
rect 27896 10056 27948 10062
rect 27896 9998 27948 10004
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 27344 9512 27396 9518
rect 26988 9438 27200 9466
rect 27344 9454 27396 9460
rect 27068 9376 27120 9382
rect 27068 9318 27120 9324
rect 27080 9178 27108 9318
rect 26976 9172 27028 9178
rect 26976 9114 27028 9120
rect 27068 9172 27120 9178
rect 27068 9114 27120 9120
rect 26988 8906 27016 9114
rect 26976 8900 27028 8906
rect 26976 8842 27028 8848
rect 26884 8356 26936 8362
rect 26884 8298 26936 8304
rect 27172 8294 27200 9438
rect 27436 9036 27488 9042
rect 27436 8978 27488 8984
rect 27080 8266 27200 8294
rect 26882 6896 26938 6905
rect 26882 6831 26938 6840
rect 26896 6497 26924 6831
rect 26882 6488 26938 6497
rect 26882 6423 26938 6432
rect 26976 5024 27028 5030
rect 26976 4966 27028 4972
rect 26988 4622 27016 4966
rect 26976 4616 27028 4622
rect 26976 4558 27028 4564
rect 27080 4434 27108 8266
rect 27158 5944 27214 5953
rect 27158 5879 27160 5888
rect 27212 5879 27214 5888
rect 27160 5850 27212 5856
rect 27342 5128 27398 5137
rect 27342 5063 27398 5072
rect 26988 4406 27108 4434
rect 27252 4480 27304 4486
rect 27252 4422 27304 4428
rect 26884 3188 26936 3194
rect 26884 3130 26936 3136
rect 26792 2984 26844 2990
rect 26792 2926 26844 2932
rect 26896 800 26924 3130
rect 26988 2774 27016 4406
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 27068 3460 27120 3466
rect 27068 3402 27120 3408
rect 27080 3194 27108 3402
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 26988 2746 27108 2774
rect 27080 1970 27108 2746
rect 27068 1964 27120 1970
rect 27068 1906 27120 1912
rect 27172 800 27200 3878
rect 27264 2378 27292 4422
rect 27356 3670 27384 5063
rect 27448 3670 27476 8978
rect 27528 3732 27580 3738
rect 27528 3674 27580 3680
rect 27344 3664 27396 3670
rect 27344 3606 27396 3612
rect 27436 3664 27488 3670
rect 27436 3606 27488 3612
rect 27344 3460 27396 3466
rect 27344 3402 27396 3408
rect 27356 3126 27384 3402
rect 27540 3194 27568 3674
rect 27632 3534 27660 9862
rect 27908 9722 27936 9998
rect 27988 9920 28040 9926
rect 27988 9862 28040 9868
rect 27896 9716 27948 9722
rect 27896 9658 27948 9664
rect 27712 8832 27764 8838
rect 27712 8774 27764 8780
rect 27724 8634 27752 8774
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27896 6724 27948 6730
rect 27896 6666 27948 6672
rect 27802 5944 27858 5953
rect 27908 5914 27936 6666
rect 27802 5879 27804 5888
rect 27856 5879 27858 5888
rect 27896 5908 27948 5914
rect 27804 5850 27856 5856
rect 27896 5850 27948 5856
rect 27712 4480 27764 4486
rect 27712 4422 27764 4428
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 27724 3126 27752 4422
rect 27816 4026 27844 5850
rect 27896 5092 27948 5098
rect 27896 5034 27948 5040
rect 27908 4554 27936 5034
rect 27896 4548 27948 4554
rect 27896 4490 27948 4496
rect 28000 4146 28028 9862
rect 28092 5370 28120 18362
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28184 18193 28212 18226
rect 28170 18184 28226 18193
rect 28170 18119 28226 18128
rect 28276 18034 28304 25735
rect 28540 23860 28592 23866
rect 28540 23802 28592 23808
rect 28448 23316 28500 23322
rect 28448 23258 28500 23264
rect 28354 20632 28410 20641
rect 28354 20567 28356 20576
rect 28408 20567 28410 20576
rect 28356 20538 28408 20544
rect 28368 19854 28396 20538
rect 28460 19990 28488 23258
rect 28448 19984 28500 19990
rect 28448 19926 28500 19932
rect 28356 19848 28408 19854
rect 28356 19790 28408 19796
rect 28448 19780 28500 19786
rect 28448 19722 28500 19728
rect 28460 19514 28488 19722
rect 28448 19508 28500 19514
rect 28448 19450 28500 19456
rect 28446 19136 28502 19145
rect 28446 19071 28502 19080
rect 28356 18216 28408 18222
rect 28356 18158 28408 18164
rect 28184 18006 28304 18034
rect 28184 12986 28212 18006
rect 28262 17912 28318 17921
rect 28262 17847 28264 17856
rect 28316 17847 28318 17856
rect 28264 17818 28316 17824
rect 28368 16794 28396 18158
rect 28356 16788 28408 16794
rect 28356 16730 28408 16736
rect 28460 15162 28488 19071
rect 28264 15156 28316 15162
rect 28264 15098 28316 15104
rect 28448 15156 28500 15162
rect 28448 15098 28500 15104
rect 28276 14822 28304 15098
rect 28448 15020 28500 15026
rect 28448 14962 28500 14968
rect 28264 14816 28316 14822
rect 28264 14758 28316 14764
rect 28356 14000 28408 14006
rect 28356 13942 28408 13948
rect 28262 13696 28318 13705
rect 28262 13631 28318 13640
rect 28276 13530 28304 13631
rect 28368 13530 28396 13942
rect 28264 13524 28316 13530
rect 28264 13466 28316 13472
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 28460 13410 28488 14962
rect 28552 14074 28580 23802
rect 28632 19712 28684 19718
rect 28632 19654 28684 19660
rect 28644 17338 28672 19654
rect 28736 19514 28764 35702
rect 29564 35494 29592 36722
rect 29644 36032 29696 36038
rect 29644 35974 29696 35980
rect 29656 35834 29684 35974
rect 29644 35828 29696 35834
rect 29644 35770 29696 35776
rect 29552 35488 29604 35494
rect 29552 35430 29604 35436
rect 29460 33856 29512 33862
rect 29460 33798 29512 33804
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 29012 28529 29040 30194
rect 28998 28520 29054 28529
rect 28998 28455 29054 28464
rect 29276 28416 29328 28422
rect 29276 28358 29328 28364
rect 29000 24200 29052 24206
rect 29000 24142 29052 24148
rect 28816 19984 28868 19990
rect 28816 19926 28868 19932
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28724 19168 28776 19174
rect 28724 19110 28776 19116
rect 28632 17332 28684 17338
rect 28632 17274 28684 17280
rect 28632 15904 28684 15910
rect 28632 15846 28684 15852
rect 28644 15366 28672 15846
rect 28632 15360 28684 15366
rect 28632 15302 28684 15308
rect 28736 14906 28764 19110
rect 28828 15026 28856 19926
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 28920 18170 28948 19314
rect 29012 18358 29040 24142
rect 29184 22568 29236 22574
rect 29184 22510 29236 22516
rect 29092 20800 29144 20806
rect 29092 20742 29144 20748
rect 29104 20466 29132 20742
rect 29092 20460 29144 20466
rect 29092 20402 29144 20408
rect 29104 20233 29132 20402
rect 29090 20224 29146 20233
rect 29090 20159 29146 20168
rect 29090 19544 29146 19553
rect 29090 19479 29146 19488
rect 29000 18352 29052 18358
rect 29000 18294 29052 18300
rect 28920 18142 29040 18170
rect 29012 17270 29040 18142
rect 29000 17264 29052 17270
rect 29000 17206 29052 17212
rect 28998 17096 29054 17105
rect 28998 17031 29054 17040
rect 28908 16992 28960 16998
rect 28908 16934 28960 16940
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 28736 14878 28856 14906
rect 28632 14816 28684 14822
rect 28632 14758 28684 14764
rect 28644 14521 28672 14758
rect 28630 14512 28686 14521
rect 28630 14447 28686 14456
rect 28540 14068 28592 14074
rect 28540 14010 28592 14016
rect 28552 13802 28580 14010
rect 28540 13796 28592 13802
rect 28540 13738 28592 13744
rect 28264 13388 28316 13394
rect 28264 13330 28316 13336
rect 28368 13382 28488 13410
rect 28172 12980 28224 12986
rect 28172 12922 28224 12928
rect 28184 12481 28212 12922
rect 28276 12889 28304 13330
rect 28262 12880 28318 12889
rect 28262 12815 28318 12824
rect 28170 12472 28226 12481
rect 28170 12407 28226 12416
rect 28276 10810 28304 12815
rect 28264 10804 28316 10810
rect 28264 10746 28316 10752
rect 28368 10130 28396 13382
rect 28448 12708 28500 12714
rect 28448 12650 28500 12656
rect 28356 10124 28408 10130
rect 28356 10066 28408 10072
rect 28356 7268 28408 7274
rect 28356 7210 28408 7216
rect 28080 5364 28132 5370
rect 28080 5306 28132 5312
rect 28264 5364 28316 5370
rect 28264 5306 28316 5312
rect 27988 4140 28040 4146
rect 27988 4082 28040 4088
rect 27816 3998 28120 4026
rect 27988 3936 28040 3942
rect 27988 3878 28040 3884
rect 28000 3534 28028 3878
rect 27988 3528 28040 3534
rect 27816 3488 27988 3516
rect 27344 3120 27396 3126
rect 27344 3062 27396 3068
rect 27436 3120 27488 3126
rect 27436 3062 27488 3068
rect 27712 3120 27764 3126
rect 27712 3062 27764 3068
rect 27344 2984 27396 2990
rect 27344 2926 27396 2932
rect 27356 2582 27384 2926
rect 27344 2576 27396 2582
rect 27344 2518 27396 2524
rect 27252 2372 27304 2378
rect 27252 2314 27304 2320
rect 27448 800 27476 3062
rect 27528 2508 27580 2514
rect 27528 2450 27580 2456
rect 27540 1358 27568 2450
rect 27528 1352 27580 1358
rect 27528 1294 27580 1300
rect 27816 800 27844 3488
rect 27988 3470 28040 3476
rect 28092 2774 28120 3998
rect 28172 3392 28224 3398
rect 28172 3334 28224 3340
rect 28000 2746 28120 2774
rect 28000 2009 28028 2746
rect 27986 2000 28042 2009
rect 27986 1935 28042 1944
rect 28184 1714 28212 3334
rect 28276 2310 28304 5306
rect 28368 3602 28396 7210
rect 28356 3596 28408 3602
rect 28356 3538 28408 3544
rect 28460 3126 28488 12650
rect 28552 12374 28580 13738
rect 28540 12368 28592 12374
rect 28540 12310 28592 12316
rect 28644 11898 28672 14447
rect 28632 11892 28684 11898
rect 28632 11834 28684 11840
rect 28644 11694 28672 11834
rect 28632 11688 28684 11694
rect 28632 11630 28684 11636
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28538 5536 28594 5545
rect 28538 5471 28594 5480
rect 28448 3120 28500 3126
rect 28448 3062 28500 3068
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 28368 2446 28396 2790
rect 28552 2582 28580 5471
rect 28644 4758 28672 8230
rect 28828 4826 28856 14878
rect 28920 12918 28948 16934
rect 29012 15008 29040 17031
rect 29104 16998 29132 19479
rect 29196 18306 29224 22510
rect 29288 18426 29316 28358
rect 29368 27668 29420 27674
rect 29368 27610 29420 27616
rect 29276 18420 29328 18426
rect 29276 18362 29328 18368
rect 29196 18278 29316 18306
rect 29184 18216 29236 18222
rect 29184 18158 29236 18164
rect 29196 17542 29224 18158
rect 29184 17536 29236 17542
rect 29184 17478 29236 17484
rect 29092 16992 29144 16998
rect 29092 16934 29144 16940
rect 29012 14980 29132 15008
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 29012 13462 29040 13806
rect 29000 13456 29052 13462
rect 29000 13398 29052 13404
rect 29012 12986 29040 13398
rect 29000 12980 29052 12986
rect 29000 12922 29052 12928
rect 28908 12912 28960 12918
rect 28908 12854 28960 12860
rect 28998 10160 29054 10169
rect 28998 10095 29054 10104
rect 29012 10062 29040 10095
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29104 6769 29132 14980
rect 29196 7818 29224 17478
rect 29288 17134 29316 18278
rect 29276 17128 29328 17134
rect 29276 17070 29328 17076
rect 29380 15706 29408 27610
rect 29472 19514 29500 33798
rect 29564 23118 29592 35430
rect 29552 23112 29604 23118
rect 29552 23054 29604 23060
rect 29748 20602 29776 37334
rect 29840 23322 29868 37742
rect 30024 37466 30052 38014
rect 30012 37460 30064 37466
rect 30012 37402 30064 37408
rect 30300 36904 30328 39222
rect 30378 39200 30434 40000
rect 30838 39200 30894 40000
rect 31206 39200 31262 40000
rect 31666 39200 31722 40000
rect 32034 39200 32090 40000
rect 32402 39200 32458 40000
rect 32862 39200 32918 40000
rect 33230 39200 33286 40000
rect 33690 39200 33746 40000
rect 34058 39200 34114 40000
rect 34426 39200 34482 40000
rect 34886 39200 34942 40000
rect 35254 39200 35310 40000
rect 35622 39200 35678 40000
rect 36082 39200 36138 40000
rect 36450 39200 36506 40000
rect 36910 39200 36966 40000
rect 37016 39222 37228 39250
rect 30392 37262 30420 39200
rect 30380 37256 30432 37262
rect 30432 37204 30512 37210
rect 30380 37198 30512 37204
rect 30392 37182 30512 37198
rect 30380 36916 30432 36922
rect 30300 36876 30380 36904
rect 30380 36858 30432 36864
rect 30380 36780 30432 36786
rect 30380 36722 30432 36728
rect 30104 36168 30156 36174
rect 30104 36110 30156 36116
rect 30116 35630 30144 36110
rect 30288 36032 30340 36038
rect 30288 35974 30340 35980
rect 30104 35624 30156 35630
rect 30104 35566 30156 35572
rect 30300 29345 30328 35974
rect 30392 34950 30420 36722
rect 30484 36378 30512 37182
rect 30748 37120 30800 37126
rect 30748 37062 30800 37068
rect 30472 36372 30524 36378
rect 30472 36314 30524 36320
rect 30380 34944 30432 34950
rect 30380 34886 30432 34892
rect 30286 29336 30342 29345
rect 30286 29271 30342 29280
rect 30196 26444 30248 26450
rect 30196 26386 30248 26392
rect 29920 24064 29972 24070
rect 29920 24006 29972 24012
rect 29828 23316 29880 23322
rect 29828 23258 29880 23264
rect 29828 22772 29880 22778
rect 29828 22714 29880 22720
rect 29736 20596 29788 20602
rect 29736 20538 29788 20544
rect 29748 19854 29776 20538
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29460 19508 29512 19514
rect 29460 19450 29512 19456
rect 29840 18578 29868 22714
rect 29748 18550 29868 18578
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29458 16824 29514 16833
rect 29458 16759 29514 16768
rect 29368 15700 29420 15706
rect 29368 15642 29420 15648
rect 29380 15502 29408 15642
rect 29368 15496 29420 15502
rect 29368 15438 29420 15444
rect 29274 14104 29330 14113
rect 29274 14039 29276 14048
rect 29328 14039 29330 14048
rect 29276 14010 29328 14016
rect 29288 13841 29316 14010
rect 29274 13832 29330 13841
rect 29274 13767 29330 13776
rect 29184 7812 29236 7818
rect 29184 7754 29236 7760
rect 29090 6760 29146 6769
rect 29090 6695 29146 6704
rect 28906 4856 28962 4865
rect 28816 4820 28868 4826
rect 28906 4791 28962 4800
rect 28816 4762 28868 4768
rect 28632 4752 28684 4758
rect 28632 4694 28684 4700
rect 28724 3936 28776 3942
rect 28724 3878 28776 3884
rect 28736 3058 28764 3878
rect 28828 3534 28856 4762
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 28920 3058 28948 4791
rect 29368 3936 29420 3942
rect 29368 3878 29420 3884
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 28724 3052 28776 3058
rect 28724 2994 28776 3000
rect 28908 3052 28960 3058
rect 28908 2994 28960 3000
rect 28540 2576 28592 2582
rect 28540 2518 28592 2524
rect 28356 2440 28408 2446
rect 28408 2400 28488 2428
rect 28356 2382 28408 2388
rect 28264 2304 28316 2310
rect 28264 2246 28316 2252
rect 28092 1686 28212 1714
rect 28092 800 28120 1686
rect 28460 800 28488 2400
rect 28736 800 28764 2994
rect 29104 800 29132 3334
rect 29380 2446 29408 3878
rect 29472 3777 29500 16759
rect 29552 16720 29604 16726
rect 29550 16688 29552 16697
rect 29604 16688 29606 16697
rect 29550 16623 29606 16632
rect 29656 15706 29684 17138
rect 29644 15700 29696 15706
rect 29644 15642 29696 15648
rect 29644 13184 29696 13190
rect 29644 13126 29696 13132
rect 29656 12986 29684 13126
rect 29748 13025 29776 18550
rect 29932 18442 29960 24006
rect 30104 23180 30156 23186
rect 30104 23122 30156 23128
rect 30012 23044 30064 23050
rect 30012 22986 30064 22992
rect 30024 22778 30052 22986
rect 30116 22778 30144 23122
rect 30012 22772 30064 22778
rect 30012 22714 30064 22720
rect 30104 22772 30156 22778
rect 30104 22714 30156 22720
rect 30208 22094 30236 26386
rect 30392 23798 30420 34886
rect 30654 29472 30710 29481
rect 30654 29407 30710 29416
rect 30380 23792 30432 23798
rect 30380 23734 30432 23740
rect 30472 23588 30524 23594
rect 30472 23530 30524 23536
rect 29840 18414 29960 18442
rect 30024 22066 30236 22094
rect 29734 13016 29790 13025
rect 29644 12980 29696 12986
rect 29734 12951 29790 12960
rect 29644 12922 29696 12928
rect 29840 12850 29868 18414
rect 29920 18284 29972 18290
rect 29920 18226 29972 18232
rect 29932 17542 29960 18226
rect 29920 17536 29972 17542
rect 29920 17478 29972 17484
rect 29828 12844 29880 12850
rect 29828 12786 29880 12792
rect 29932 12434 29960 17478
rect 30024 14618 30052 22066
rect 30196 19780 30248 19786
rect 30196 19722 30248 19728
rect 30208 19553 30236 19722
rect 30194 19544 30250 19553
rect 30194 19479 30250 19488
rect 30196 19372 30248 19378
rect 30196 19314 30248 19320
rect 30208 19174 30236 19314
rect 30286 19272 30342 19281
rect 30286 19207 30342 19216
rect 30196 19168 30248 19174
rect 30196 19110 30248 19116
rect 30104 18896 30156 18902
rect 30104 18838 30156 18844
rect 30012 14612 30064 14618
rect 30012 14554 30064 14560
rect 29840 12406 29960 12434
rect 29550 12336 29606 12345
rect 29550 12271 29552 12280
rect 29604 12271 29606 12280
rect 29552 12242 29604 12248
rect 29552 7540 29604 7546
rect 29552 7482 29604 7488
rect 29458 3768 29514 3777
rect 29458 3703 29514 3712
rect 29564 3534 29592 7482
rect 29840 6254 29868 12406
rect 29918 11520 29974 11529
rect 29918 11455 29974 11464
rect 29828 6248 29880 6254
rect 29828 6190 29880 6196
rect 29552 3528 29604 3534
rect 29552 3470 29604 3476
rect 29644 3120 29696 3126
rect 29644 3062 29696 3068
rect 29368 2440 29420 2446
rect 29368 2382 29420 2388
rect 29380 800 29408 2382
rect 29656 800 29684 3062
rect 29932 2378 29960 11455
rect 30116 3670 30144 18838
rect 30208 18698 30236 19110
rect 30196 18692 30248 18698
rect 30196 18634 30248 18640
rect 30300 18358 30328 19207
rect 30288 18352 30340 18358
rect 30288 18294 30340 18300
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30392 13569 30420 17070
rect 30378 13560 30434 13569
rect 30378 13495 30434 13504
rect 30484 13433 30512 23530
rect 30564 23044 30616 23050
rect 30564 22986 30616 22992
rect 30576 22438 30604 22986
rect 30564 22432 30616 22438
rect 30562 22400 30564 22409
rect 30616 22400 30618 22409
rect 30562 22335 30618 22344
rect 30668 19990 30696 29407
rect 30656 19984 30708 19990
rect 30656 19926 30708 19932
rect 30564 18828 30616 18834
rect 30564 18770 30616 18776
rect 30470 13424 30526 13433
rect 30470 13359 30526 13368
rect 30576 10538 30604 18770
rect 30760 18766 30788 37062
rect 30852 36922 30880 39200
rect 30840 36916 30892 36922
rect 30840 36858 30892 36864
rect 31024 36780 31076 36786
rect 31024 36722 31076 36728
rect 31036 35494 31064 36722
rect 31220 36378 31248 39200
rect 31680 37346 31708 39200
rect 31680 37318 31800 37346
rect 31772 37262 31800 37318
rect 31760 37256 31812 37262
rect 31760 37198 31812 37204
rect 32048 36922 32076 39200
rect 32416 36922 32444 39200
rect 32876 37262 32904 39200
rect 32864 37256 32916 37262
rect 32864 37198 32916 37204
rect 33140 37256 33192 37262
rect 33140 37198 33192 37204
rect 32036 36916 32088 36922
rect 32036 36858 32088 36864
rect 32404 36916 32456 36922
rect 32404 36858 32456 36864
rect 32128 36780 32180 36786
rect 32128 36722 32180 36728
rect 32680 36780 32732 36786
rect 32680 36722 32732 36728
rect 31208 36372 31260 36378
rect 31208 36314 31260 36320
rect 31116 36168 31168 36174
rect 31116 36110 31168 36116
rect 31024 35488 31076 35494
rect 31024 35430 31076 35436
rect 30932 22976 30984 22982
rect 30932 22918 30984 22924
rect 30748 18760 30800 18766
rect 30748 18702 30800 18708
rect 30840 18080 30892 18086
rect 30840 18022 30892 18028
rect 30656 14272 30708 14278
rect 30656 14214 30708 14220
rect 30564 10532 30616 10538
rect 30564 10474 30616 10480
rect 30668 10266 30696 14214
rect 30852 14074 30880 18022
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 30944 11665 30972 22918
rect 31036 19242 31064 35430
rect 31128 34950 31156 36110
rect 32140 36038 32168 36722
rect 32128 36032 32180 36038
rect 32128 35974 32180 35980
rect 32692 35494 32720 36722
rect 33152 36378 33180 37198
rect 33244 36922 33272 39200
rect 33324 37732 33376 37738
rect 33324 37674 33376 37680
rect 33336 37466 33364 37674
rect 33324 37460 33376 37466
rect 33324 37402 33376 37408
rect 33232 36916 33284 36922
rect 33232 36858 33284 36864
rect 33508 36780 33560 36786
rect 33508 36722 33560 36728
rect 33140 36372 33192 36378
rect 33140 36314 33192 36320
rect 33520 35698 33548 36722
rect 33704 36378 33732 39200
rect 34072 37262 34100 39200
rect 34060 37256 34112 37262
rect 34060 37198 34112 37204
rect 34440 36904 34468 39200
rect 34900 37754 34928 39200
rect 34808 37726 34928 37754
rect 35268 37754 35296 39200
rect 35268 37726 35388 37754
rect 34704 37664 34756 37670
rect 34704 37606 34756 37612
rect 34716 37466 34744 37606
rect 34704 37460 34756 37466
rect 34704 37402 34756 37408
rect 34520 36916 34572 36922
rect 34440 36876 34520 36904
rect 34520 36858 34572 36864
rect 34244 36780 34296 36786
rect 34244 36722 34296 36728
rect 33692 36372 33744 36378
rect 33692 36314 33744 36320
rect 33600 36168 33652 36174
rect 33600 36110 33652 36116
rect 33508 35692 33560 35698
rect 33508 35634 33560 35640
rect 32680 35488 32732 35494
rect 32680 35430 32732 35436
rect 32692 35154 32720 35430
rect 32680 35148 32732 35154
rect 32680 35090 32732 35096
rect 33612 34950 33640 36110
rect 34256 35494 34284 36722
rect 34808 36378 34836 37726
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 35360 37262 35388 37726
rect 35348 37256 35400 37262
rect 35348 37198 35400 37204
rect 35636 36922 35664 39200
rect 35808 37868 35860 37874
rect 35808 37810 35860 37816
rect 35820 37398 35848 37810
rect 35808 37392 35860 37398
rect 35808 37334 35860 37340
rect 35716 37256 35768 37262
rect 35716 37198 35768 37204
rect 35624 36916 35676 36922
rect 35624 36858 35676 36864
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35728 36378 35756 37198
rect 36096 36922 36124 39200
rect 36084 36916 36136 36922
rect 36084 36858 36136 36864
rect 36464 36802 36492 39200
rect 36924 39114 36952 39200
rect 37016 39114 37044 39222
rect 36924 39086 37044 39114
rect 37200 36904 37228 39222
rect 37278 39200 37334 40000
rect 37646 39200 37702 40000
rect 38106 39200 38162 40000
rect 38474 39200 38530 40000
rect 38934 39200 38990 40000
rect 39302 39200 39358 40000
rect 39670 39200 39726 40000
rect 39776 39222 39988 39250
rect 37292 37074 37320 39200
rect 37660 37262 37688 39200
rect 37832 37800 37884 37806
rect 37832 37742 37884 37748
rect 37844 37466 37872 37742
rect 37832 37460 37884 37466
rect 37832 37402 37884 37408
rect 37648 37256 37700 37262
rect 37648 37198 37700 37204
rect 37292 37046 37412 37074
rect 37280 36916 37332 36922
rect 37200 36876 37280 36904
rect 37280 36858 37332 36864
rect 36464 36786 36584 36802
rect 35992 36780 36044 36786
rect 35992 36722 36044 36728
rect 36268 36780 36320 36786
rect 36464 36780 36596 36786
rect 36464 36774 36544 36780
rect 36268 36722 36320 36728
rect 36544 36722 36596 36728
rect 37096 36780 37148 36786
rect 37096 36722 37148 36728
rect 36004 36378 36032 36722
rect 34796 36372 34848 36378
rect 34796 36314 34848 36320
rect 35716 36372 35768 36378
rect 35716 36314 35768 36320
rect 35992 36372 36044 36378
rect 35992 36314 36044 36320
rect 34704 36168 34756 36174
rect 34704 36110 34756 36116
rect 34716 35494 34744 36110
rect 34244 35488 34296 35494
rect 34244 35430 34296 35436
rect 34704 35488 34756 35494
rect 34704 35430 34756 35436
rect 31116 34944 31168 34950
rect 31116 34886 31168 34892
rect 33600 34944 33652 34950
rect 33600 34886 33652 34892
rect 31128 30433 31156 34886
rect 33612 34746 33640 34886
rect 33600 34740 33652 34746
rect 33600 34682 33652 34688
rect 32772 32428 32824 32434
rect 32772 32370 32824 32376
rect 31114 30424 31170 30433
rect 31114 30359 31170 30368
rect 31116 27872 31168 27878
rect 31116 27814 31168 27820
rect 31024 19236 31076 19242
rect 31024 19178 31076 19184
rect 31128 14793 31156 27814
rect 31850 26752 31906 26761
rect 31850 26687 31906 26696
rect 31576 26512 31628 26518
rect 31576 26454 31628 26460
rect 31300 23044 31352 23050
rect 31300 22986 31352 22992
rect 31312 22438 31340 22986
rect 31300 22432 31352 22438
rect 31298 22400 31300 22409
rect 31352 22400 31354 22409
rect 31298 22335 31354 22344
rect 31300 22024 31352 22030
rect 31300 21966 31352 21972
rect 31208 21548 31260 21554
rect 31208 21490 31260 21496
rect 31114 14784 31170 14793
rect 31114 14719 31170 14728
rect 30930 11656 30986 11665
rect 30930 11591 30986 11600
rect 30656 10260 30708 10266
rect 30656 10202 30708 10208
rect 31220 9110 31248 21490
rect 31312 11626 31340 21966
rect 31392 19712 31444 19718
rect 31390 19680 31392 19689
rect 31444 19680 31446 19689
rect 31390 19615 31446 19624
rect 31588 16289 31616 26454
rect 31760 25356 31812 25362
rect 31760 25298 31812 25304
rect 31666 21448 31722 21457
rect 31666 21383 31722 21392
rect 31680 19281 31708 21383
rect 31772 19378 31800 25298
rect 31760 19372 31812 19378
rect 31760 19314 31812 19320
rect 31666 19272 31722 19281
rect 31666 19207 31722 19216
rect 31666 18320 31722 18329
rect 31666 18255 31722 18264
rect 31574 16280 31630 16289
rect 31574 16215 31630 16224
rect 31680 12481 31708 18255
rect 31760 18148 31812 18154
rect 31760 18090 31812 18096
rect 31666 12472 31722 12481
rect 31666 12407 31722 12416
rect 31666 12336 31722 12345
rect 31666 12271 31722 12280
rect 31300 11620 31352 11626
rect 31300 11562 31352 11568
rect 31680 9353 31708 12271
rect 31666 9344 31722 9353
rect 31666 9279 31722 9288
rect 31208 9104 31260 9110
rect 31208 9046 31260 9052
rect 31024 6928 31076 6934
rect 31024 6870 31076 6876
rect 30196 5568 30248 5574
rect 30196 5510 30248 5516
rect 30104 3664 30156 3670
rect 30104 3606 30156 3612
rect 30012 3392 30064 3398
rect 30012 3334 30064 3340
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 30024 800 30052 3334
rect 30208 3058 30236 5510
rect 30288 3936 30340 3942
rect 30288 3878 30340 3884
rect 30748 3936 30800 3942
rect 30748 3878 30800 3884
rect 30300 3126 30328 3878
rect 30288 3120 30340 3126
rect 30288 3062 30340 3068
rect 30656 3120 30708 3126
rect 30656 3062 30708 3068
rect 30196 3052 30248 3058
rect 30196 2994 30248 3000
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 30288 2372 30340 2378
rect 30288 2314 30340 2320
rect 30300 800 30328 2314
rect 30392 1465 30420 2382
rect 30378 1456 30434 1465
rect 30378 1391 30434 1400
rect 30668 800 30696 3062
rect 30760 2378 30788 3878
rect 31036 3534 31064 6870
rect 31116 6860 31168 6866
rect 31116 6802 31168 6808
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 30932 3392 30984 3398
rect 30932 3334 30984 3340
rect 30748 2372 30800 2378
rect 30748 2314 30800 2320
rect 30944 800 30972 3334
rect 31128 2038 31156 6802
rect 31772 6458 31800 18090
rect 31864 9897 31892 26687
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32126 23352 32182 23361
rect 32126 23287 32182 23296
rect 31942 21992 31998 22001
rect 31942 21927 31998 21936
rect 31850 9888 31906 9897
rect 31850 9823 31906 9832
rect 31956 7993 31984 21927
rect 32036 19712 32088 19718
rect 32036 19654 32088 19660
rect 32048 19553 32076 19654
rect 32034 19544 32090 19553
rect 32034 19479 32090 19488
rect 32036 19372 32088 19378
rect 32036 19314 32088 19320
rect 32048 11286 32076 19314
rect 32036 11280 32088 11286
rect 32036 11222 32088 11228
rect 32140 10742 32168 23287
rect 32324 22982 32352 23666
rect 32312 22976 32364 22982
rect 32312 22918 32364 22924
rect 32220 21004 32272 21010
rect 32220 20946 32272 20952
rect 32128 10736 32180 10742
rect 32128 10678 32180 10684
rect 32232 10606 32260 20946
rect 32324 12753 32352 22918
rect 32586 20224 32642 20233
rect 32586 20159 32642 20168
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 32416 19174 32444 19314
rect 32404 19168 32456 19174
rect 32404 19110 32456 19116
rect 32310 12744 32366 12753
rect 32310 12679 32366 12688
rect 32220 10600 32272 10606
rect 32220 10542 32272 10548
rect 31942 7984 31998 7993
rect 31942 7919 31998 7928
rect 31760 6452 31812 6458
rect 31760 6394 31812 6400
rect 31208 3936 31260 3942
rect 31208 3878 31260 3884
rect 31668 3936 31720 3942
rect 31668 3878 31720 3884
rect 31220 3126 31248 3878
rect 31208 3120 31260 3126
rect 31208 3062 31260 3068
rect 31680 3058 31708 3878
rect 31942 3632 31998 3641
rect 31942 3567 31998 3576
rect 31956 3534 31984 3567
rect 31944 3528 31996 3534
rect 31944 3470 31996 3476
rect 32416 3466 32444 19110
rect 32600 7410 32628 20159
rect 32784 20058 32812 32370
rect 33140 29708 33192 29714
rect 33140 29650 33192 29656
rect 32862 26616 32918 26625
rect 32862 26551 32918 26560
rect 32772 20052 32824 20058
rect 32772 19994 32824 20000
rect 32678 8800 32734 8809
rect 32678 8735 32734 8744
rect 32588 7404 32640 7410
rect 32588 7346 32640 7352
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 31852 3392 31904 3398
rect 31852 3334 31904 3340
rect 31668 3052 31720 3058
rect 31668 2994 31720 3000
rect 31680 2774 31708 2994
rect 31588 2746 31708 2774
rect 31300 2372 31352 2378
rect 31300 2314 31352 2320
rect 31116 2032 31168 2038
rect 31116 1974 31168 1980
rect 31312 800 31340 2314
rect 31588 800 31616 2746
rect 31864 800 31892 3334
rect 32496 3120 32548 3126
rect 32496 3062 32548 3068
rect 32220 2508 32272 2514
rect 32220 2450 32272 2456
rect 32232 800 32260 2450
rect 32508 800 32536 3062
rect 32692 2582 32720 8735
rect 32876 7449 32904 26551
rect 33152 19514 33180 29650
rect 33232 26376 33284 26382
rect 33232 26318 33284 26324
rect 33140 19508 33192 19514
rect 33140 19450 33192 19456
rect 33244 11937 33272 26318
rect 33508 24880 33560 24886
rect 33508 24822 33560 24828
rect 33416 19848 33468 19854
rect 33416 19790 33468 19796
rect 33324 19440 33376 19446
rect 33324 19382 33376 19388
rect 33230 11928 33286 11937
rect 33230 11863 33286 11872
rect 33336 9110 33364 19382
rect 33324 9104 33376 9110
rect 33324 9046 33376 9052
rect 33428 8537 33456 19790
rect 33520 14278 33548 24822
rect 33600 20392 33652 20398
rect 33600 20334 33652 20340
rect 33508 14272 33560 14278
rect 33508 14214 33560 14220
rect 33612 9217 33640 20334
rect 33784 20256 33836 20262
rect 33784 20198 33836 20204
rect 33796 19786 33824 20198
rect 33784 19780 33836 19786
rect 33784 19722 33836 19728
rect 33796 19689 33824 19722
rect 33782 19680 33838 19689
rect 33782 19615 33838 19624
rect 33968 19372 34020 19378
rect 33968 19314 34020 19320
rect 33980 18630 34008 19314
rect 34256 19242 34284 35430
rect 34520 34944 34572 34950
rect 34520 34886 34572 34892
rect 34532 30569 34560 34886
rect 34716 34649 34744 35430
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34702 34640 34758 34649
rect 34702 34575 34758 34584
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 35348 32496 35400 32502
rect 35348 32438 35400 32444
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34518 30560 34574 30569
rect 34518 30495 34574 30504
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34518 29064 34574 29073
rect 34518 28999 34574 29008
rect 34244 19236 34296 19242
rect 34244 19178 34296 19184
rect 33968 18624 34020 18630
rect 33968 18566 34020 18572
rect 33980 16574 34008 18566
rect 33980 16546 34100 16574
rect 33690 10432 33746 10441
rect 33690 10367 33746 10376
rect 33598 9208 33654 9217
rect 33598 9143 33654 9152
rect 33414 8528 33470 8537
rect 33414 8463 33470 8472
rect 32954 7848 33010 7857
rect 32954 7783 33010 7792
rect 32862 7440 32918 7449
rect 32862 7375 32918 7384
rect 32770 6216 32826 6225
rect 32770 6151 32826 6160
rect 32784 3194 32812 6151
rect 32968 3534 32996 7783
rect 33508 4480 33560 4486
rect 33508 4422 33560 4428
rect 33048 4072 33100 4078
rect 33048 4014 33100 4020
rect 32956 3528 33008 3534
rect 32956 3470 33008 3476
rect 32864 3392 32916 3398
rect 32864 3334 32916 3340
rect 32772 3188 32824 3194
rect 32772 3130 32824 3136
rect 32680 2576 32732 2582
rect 32680 2518 32732 2524
rect 32876 800 32904 3334
rect 33060 3126 33088 4014
rect 33324 3936 33376 3942
rect 33324 3878 33376 3884
rect 33048 3120 33100 3126
rect 33048 3062 33100 3068
rect 33230 2952 33286 2961
rect 33230 2887 33232 2896
rect 33284 2887 33286 2896
rect 33232 2858 33284 2864
rect 33336 2514 33364 3878
rect 33520 3058 33548 4422
rect 33508 3052 33560 3058
rect 33508 2994 33560 3000
rect 33324 2508 33376 2514
rect 33324 2450 33376 2456
rect 33140 2372 33192 2378
rect 33140 2314 33192 2320
rect 33152 800 33180 2314
rect 33520 800 33548 2994
rect 33704 2650 33732 10367
rect 33874 5264 33930 5273
rect 33874 5199 33930 5208
rect 33888 3534 33916 5199
rect 34072 5137 34100 16546
rect 34532 8129 34560 28999
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34794 27704 34850 27713
rect 34934 27696 35242 27716
rect 34794 27639 34850 27648
rect 34704 22772 34756 22778
rect 34704 22714 34756 22720
rect 34612 19780 34664 19786
rect 34612 19722 34664 19728
rect 34624 19174 34652 19722
rect 34612 19168 34664 19174
rect 34612 19110 34664 19116
rect 34624 12646 34652 19110
rect 34612 12640 34664 12646
rect 34612 12582 34664 12588
rect 34716 9081 34744 22714
rect 34808 12073 34836 27639
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 35360 19310 35388 32438
rect 36004 24138 36032 36314
rect 36280 35494 36308 36722
rect 37108 36378 37136 36722
rect 37280 36644 37332 36650
rect 37280 36586 37332 36592
rect 37096 36372 37148 36378
rect 37096 36314 37148 36320
rect 36268 35488 36320 35494
rect 36268 35430 36320 35436
rect 35992 24132 36044 24138
rect 35992 24074 36044 24080
rect 35438 21040 35494 21049
rect 35438 20975 35494 20984
rect 35348 19304 35400 19310
rect 35348 19246 35400 19252
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34794 12064 34850 12073
rect 34794 11999 34850 12008
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 35452 10577 35480 20975
rect 35530 20496 35586 20505
rect 35530 20431 35586 20440
rect 35438 10568 35494 10577
rect 35438 10503 35494 10512
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34702 9072 34758 9081
rect 34702 9007 34758 9016
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34518 8120 34574 8129
rect 34934 8112 35242 8132
rect 34518 8055 34574 8064
rect 34150 7576 34206 7585
rect 34150 7511 34206 7520
rect 34058 5128 34114 5137
rect 34058 5063 34114 5072
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 33796 800 33824 3334
rect 34164 2922 34192 7511
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34520 5908 34572 5914
rect 34520 5850 34572 5856
rect 34532 3534 34560 5850
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34796 4480 34848 4486
rect 34796 4422 34848 4428
rect 35348 4480 35400 4486
rect 35348 4422 35400 4428
rect 34612 3936 34664 3942
rect 34612 3878 34664 3884
rect 34520 3528 34572 3534
rect 34520 3470 34572 3476
rect 34520 3120 34572 3126
rect 34518 3088 34520 3097
rect 34572 3088 34574 3097
rect 34428 3052 34480 3058
rect 34518 3023 34574 3032
rect 34428 2994 34480 3000
rect 34152 2916 34204 2922
rect 34152 2858 34204 2864
rect 34060 2440 34112 2446
rect 34060 2382 34112 2388
rect 34072 800 34100 2382
rect 34440 800 34468 2994
rect 34624 2378 34652 3878
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 34612 2372 34664 2378
rect 34612 2314 34664 2320
rect 34716 800 34744 3334
rect 34808 3058 34836 4422
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35360 3058 35388 4422
rect 35440 3936 35492 3942
rect 35440 3878 35492 3884
rect 34796 3052 34848 3058
rect 34796 2994 34848 3000
rect 35348 3052 35400 3058
rect 35348 2994 35400 3000
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35072 2576 35124 2582
rect 35070 2544 35072 2553
rect 35124 2544 35126 2553
rect 34980 2508 35032 2514
rect 35070 2479 35126 2488
rect 34980 2450 35032 2456
rect 34992 2038 35020 2450
rect 35072 2440 35124 2446
rect 35072 2382 35124 2388
rect 34980 2032 35032 2038
rect 34980 1974 35032 1980
rect 35084 800 35112 2382
rect 35360 800 35388 2994
rect 35452 2378 35480 3878
rect 35544 3194 35572 20431
rect 35624 19780 35676 19786
rect 35624 19722 35676 19728
rect 35636 19174 35664 19722
rect 35624 19168 35676 19174
rect 35624 19110 35676 19116
rect 35636 18902 35664 19110
rect 36280 18970 36308 35430
rect 37292 32473 37320 36586
rect 37384 36378 37412 37046
rect 37832 36780 37884 36786
rect 37832 36722 37884 36728
rect 37372 36372 37424 36378
rect 37372 36314 37424 36320
rect 37844 35494 37872 36722
rect 38016 36168 38068 36174
rect 38016 36110 38068 36116
rect 37832 35488 37884 35494
rect 37832 35430 37884 35436
rect 37278 32464 37334 32473
rect 37278 32399 37334 32408
rect 37844 20058 37872 35430
rect 38028 35290 38056 36110
rect 38120 35834 38148 39200
rect 38384 37256 38436 37262
rect 38384 37198 38436 37204
rect 38396 36922 38424 37198
rect 38384 36916 38436 36922
rect 38384 36858 38436 36864
rect 38108 35828 38160 35834
rect 38108 35770 38160 35776
rect 38488 35766 38516 39200
rect 38948 37262 38976 39200
rect 38568 37256 38620 37262
rect 38568 37198 38620 37204
rect 38936 37256 38988 37262
rect 38936 37198 38988 37204
rect 38476 35760 38528 35766
rect 38476 35702 38528 35708
rect 38580 35494 38608 37198
rect 38844 37120 38896 37126
rect 38844 37062 38896 37068
rect 38660 36168 38712 36174
rect 38660 36110 38712 36116
rect 38568 35488 38620 35494
rect 38568 35430 38620 35436
rect 38016 35284 38068 35290
rect 38016 35226 38068 35232
rect 38028 34950 38056 35226
rect 38016 34944 38068 34950
rect 38016 34886 38068 34892
rect 38580 26234 38608 35430
rect 38672 34950 38700 36110
rect 38856 35834 38884 37062
rect 39316 36922 39344 39200
rect 39684 39114 39712 39200
rect 39776 39114 39804 39222
rect 39684 39086 39804 39114
rect 39304 36916 39356 36922
rect 39304 36858 39356 36864
rect 39212 36780 39264 36786
rect 39212 36722 39264 36728
rect 38936 36032 38988 36038
rect 38936 35974 38988 35980
rect 38844 35828 38896 35834
rect 38844 35770 38896 35776
rect 38948 35766 38976 35974
rect 38936 35760 38988 35766
rect 38936 35702 38988 35708
rect 39224 35494 39252 36722
rect 39960 36360 39988 39222
rect 40130 39200 40186 40000
rect 40498 39200 40554 40000
rect 40866 39200 40922 40000
rect 41326 39200 41382 40000
rect 41694 39200 41750 40000
rect 42154 39200 42210 40000
rect 42522 39200 42578 40000
rect 42890 39200 42946 40000
rect 43350 39200 43406 40000
rect 43718 39200 43774 40000
rect 44178 39200 44234 40000
rect 44546 39200 44602 40000
rect 44914 39200 44970 40000
rect 45374 39200 45430 40000
rect 45742 39200 45798 40000
rect 40144 37346 40172 39200
rect 40408 37460 40460 37466
rect 40408 37402 40460 37408
rect 40420 37369 40448 37402
rect 40406 37360 40462 37369
rect 40144 37318 40264 37346
rect 40132 37256 40184 37262
rect 40132 37198 40184 37204
rect 40040 36372 40092 36378
rect 39960 36332 40040 36360
rect 40040 36314 40092 36320
rect 39856 36168 39908 36174
rect 39856 36110 39908 36116
rect 39212 35488 39264 35494
rect 39212 35430 39264 35436
rect 38660 34944 38712 34950
rect 38660 34886 38712 34892
rect 38488 26206 38608 26234
rect 38488 23254 38516 26206
rect 38672 24206 38700 34886
rect 38660 24200 38712 24206
rect 38660 24142 38712 24148
rect 38476 23248 38528 23254
rect 38476 23190 38528 23196
rect 39224 23186 39252 35430
rect 39868 34950 39896 36110
rect 40144 35834 40172 37198
rect 40236 37194 40264 37318
rect 40406 37295 40462 37304
rect 40224 37188 40276 37194
rect 40224 37130 40276 37136
rect 40512 36922 40540 39200
rect 40500 36916 40552 36922
rect 40500 36858 40552 36864
rect 40592 36780 40644 36786
rect 40592 36722 40644 36728
rect 40132 35828 40184 35834
rect 40132 35770 40184 35776
rect 40604 35494 40632 36722
rect 40880 36378 40908 39200
rect 41234 37904 41290 37913
rect 41234 37839 41290 37848
rect 41248 37466 41276 37839
rect 41236 37460 41288 37466
rect 41236 37402 41288 37408
rect 41340 36802 41368 39200
rect 41512 37188 41564 37194
rect 41512 37130 41564 37136
rect 41340 36786 41460 36802
rect 41340 36780 41472 36786
rect 41340 36774 41420 36780
rect 41420 36722 41472 36728
rect 40868 36372 40920 36378
rect 40868 36314 40920 36320
rect 40776 36168 40828 36174
rect 40776 36110 40828 36116
rect 40592 35488 40644 35494
rect 40592 35430 40644 35436
rect 39856 34944 39908 34950
rect 39856 34886 39908 34892
rect 39868 28422 39896 34886
rect 39856 28416 39908 28422
rect 39856 28358 39908 28364
rect 39212 23180 39264 23186
rect 39212 23122 39264 23128
rect 40604 23118 40632 35430
rect 40788 34950 40816 36110
rect 41432 35834 41460 36722
rect 41524 36378 41552 37130
rect 41708 37126 41736 39200
rect 41696 37120 41748 37126
rect 41696 37062 41748 37068
rect 42168 36922 42196 39200
rect 42340 37256 42392 37262
rect 42340 37198 42392 37204
rect 42156 36916 42208 36922
rect 42156 36858 42208 36864
rect 41604 36576 41656 36582
rect 41604 36518 41656 36524
rect 41512 36372 41564 36378
rect 41512 36314 41564 36320
rect 41420 35828 41472 35834
rect 41420 35770 41472 35776
rect 40776 34944 40828 34950
rect 40776 34886 40828 34892
rect 41328 34944 41380 34950
rect 41328 34886 41380 34892
rect 40592 23112 40644 23118
rect 40592 23054 40644 23060
rect 40788 21457 40816 34886
rect 41340 29714 41368 34886
rect 41328 29708 41380 29714
rect 41328 29650 41380 29656
rect 41616 29646 41644 36518
rect 42352 36378 42380 37198
rect 42904 37126 42932 39200
rect 43076 37256 43128 37262
rect 43076 37198 43128 37204
rect 42892 37120 42944 37126
rect 42892 37062 42944 37068
rect 42432 36780 42484 36786
rect 42432 36722 42484 36728
rect 42340 36372 42392 36378
rect 42340 36314 42392 36320
rect 41604 29640 41656 29646
rect 41604 29582 41656 29588
rect 42352 26234 42380 36314
rect 42444 35494 42472 36722
rect 43088 36378 43116 37198
rect 43364 36922 43392 39200
rect 43444 37256 43496 37262
rect 43444 37198 43496 37204
rect 43352 36916 43404 36922
rect 43352 36858 43404 36864
rect 43168 36780 43220 36786
rect 43168 36722 43220 36728
rect 43076 36372 43128 36378
rect 43076 36314 43128 36320
rect 42432 35488 42484 35494
rect 42432 35430 42484 35436
rect 42260 26206 42380 26234
rect 42260 23526 42288 26206
rect 42248 23520 42300 23526
rect 42248 23462 42300 23468
rect 42444 23050 42472 35430
rect 43088 32434 43116 36314
rect 43180 34950 43208 36722
rect 43456 35894 43484 37198
rect 44192 37126 44220 39200
rect 44180 37120 44232 37126
rect 44180 37062 44232 37068
rect 43536 36780 43588 36786
rect 43536 36722 43588 36728
rect 43364 35866 43484 35894
rect 43364 35494 43392 35866
rect 43352 35488 43404 35494
rect 43352 35430 43404 35436
rect 43168 34944 43220 34950
rect 43168 34886 43220 34892
rect 43076 32428 43128 32434
rect 43076 32370 43128 32376
rect 42432 23044 42484 23050
rect 42432 22986 42484 22992
rect 40774 21448 40830 21457
rect 40774 21383 40830 21392
rect 37832 20052 37884 20058
rect 37832 19994 37884 20000
rect 43364 19854 43392 35430
rect 43548 34950 43576 36722
rect 44560 36378 44588 39200
rect 45388 36922 45416 39200
rect 45376 36916 45428 36922
rect 45376 36858 45428 36864
rect 44548 36372 44600 36378
rect 44548 36314 44600 36320
rect 43720 36168 43772 36174
rect 43720 36110 43772 36116
rect 43628 35692 43680 35698
rect 43628 35634 43680 35640
rect 43536 34944 43588 34950
rect 43536 34886 43588 34892
rect 43548 19922 43576 34886
rect 43640 33862 43668 35634
rect 43732 34542 43760 36110
rect 45756 35834 45784 39200
rect 45744 35828 45796 35834
rect 45744 35770 45796 35776
rect 43720 34536 43772 34542
rect 43720 34478 43772 34484
rect 43628 33856 43680 33862
rect 43628 33798 43680 33804
rect 43640 19990 43668 33798
rect 43732 32502 43760 34478
rect 43720 32496 43772 32502
rect 43720 32438 43772 32444
rect 44088 30048 44140 30054
rect 44086 30016 44088 30025
rect 44140 30016 44142 30025
rect 44086 29951 44142 29960
rect 43628 19984 43680 19990
rect 43628 19926 43680 19932
rect 43536 19916 43588 19922
rect 43536 19858 43588 19864
rect 43352 19848 43404 19854
rect 43352 19790 43404 19796
rect 36268 18964 36320 18970
rect 36268 18906 36320 18912
rect 35624 18896 35676 18902
rect 35624 18838 35676 18844
rect 43996 18692 44048 18698
rect 43996 18634 44048 18640
rect 41604 17332 41656 17338
rect 41604 17274 41656 17280
rect 37924 16992 37976 16998
rect 37924 16934 37976 16940
rect 35898 14376 35954 14385
rect 35898 14311 35954 14320
rect 35912 4826 35940 14311
rect 37462 6624 37518 6633
rect 37462 6559 37518 6568
rect 35900 4820 35952 4826
rect 35900 4762 35952 4768
rect 35912 3534 35940 4762
rect 37096 4752 37148 4758
rect 37096 4694 37148 4700
rect 36636 4480 36688 4486
rect 36636 4422 36688 4428
rect 36084 3936 36136 3942
rect 36084 3878 36136 3884
rect 36268 3936 36320 3942
rect 36268 3878 36320 3884
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 35624 3392 35676 3398
rect 35624 3334 35676 3340
rect 35532 3188 35584 3194
rect 35532 3130 35584 3136
rect 35440 2372 35492 2378
rect 35440 2314 35492 2320
rect 35532 2304 35584 2310
rect 35532 2246 35584 2252
rect 35544 1766 35572 2246
rect 35532 1760 35584 1766
rect 35532 1702 35584 1708
rect 35636 800 35664 3334
rect 35992 3120 36044 3126
rect 35992 3062 36044 3068
rect 36004 800 36032 3062
rect 36096 2446 36124 3878
rect 36280 3058 36308 3878
rect 36648 3534 36676 4422
rect 36912 4072 36964 4078
rect 36912 4014 36964 4020
rect 36636 3528 36688 3534
rect 36636 3470 36688 3476
rect 36636 3392 36688 3398
rect 36636 3334 36688 3340
rect 36268 3052 36320 3058
rect 36268 2994 36320 3000
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36280 800 36308 2994
rect 36648 800 36676 3334
rect 36924 2990 36952 4014
rect 36912 2984 36964 2990
rect 36912 2926 36964 2932
rect 36924 800 36952 2926
rect 37108 2582 37136 4694
rect 37280 4480 37332 4486
rect 37280 4422 37332 4428
rect 37188 3936 37240 3942
rect 37188 3878 37240 3884
rect 37200 3126 37228 3878
rect 37292 3466 37320 4422
rect 37372 4004 37424 4010
rect 37372 3946 37424 3952
rect 37280 3460 37332 3466
rect 37280 3402 37332 3408
rect 37188 3120 37240 3126
rect 37188 3062 37240 3068
rect 37096 2576 37148 2582
rect 37096 2518 37148 2524
rect 37292 800 37320 3402
rect 37384 3194 37412 3946
rect 37476 3738 37504 6559
rect 37936 4826 37964 16934
rect 41616 16574 41644 17274
rect 43904 17264 43956 17270
rect 43904 17206 43956 17212
rect 41616 16546 41736 16574
rect 38014 10024 38070 10033
rect 38014 9959 38070 9968
rect 37924 4820 37976 4826
rect 37924 4762 37976 4768
rect 37464 3732 37516 3738
rect 37464 3674 37516 3680
rect 37936 3534 37964 4762
rect 37924 3528 37976 3534
rect 37924 3470 37976 3476
rect 37648 3392 37700 3398
rect 37568 3352 37648 3380
rect 37372 3188 37424 3194
rect 37372 3130 37424 3136
rect 37568 800 37596 3352
rect 37648 3334 37700 3340
rect 38028 3126 38056 9959
rect 41420 9172 41472 9178
rect 41420 9114 41472 9120
rect 40776 8560 40828 8566
rect 40776 8502 40828 8508
rect 40788 4826 40816 8502
rect 41432 5370 41460 9114
rect 41708 5574 41736 16546
rect 42062 14920 42118 14929
rect 42062 14855 42118 14864
rect 42076 6866 42104 14855
rect 42522 11792 42578 11801
rect 42522 11727 42578 11736
rect 42246 11656 42302 11665
rect 42246 11591 42302 11600
rect 42156 9376 42208 9382
rect 42156 9318 42208 9324
rect 42064 6860 42116 6866
rect 42064 6802 42116 6808
rect 42168 5574 42196 9318
rect 41696 5568 41748 5574
rect 41696 5510 41748 5516
rect 42156 5568 42208 5574
rect 42156 5510 42208 5516
rect 41420 5364 41472 5370
rect 41420 5306 41472 5312
rect 40776 4820 40828 4826
rect 40776 4762 40828 4768
rect 39120 4616 39172 4622
rect 39120 4558 39172 4564
rect 38660 4480 38712 4486
rect 38660 4422 38712 4428
rect 38476 3392 38528 3398
rect 38476 3334 38528 3340
rect 38016 3120 38068 3126
rect 38016 3062 38068 3068
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 38304 2938 38332 2994
rect 38212 2910 38332 2938
rect 37832 2372 37884 2378
rect 37832 2314 37884 2320
rect 37844 800 37872 2314
rect 38212 800 38240 2910
rect 38488 800 38516 3334
rect 38672 3058 38700 4422
rect 38844 3936 38896 3942
rect 38844 3878 38896 3884
rect 38660 3052 38712 3058
rect 38660 2994 38712 3000
rect 38856 2378 38884 3878
rect 39132 3534 39160 4558
rect 39856 4480 39908 4486
rect 39856 4422 39908 4428
rect 39868 4321 39896 4422
rect 39854 4312 39910 4321
rect 39854 4247 39910 4256
rect 39394 4176 39450 4185
rect 39394 4111 39450 4120
rect 39120 3528 39172 3534
rect 39120 3470 39172 3476
rect 39408 3126 39436 4111
rect 39764 3936 39816 3942
rect 39764 3878 39816 3884
rect 39488 3392 39540 3398
rect 39488 3334 39540 3340
rect 39396 3120 39448 3126
rect 39396 3062 39448 3068
rect 39120 3052 39172 3058
rect 39120 2994 39172 3000
rect 38844 2372 38896 2378
rect 38844 2314 38896 2320
rect 38856 800 38884 2314
rect 39132 800 39160 2994
rect 39500 800 39528 3334
rect 39776 2446 39804 3878
rect 39868 3534 39896 4247
rect 39948 3936 40000 3942
rect 39948 3878 40000 3884
rect 40408 3936 40460 3942
rect 40408 3878 40460 3884
rect 39856 3528 39908 3534
rect 39856 3470 39908 3476
rect 39960 3058 39988 3878
rect 40222 3224 40278 3233
rect 40222 3159 40278 3168
rect 40236 3126 40264 3159
rect 40224 3120 40276 3126
rect 40224 3062 40276 3068
rect 40420 3058 40448 3878
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 39948 3052 40000 3058
rect 39948 2994 40000 3000
rect 40040 3052 40092 3058
rect 40040 2994 40092 3000
rect 40408 3052 40460 3058
rect 40408 2994 40460 3000
rect 39764 2440 39816 2446
rect 40052 2394 40080 2994
rect 40408 2848 40460 2854
rect 40408 2790 40460 2796
rect 39764 2382 39816 2388
rect 39776 800 39804 2382
rect 39960 2366 40080 2394
rect 39960 1850 39988 2366
rect 40040 2304 40092 2310
rect 40040 2246 40092 2252
rect 40132 2304 40184 2310
rect 40132 2246 40184 2252
rect 40052 1970 40080 2246
rect 40040 1964 40092 1970
rect 40040 1906 40092 1912
rect 39960 1822 40080 1850
rect 40052 800 40080 1822
rect 26608 128 26660 134
rect 26608 70 26660 76
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28078 0 28134 800
rect 28446 0 28502 800
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34702 0 34758 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 36910 0 36966 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 40038 0 40094 800
rect 40144 649 40172 2246
rect 40420 800 40448 2790
rect 40696 2378 40724 3334
rect 40788 3058 40816 4762
rect 41432 3534 41460 5306
rect 41512 4480 41564 4486
rect 41512 4422 41564 4428
rect 41420 3528 41472 3534
rect 41420 3470 41472 3476
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 40776 3052 40828 3058
rect 40776 2994 40828 3000
rect 40684 2372 40736 2378
rect 40684 2314 40736 2320
rect 41052 2372 41104 2378
rect 41052 2314 41104 2320
rect 40696 800 40724 2314
rect 41064 800 41092 2314
rect 41340 800 41368 3334
rect 41524 2378 41552 4422
rect 41708 4146 41736 5510
rect 42260 5302 42288 11591
rect 42340 5568 42392 5574
rect 42340 5510 42392 5516
rect 42248 5296 42300 5302
rect 42248 5238 42300 5244
rect 41696 4140 41748 4146
rect 41696 4082 41748 4088
rect 42352 3534 42380 5510
rect 42536 4758 42564 11727
rect 43258 10976 43314 10985
rect 43258 10911 43314 10920
rect 43074 8936 43130 8945
rect 43074 8871 43130 8880
rect 42984 8628 43036 8634
rect 42984 8570 43036 8576
rect 42708 6860 42760 6866
rect 42708 6802 42760 6808
rect 42720 5710 42748 6802
rect 42800 6180 42852 6186
rect 42800 6122 42852 6128
rect 42708 5704 42760 5710
rect 42708 5646 42760 5652
rect 42616 5024 42668 5030
rect 42616 4966 42668 4972
rect 42524 4752 42576 4758
rect 42524 4694 42576 4700
rect 42340 3528 42392 3534
rect 42340 3470 42392 3476
rect 42248 3392 42300 3398
rect 42248 3334 42300 3340
rect 41972 3052 42024 3058
rect 41972 2994 42024 3000
rect 41696 2848 41748 2854
rect 41696 2790 41748 2796
rect 41512 2372 41564 2378
rect 41512 2314 41564 2320
rect 41604 2304 41656 2310
rect 41604 2246 41656 2252
rect 41616 2106 41644 2246
rect 41604 2100 41656 2106
rect 41604 2042 41656 2048
rect 41708 800 41736 2790
rect 41984 800 42012 2994
rect 42260 800 42288 3334
rect 42628 3058 42656 4966
rect 42812 3126 42840 6122
rect 42996 6118 43024 8570
rect 42984 6112 43036 6118
rect 42984 6054 43036 6060
rect 42892 5568 42944 5574
rect 42892 5510 42944 5516
rect 42904 5234 42932 5510
rect 42892 5228 42944 5234
rect 42892 5170 42944 5176
rect 42984 4548 43036 4554
rect 42984 4490 43036 4496
rect 42996 3466 43024 4490
rect 43088 3670 43116 8871
rect 43168 6112 43220 6118
rect 43168 6054 43220 6060
rect 43180 4622 43208 6054
rect 43168 4616 43220 4622
rect 43168 4558 43220 4564
rect 43168 4480 43220 4486
rect 43168 4422 43220 4428
rect 43076 3664 43128 3670
rect 43076 3606 43128 3612
rect 42984 3460 43036 3466
rect 42984 3402 43036 3408
rect 42800 3120 42852 3126
rect 42800 3062 42852 3068
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 42800 2848 42852 2854
rect 42800 2790 42852 2796
rect 42812 2446 42840 2790
rect 42800 2440 42852 2446
rect 42800 2382 42852 2388
rect 42890 2408 42946 2417
rect 42616 2372 42668 2378
rect 42890 2343 42946 2352
rect 42616 2314 42668 2320
rect 42628 800 42656 2314
rect 42904 2310 42932 2343
rect 42892 2304 42944 2310
rect 42892 2246 42944 2252
rect 42996 2122 43024 3402
rect 43180 3126 43208 4422
rect 43272 4146 43300 10911
rect 43350 10568 43406 10577
rect 43350 10503 43406 10512
rect 43364 10266 43392 10503
rect 43352 10260 43404 10266
rect 43352 10202 43404 10208
rect 43364 10062 43392 10202
rect 43352 10056 43404 10062
rect 43352 9998 43404 10004
rect 43812 6112 43864 6118
rect 43812 6054 43864 6060
rect 43536 5568 43588 5574
rect 43536 5510 43588 5516
rect 43444 5024 43496 5030
rect 43444 4966 43496 4972
rect 43352 4480 43404 4486
rect 43352 4422 43404 4428
rect 43260 4140 43312 4146
rect 43260 4082 43312 4088
rect 43168 3120 43220 3126
rect 43168 3062 43220 3068
rect 43364 2258 43392 4422
rect 43456 2378 43484 4966
rect 43548 4282 43576 5510
rect 43536 4276 43588 4282
rect 43536 4218 43588 4224
rect 43824 4214 43852 6054
rect 43812 4208 43864 4214
rect 43812 4150 43864 4156
rect 43824 3380 43852 4150
rect 43916 3670 43944 17206
rect 44008 4146 44036 18634
rect 44086 10024 44142 10033
rect 44086 9959 44142 9968
rect 44100 9926 44128 9959
rect 44088 9920 44140 9926
rect 44088 9862 44140 9868
rect 44180 6112 44232 6118
rect 44180 6054 44232 6060
rect 44192 4554 44220 6054
rect 45100 5568 45152 5574
rect 45100 5510 45152 5516
rect 44180 4548 44232 4554
rect 44180 4490 44232 4496
rect 44824 4548 44876 4554
rect 44824 4490 44876 4496
rect 43996 4140 44048 4146
rect 43996 4082 44048 4088
rect 44456 4004 44508 4010
rect 44456 3946 44508 3952
rect 44180 3936 44232 3942
rect 44180 3878 44232 3884
rect 43904 3664 43956 3670
rect 43904 3606 43956 3612
rect 43996 3596 44048 3602
rect 43996 3538 44048 3544
rect 43824 3352 43944 3380
rect 43536 3120 43588 3126
rect 43536 3062 43588 3068
rect 43444 2372 43496 2378
rect 43444 2314 43496 2320
rect 42904 2094 43024 2122
rect 43272 2230 43392 2258
rect 42904 800 42932 2094
rect 43272 800 43300 2230
rect 43548 800 43576 3062
rect 43916 800 43944 3352
rect 44008 3194 44036 3538
rect 43996 3188 44048 3194
rect 43996 3130 44048 3136
rect 44192 800 44220 3878
rect 44468 3466 44496 3946
rect 44456 3460 44508 3466
rect 44456 3402 44508 3408
rect 44468 800 44496 3402
rect 44836 800 44864 4490
rect 45112 800 45140 5510
rect 45744 5228 45796 5234
rect 45744 5170 45796 5176
rect 45468 4208 45520 4214
rect 45468 4150 45520 4156
rect 45480 800 45508 4150
rect 45756 800 45784 5170
rect 40130 640 40186 649
rect 40130 575 40186 584
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41326 0 41382 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44454 0 44510 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45742 0 45798 800
<< via2 >>
rect 3974 39616 4030 39672
rect 938 27376 994 27432
rect 18 17040 74 17096
rect 570 21120 626 21176
rect 662 20576 718 20632
rect 846 23432 902 23488
rect 2870 39072 2926 39128
rect 1398 35536 1454 35592
rect 1398 34312 1454 34368
rect 1490 33224 1546 33280
rect 1490 32000 1546 32056
rect 1398 30776 1454 30832
rect 1398 29688 1454 29744
rect 1490 28500 1492 28520
rect 1492 28500 1544 28520
rect 1544 28500 1546 28520
rect 1490 28464 1546 28500
rect 1398 27240 1454 27296
rect 2778 36760 2834 36816
rect 3146 37848 3202 37904
rect 3514 38528 3570 38584
rect 3698 37324 3754 37360
rect 3698 37304 3700 37324
rect 3700 37304 3752 37324
rect 3752 37304 3754 37324
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 3514 34992 3570 35048
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4710 37440 4766 37496
rect 5354 37576 5410 37632
rect 4066 36080 4122 36136
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 3606 33768 3662 33824
rect 3422 32544 3478 32600
rect 1398 26152 1454 26208
rect 1398 24928 1454 24984
rect 1490 23724 1546 23760
rect 1490 23704 1492 23724
rect 1492 23704 1544 23724
rect 1544 23704 1546 23724
rect 1490 22752 1546 22808
rect 1398 22616 1454 22672
rect 1306 16108 1362 16144
rect 1306 16088 1308 16108
rect 1308 16088 1360 16108
rect 1360 16088 1362 16108
rect 1306 14864 1362 14920
rect 1030 14048 1086 14104
rect 846 11736 902 11792
rect 662 5208 718 5264
rect 2042 23432 2098 23488
rect 1950 21664 2006 21720
rect 2410 24556 2412 24576
rect 2412 24556 2464 24576
rect 2464 24556 2466 24576
rect 2410 24520 2466 24556
rect 2410 24012 2412 24032
rect 2412 24012 2464 24032
rect 2464 24012 2466 24032
rect 2410 23976 2466 24012
rect 2042 19216 2098 19272
rect 1766 19080 1822 19136
rect 1674 17196 1730 17232
rect 1674 17176 1676 17196
rect 1676 17176 1728 17196
rect 1728 17176 1730 17196
rect 1674 16244 1730 16280
rect 1674 16224 1676 16244
rect 1676 16224 1728 16244
rect 1728 16224 1730 16244
rect 1582 15988 1584 16008
rect 1584 15988 1636 16008
rect 1636 15988 1638 16008
rect 1582 15952 1638 15988
rect 1674 14456 1730 14512
rect 1122 6296 1178 6352
rect 2042 18808 2098 18864
rect 2134 17060 2190 17096
rect 2134 17040 2136 17060
rect 2136 17040 2188 17060
rect 2188 17040 2190 17060
rect 1766 13640 1822 13696
rect 1674 12688 1730 12744
rect 1582 10668 1638 10704
rect 1582 10648 1584 10668
rect 1584 10648 1636 10668
rect 1636 10648 1638 10668
rect 1582 10532 1638 10568
rect 1582 10512 1584 10532
rect 1584 10512 1636 10532
rect 1636 10512 1638 10532
rect 1490 9560 1546 9616
rect 1398 8880 1454 8936
rect 1858 12316 1860 12336
rect 1860 12316 1912 12336
rect 1912 12316 1914 12336
rect 1858 12280 1914 12316
rect 2134 16360 2190 16416
rect 2134 15408 2190 15464
rect 1858 10240 1914 10296
rect 1950 8744 2006 8800
rect 2870 31456 2926 31512
rect 3514 30232 3570 30288
rect 3422 27920 3478 27976
rect 2870 23860 2926 23896
rect 2870 23840 2872 23860
rect 2872 23840 2924 23860
rect 2924 23840 2926 23860
rect 2962 23432 3018 23488
rect 2594 20984 2650 21040
rect 3054 22072 3110 22128
rect 2870 21392 2926 21448
rect 2870 20848 2926 20904
rect 2778 20304 2834 20360
rect 2318 13932 2374 13968
rect 2318 13912 2320 13932
rect 2320 13912 2372 13932
rect 2372 13912 2374 13932
rect 2686 18128 2742 18184
rect 2962 17856 3018 17912
rect 4986 35944 5042 36000
rect 4710 34584 4766 34640
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 3882 29008 3938 29064
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 26696 4122 26752
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4158 24676 4214 24712
rect 4158 24656 4160 24676
rect 4160 24656 4212 24676
rect 4212 24656 4214 24676
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4066 24384 4122 24440
rect 4066 23432 4122 23488
rect 4710 23432 4766 23488
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 3974 22888 4030 22944
rect 3238 19760 3294 19816
rect 3330 19660 3332 19680
rect 3332 19660 3384 19680
rect 3384 19660 3386 19680
rect 3330 19624 3386 19660
rect 3422 19216 3478 19272
rect 3146 18400 3202 18456
rect 2686 16496 2742 16552
rect 2778 13912 2834 13968
rect 2870 13776 2926 13832
rect 2134 10104 2190 10160
rect 2410 11872 2466 11928
rect 1766 8472 1822 8528
rect 2042 8336 2098 8392
rect 1398 7248 1454 7304
rect 1490 6160 1546 6216
rect 1490 4936 1546 4992
rect 2226 8608 2282 8664
rect 3238 17176 3294 17232
rect 3238 16632 3294 16688
rect 3606 21800 3662 21856
rect 3514 16768 3570 16824
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 3698 20168 3754 20224
rect 3698 20032 3754 20088
rect 3882 21120 3938 21176
rect 3882 20984 3938 21040
rect 3698 18536 3754 18592
rect 3698 17992 3754 18048
rect 3974 18284 4030 18320
rect 3974 18264 3976 18284
rect 3976 18264 4028 18284
rect 4028 18264 4030 18284
rect 8114 37340 8116 37360
rect 8116 37340 8168 37360
rect 8168 37340 8170 37360
rect 8114 37304 8170 37340
rect 4986 23840 5042 23896
rect 4894 23160 4950 23216
rect 4802 21528 4858 21584
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4250 20984 4306 21040
rect 4342 20868 4398 20904
rect 4342 20848 4344 20868
rect 4344 20848 4396 20868
rect 4396 20848 4398 20868
rect 4526 20340 4528 20360
rect 4528 20340 4580 20360
rect 4580 20340 4582 20360
rect 4526 20304 4582 20340
rect 4618 20168 4674 20224
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4250 19896 4306 19952
rect 4526 19352 4582 19408
rect 4710 19352 4766 19408
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4526 18808 4582 18864
rect 4158 18536 4214 18592
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4066 17312 4122 17368
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 5170 23432 5226 23488
rect 5170 22208 5226 22264
rect 5354 21664 5410 21720
rect 5630 23588 5686 23624
rect 5630 23568 5632 23588
rect 5632 23568 5684 23588
rect 5684 23568 5686 23588
rect 5538 23196 5540 23216
rect 5540 23196 5592 23216
rect 5592 23196 5594 23216
rect 5538 23160 5594 23196
rect 5446 21392 5502 21448
rect 4986 17448 5042 17504
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 3606 15544 3662 15600
rect 4618 15564 4674 15600
rect 4618 15544 4620 15564
rect 4620 15544 4672 15564
rect 4672 15544 4674 15564
rect 4066 15000 4122 15056
rect 4710 15408 4766 15464
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 3422 14320 3478 14376
rect 3146 12008 3202 12064
rect 2870 11328 2926 11384
rect 2594 10140 2596 10160
rect 2596 10140 2648 10160
rect 2648 10140 2650 10160
rect 2594 10104 2650 10140
rect 2594 8200 2650 8256
rect 2686 8064 2742 8120
rect 2042 4664 2098 4720
rect 938 2488 994 2544
rect 1398 3712 1454 3768
rect 2870 9696 2926 9752
rect 3146 10784 3202 10840
rect 3882 14220 3884 14240
rect 3884 14220 3936 14240
rect 3936 14220 3938 14240
rect 3882 14184 3938 14220
rect 4342 14492 4344 14512
rect 4344 14492 4396 14512
rect 4396 14492 4398 14512
rect 4342 14456 4398 14492
rect 5446 20848 5502 20904
rect 5354 19624 5410 19680
rect 5354 19352 5410 19408
rect 5538 20712 5594 20768
rect 5538 20576 5594 20632
rect 6182 22752 6238 22808
rect 6274 22480 6330 22536
rect 5814 20460 5870 20496
rect 5814 20440 5816 20460
rect 5816 20440 5868 20460
rect 5868 20440 5870 20460
rect 5446 18808 5502 18864
rect 5354 17992 5410 18048
rect 4066 14320 4122 14376
rect 3882 13388 3938 13424
rect 3882 13368 3884 13388
rect 3884 13368 3936 13388
rect 3936 13368 3938 13388
rect 3882 13232 3938 13288
rect 3514 13096 3570 13152
rect 3514 12980 3570 13016
rect 3514 12960 3516 12980
rect 3516 12960 3568 12980
rect 3568 12960 3570 12980
rect 3514 12688 3570 12744
rect 3790 12552 3846 12608
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4158 13096 4214 13152
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3790 11464 3846 11520
rect 3974 11600 4030 11656
rect 4526 12144 4582 12200
rect 3606 9968 3662 10024
rect 3606 9716 3662 9752
rect 3606 9696 3608 9716
rect 3608 9696 3660 9716
rect 3660 9696 3662 9716
rect 3514 9444 3570 9480
rect 3514 9424 3516 9444
rect 3516 9424 3568 9444
rect 3568 9424 3570 9444
rect 3054 2624 3110 2680
rect 3054 2080 3110 2136
rect 2962 1536 3018 1592
rect 2870 1400 2926 1456
rect 2778 856 2834 912
rect 3422 8628 3478 8664
rect 3422 8608 3424 8628
rect 3424 8608 3476 8628
rect 3476 8608 3478 8628
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4158 10784 4214 10840
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4710 11056 4766 11112
rect 3882 9696 3938 9752
rect 3882 9560 3938 9616
rect 4526 9560 4582 9616
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 5262 13776 5318 13832
rect 5538 17720 5594 17776
rect 6090 19352 6146 19408
rect 5998 17992 6054 18048
rect 6642 23568 6698 23624
rect 6550 23432 6606 23488
rect 6642 21800 6698 21856
rect 6642 20304 6698 20360
rect 6550 20032 6606 20088
rect 7378 27104 7434 27160
rect 6918 26832 6974 26888
rect 6918 26152 6974 26208
rect 6826 20712 6882 20768
rect 5538 16904 5594 16960
rect 5538 14456 5594 14512
rect 4986 12416 5042 12472
rect 5538 13640 5594 13696
rect 5814 14184 5870 14240
rect 5906 12824 5962 12880
rect 4986 11620 5042 11656
rect 4986 11600 4988 11620
rect 4988 11600 5040 11620
rect 5040 11600 5042 11620
rect 4894 11328 4950 11384
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4342 7792 4398 7848
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4618 6976 4674 7032
rect 3882 6452 3938 6488
rect 4434 6860 4490 6896
rect 4434 6840 4436 6860
rect 4436 6840 4488 6860
rect 4488 6840 4490 6860
rect 4618 6704 4674 6760
rect 3882 6432 3884 6452
rect 3884 6432 3936 6452
rect 3936 6432 3938 6452
rect 3330 6160 3386 6216
rect 3146 856 3202 912
rect 3422 3052 3478 3088
rect 3422 3032 3424 3052
rect 3424 3032 3476 3052
rect 3476 3032 3478 3052
rect 3330 1264 3386 1320
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 3974 5480 4030 5536
rect 4066 5344 4122 5400
rect 4618 5480 4674 5536
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4066 4392 4122 4448
rect 5722 11892 5778 11928
rect 5722 11872 5724 11892
rect 5724 11872 5776 11892
rect 5776 11872 5778 11892
rect 5538 9560 5594 9616
rect 5354 9324 5356 9344
rect 5356 9324 5408 9344
rect 5408 9324 5410 9344
rect 5354 9288 5410 9324
rect 5078 7248 5134 7304
rect 5170 6860 5226 6896
rect 5170 6840 5172 6860
rect 5172 6840 5224 6860
rect 5224 6840 5226 6860
rect 5078 6704 5134 6760
rect 4986 5888 5042 5944
rect 4894 4936 4950 4992
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3974 3612 3976 3632
rect 3976 3612 4028 3632
rect 4028 3612 4030 3632
rect 4710 3848 4766 3904
rect 3974 3576 4030 3612
rect 3882 3168 3938 3224
rect 4066 3188 4122 3224
rect 4066 3168 4068 3188
rect 4068 3168 4120 3188
rect 4120 3168 4122 3188
rect 4618 3440 4674 3496
rect 938 312 994 368
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4066 1944 4122 2000
rect 4618 1128 4674 1184
rect 4250 40 4306 96
rect 5170 2760 5226 2816
rect 5354 6704 5410 6760
rect 6274 16768 6330 16824
rect 6550 18536 6606 18592
rect 6734 17740 6790 17776
rect 6734 17720 6736 17740
rect 6736 17720 6788 17740
rect 6788 17720 6790 17740
rect 7010 20712 7066 20768
rect 6734 15952 6790 16008
rect 6458 15272 6514 15328
rect 6458 14456 6514 14512
rect 6734 14320 6790 14376
rect 6550 13640 6606 13696
rect 5998 11192 6054 11248
rect 6274 12144 6330 12200
rect 6550 12008 6606 12064
rect 6550 11736 6606 11792
rect 6274 11328 6330 11384
rect 6366 10920 6422 10976
rect 6274 10784 6330 10840
rect 6458 10784 6514 10840
rect 6090 9560 6146 9616
rect 6090 9152 6146 9208
rect 5814 6568 5870 6624
rect 5538 4528 5594 4584
rect 6182 8900 6238 8936
rect 6182 8880 6184 8900
rect 6184 8880 6236 8900
rect 6236 8880 6238 8900
rect 6182 8336 6238 8392
rect 6642 11076 6698 11112
rect 6642 11056 6644 11076
rect 6644 11056 6696 11076
rect 6696 11056 6698 11076
rect 6642 9152 6698 9208
rect 7194 22072 7250 22128
rect 7194 19760 7250 19816
rect 7286 18672 7342 18728
rect 7102 17856 7158 17912
rect 7194 16496 7250 16552
rect 6366 6976 6422 7032
rect 6550 7656 6606 7712
rect 7194 12144 7250 12200
rect 7378 16632 7434 16688
rect 7930 23432 7986 23488
rect 7654 20304 7710 20360
rect 7562 18128 7618 18184
rect 7562 17312 7618 17368
rect 7562 16632 7618 16688
rect 8574 26732 8576 26752
rect 8576 26732 8628 26752
rect 8628 26732 8630 26752
rect 8574 26696 8630 26732
rect 7930 21972 7932 21992
rect 7932 21972 7984 21992
rect 7984 21972 7986 21992
rect 7930 21936 7986 21972
rect 8298 23976 8354 24032
rect 8666 24792 8722 24848
rect 8114 20576 8170 20632
rect 8022 16904 8078 16960
rect 7378 12824 7434 12880
rect 6918 9968 6974 10024
rect 6918 9560 6974 9616
rect 7010 9016 7066 9072
rect 7102 8880 7158 8936
rect 8390 20032 8446 20088
rect 8758 23160 8814 23216
rect 8574 19896 8630 19952
rect 9218 24112 9274 24168
rect 9034 22888 9090 22944
rect 9034 21800 9090 21856
rect 8942 20440 8998 20496
rect 8666 19624 8722 19680
rect 8666 18672 8722 18728
rect 8574 18128 8630 18184
rect 8390 15272 8446 15328
rect 8206 15036 8208 15056
rect 8208 15036 8260 15056
rect 8260 15036 8262 15056
rect 8206 15000 8262 15036
rect 8114 14864 8170 14920
rect 7746 14456 7802 14512
rect 7654 11328 7710 11384
rect 7930 12960 7986 13016
rect 7838 11600 7894 11656
rect 8574 12416 8630 12472
rect 8206 10784 8262 10840
rect 8022 10240 8078 10296
rect 8022 9968 8078 10024
rect 8022 9560 8078 9616
rect 7746 9152 7802 9208
rect 7378 8880 7434 8936
rect 6642 7112 6698 7168
rect 6734 3304 6790 3360
rect 6550 1808 6606 1864
rect 7194 7928 7250 7984
rect 8114 9152 8170 9208
rect 7746 8744 7802 8800
rect 7654 7248 7710 7304
rect 7470 6704 7526 6760
rect 7470 6432 7526 6488
rect 7010 2624 7066 2680
rect 8942 18400 8998 18456
rect 9494 28872 9550 28928
rect 9494 26460 9496 26480
rect 9496 26460 9548 26480
rect 9548 26460 9550 26480
rect 9494 26424 9550 26460
rect 9678 22480 9734 22536
rect 9954 24556 9956 24576
rect 9956 24556 10008 24576
rect 10008 24556 10010 24576
rect 9954 24520 10010 24556
rect 10046 24248 10102 24304
rect 10138 23976 10194 24032
rect 10046 23704 10102 23760
rect 9770 21120 9826 21176
rect 9402 19488 9458 19544
rect 9034 16496 9090 16552
rect 8758 12280 8814 12336
rect 8482 9152 8538 9208
rect 8666 9152 8722 9208
rect 8942 12552 8998 12608
rect 9126 15952 9182 16008
rect 9218 15680 9274 15736
rect 9218 14592 9274 14648
rect 9678 19624 9734 19680
rect 9402 15136 9458 15192
rect 8942 10260 8998 10296
rect 8942 10240 8944 10260
rect 8944 10240 8996 10260
rect 8996 10240 8998 10260
rect 9310 10784 9366 10840
rect 9126 10512 9182 10568
rect 9034 9988 9090 10024
rect 9034 9968 9036 9988
rect 9036 9968 9088 9988
rect 9088 9968 9090 9988
rect 8942 9832 8998 9888
rect 9218 9832 9274 9888
rect 8850 9288 8906 9344
rect 8206 6976 8262 7032
rect 8298 6704 8354 6760
rect 9126 9288 9182 9344
rect 9494 11736 9550 11792
rect 9402 9288 9458 9344
rect 8942 7792 8998 7848
rect 8850 7656 8906 7712
rect 9034 7656 9090 7712
rect 8574 6024 8630 6080
rect 10874 32408 10930 32464
rect 10414 27648 10470 27704
rect 10598 24812 10654 24848
rect 10598 24792 10600 24812
rect 10600 24792 10652 24812
rect 10652 24792 10654 24812
rect 10414 23840 10470 23896
rect 10506 23432 10562 23488
rect 10230 22888 10286 22944
rect 10414 22652 10416 22672
rect 10416 22652 10468 22672
rect 10468 22652 10470 22672
rect 10414 22616 10470 22652
rect 10322 22480 10378 22536
rect 10138 22208 10194 22264
rect 10230 22072 10286 22128
rect 10322 21936 10378 21992
rect 10966 24656 11022 24712
rect 10782 22636 10838 22672
rect 10782 22616 10784 22636
rect 10784 22616 10836 22636
rect 10836 22616 10838 22636
rect 10782 22072 10838 22128
rect 10138 17584 10194 17640
rect 10322 19488 10378 19544
rect 10230 16632 10286 16688
rect 9862 13812 9864 13832
rect 9864 13812 9916 13832
rect 9916 13812 9918 13832
rect 9862 13776 9918 13812
rect 9678 13368 9734 13424
rect 9862 12416 9918 12472
rect 9770 11056 9826 11112
rect 9494 7928 9550 7984
rect 9494 7656 9550 7712
rect 9586 7520 9642 7576
rect 9494 6976 9550 7032
rect 9126 4820 9182 4856
rect 9126 4800 9128 4820
rect 9128 4800 9180 4820
rect 9180 4800 9182 4820
rect 8942 4392 8998 4448
rect 9402 6860 9458 6896
rect 9402 6840 9404 6860
rect 9404 6840 9456 6860
rect 9456 6840 9458 6860
rect 9310 6160 9366 6216
rect 9402 5908 9458 5944
rect 9402 5888 9404 5908
rect 9404 5888 9456 5908
rect 9456 5888 9458 5908
rect 9586 6704 9642 6760
rect 9586 6160 9642 6216
rect 9494 3732 9550 3768
rect 9494 3712 9496 3732
rect 9496 3712 9548 3732
rect 9548 3712 9550 3732
rect 9770 6316 9826 6352
rect 9770 6296 9772 6316
rect 9772 6296 9824 6316
rect 9824 6296 9826 6316
rect 9678 5480 9734 5536
rect 9954 11192 10010 11248
rect 9954 9832 10010 9888
rect 9954 8472 10010 8528
rect 9954 8200 10010 8256
rect 9954 8084 10010 8120
rect 9954 8064 9956 8084
rect 9956 8064 10008 8084
rect 10008 8064 10010 8084
rect 9954 6568 10010 6624
rect 10782 21392 10838 21448
rect 10782 20440 10838 20496
rect 10690 19760 10746 19816
rect 10690 19488 10746 19544
rect 10690 19352 10746 19408
rect 10322 13640 10378 13696
rect 10690 16768 10746 16824
rect 10598 12960 10654 13016
rect 10506 12280 10562 12336
rect 10230 10512 10286 10568
rect 10322 9696 10378 9752
rect 10138 9016 10194 9072
rect 11058 22072 11114 22128
rect 10966 18536 11022 18592
rect 11518 25644 11520 25664
rect 11520 25644 11572 25664
rect 11572 25644 11574 25664
rect 11518 25608 11574 25644
rect 11426 25064 11482 25120
rect 11518 24928 11574 24984
rect 11334 22616 11390 22672
rect 11334 18808 11390 18864
rect 11610 23296 11666 23352
rect 12162 23296 12218 23352
rect 11886 21836 11888 21856
rect 11888 21836 11940 21856
rect 11940 21836 11942 21856
rect 11886 21800 11942 21836
rect 11702 21528 11758 21584
rect 11334 17856 11390 17912
rect 10874 16496 10930 16552
rect 10874 15680 10930 15736
rect 10782 14456 10838 14512
rect 10782 13912 10838 13968
rect 11150 17040 11206 17096
rect 11334 16360 11390 16416
rect 11702 18536 11758 18592
rect 11610 16244 11666 16280
rect 11610 16224 11612 16244
rect 11612 16224 11664 16244
rect 11664 16224 11666 16244
rect 11702 15136 11758 15192
rect 11610 14884 11666 14920
rect 11610 14864 11612 14884
rect 11612 14864 11664 14884
rect 11664 14864 11666 14884
rect 11058 14048 11114 14104
rect 10874 12824 10930 12880
rect 10782 10648 10838 10704
rect 10230 6160 10286 6216
rect 10230 5652 10232 5672
rect 10232 5652 10284 5672
rect 10284 5652 10286 5672
rect 10230 5616 10286 5652
rect 11058 10240 11114 10296
rect 11518 14184 11574 14240
rect 11426 12416 11482 12472
rect 11334 11872 11390 11928
rect 11426 11192 11482 11248
rect 11334 11056 11390 11112
rect 11150 10104 11206 10160
rect 10874 8608 10930 8664
rect 11058 8608 11114 8664
rect 10506 6976 10562 7032
rect 10874 8472 10930 8528
rect 10782 7384 10838 7440
rect 10506 6704 10562 6760
rect 10598 6568 10654 6624
rect 10598 5652 10600 5672
rect 10600 5652 10652 5672
rect 10652 5652 10654 5672
rect 10598 5616 10654 5652
rect 10138 4528 10194 4584
rect 10782 5108 10784 5128
rect 10784 5108 10836 5128
rect 10836 5108 10838 5128
rect 10782 5072 10838 5108
rect 10782 4528 10838 4584
rect 10506 4120 10562 4176
rect 9770 2488 9826 2544
rect 6182 176 6238 232
rect 9586 2216 9642 2272
rect 10138 2508 10194 2544
rect 10138 2488 10140 2508
rect 10140 2488 10192 2508
rect 10192 2488 10194 2508
rect 11150 7112 11206 7168
rect 11058 5888 11114 5944
rect 10966 5480 11022 5536
rect 11150 5208 11206 5264
rect 11518 9832 11574 9888
rect 11610 9560 11666 9616
rect 12714 26968 12770 27024
rect 12622 26460 12624 26480
rect 12624 26460 12676 26480
rect 12676 26460 12678 26480
rect 12622 26424 12678 26460
rect 12714 25880 12770 25936
rect 12530 25608 12586 25664
rect 12346 23468 12348 23488
rect 12348 23468 12400 23488
rect 12400 23468 12402 23488
rect 12346 23432 12402 23468
rect 12530 25200 12586 25256
rect 12346 22888 12402 22944
rect 12530 22888 12586 22944
rect 12438 22072 12494 22128
rect 12070 20712 12126 20768
rect 12162 18808 12218 18864
rect 12898 23588 12954 23624
rect 12898 23568 12900 23588
rect 12900 23568 12952 23588
rect 12952 23568 12954 23588
rect 12898 21936 12954 21992
rect 12530 20712 12586 20768
rect 12438 17740 12494 17776
rect 12438 17720 12440 17740
rect 12440 17720 12492 17740
rect 12492 17720 12494 17740
rect 11886 11464 11942 11520
rect 11886 9968 11942 10024
rect 11794 9424 11850 9480
rect 11978 9696 12034 9752
rect 11978 9560 12034 9616
rect 11426 7692 11428 7712
rect 11428 7692 11480 7712
rect 11480 7692 11482 7712
rect 11426 7656 11482 7692
rect 11518 7520 11574 7576
rect 11426 7148 11428 7168
rect 11428 7148 11480 7168
rect 11480 7148 11482 7168
rect 11426 7112 11482 7148
rect 11334 5752 11390 5808
rect 11150 3168 11206 3224
rect 11610 7268 11666 7304
rect 11610 7248 11612 7268
rect 11612 7248 11664 7268
rect 11664 7248 11666 7268
rect 11610 7112 11666 7168
rect 12806 19624 12862 19680
rect 12806 16496 12862 16552
rect 13174 30504 13230 30560
rect 13082 26308 13138 26344
rect 13082 26288 13084 26308
rect 13084 26288 13136 26308
rect 13136 26288 13138 26308
rect 13082 25200 13138 25256
rect 13174 22480 13230 22536
rect 13082 22344 13138 22400
rect 12990 19624 13046 19680
rect 13174 21684 13230 21720
rect 13174 21664 13176 21684
rect 13176 21664 13228 21684
rect 13228 21664 13230 21684
rect 13174 21412 13230 21448
rect 13174 21392 13176 21412
rect 13176 21392 13228 21412
rect 13228 21392 13230 21412
rect 13174 21256 13230 21312
rect 14370 35944 14426 36000
rect 13726 34584 13782 34640
rect 13358 30368 13414 30424
rect 13726 26288 13782 26344
rect 13634 24284 13636 24304
rect 13636 24284 13688 24304
rect 13688 24284 13690 24304
rect 13634 24248 13690 24284
rect 13542 23568 13598 23624
rect 13450 22752 13506 22808
rect 13450 21664 13506 21720
rect 13358 19352 13414 19408
rect 13174 17992 13230 18048
rect 13174 16652 13230 16688
rect 13174 16632 13176 16652
rect 13176 16632 13228 16652
rect 13228 16632 13230 16652
rect 13174 16396 13176 16416
rect 13176 16396 13228 16416
rect 13228 16396 13230 16416
rect 13174 16360 13230 16396
rect 12622 14492 12624 14512
rect 12624 14492 12676 14512
rect 12676 14492 12678 14512
rect 12622 14456 12678 14492
rect 12254 13504 12310 13560
rect 12346 13096 12402 13152
rect 11886 6976 11942 7032
rect 11886 6704 11942 6760
rect 11794 5616 11850 5672
rect 11794 3304 11850 3360
rect 12438 10512 12494 10568
rect 12438 10104 12494 10160
rect 12346 8372 12348 8392
rect 12348 8372 12400 8392
rect 12400 8372 12402 8392
rect 12346 8336 12402 8372
rect 12346 7928 12402 7984
rect 12254 5752 12310 5808
rect 12162 5208 12218 5264
rect 12162 4800 12218 4856
rect 12438 4256 12494 4312
rect 11610 720 11666 776
rect 12806 13640 12862 13696
rect 12806 13096 12862 13152
rect 13174 14612 13230 14648
rect 13910 22480 13966 22536
rect 13542 19896 13598 19952
rect 13542 19796 13544 19816
rect 13544 19796 13596 19816
rect 13596 19796 13598 19816
rect 13542 19760 13598 19796
rect 13634 19352 13690 19408
rect 13450 19216 13506 19272
rect 13358 17992 13414 18048
rect 13450 15272 13506 15328
rect 13174 14592 13176 14612
rect 13176 14592 13228 14612
rect 13228 14592 13230 14612
rect 13082 14456 13138 14512
rect 12990 13640 13046 13696
rect 12622 9152 12678 9208
rect 12898 12960 12954 13016
rect 12990 12416 13046 12472
rect 12898 11212 12954 11248
rect 12898 11192 12900 11212
rect 12900 11192 12952 11212
rect 12952 11192 12954 11212
rect 12990 9968 13046 10024
rect 12898 9288 12954 9344
rect 13174 14184 13230 14240
rect 13358 13776 13414 13832
rect 13542 13776 13598 13832
rect 13358 11892 13414 11928
rect 13358 11872 13360 11892
rect 13360 11872 13412 11892
rect 13412 11872 13414 11892
rect 13174 10920 13230 10976
rect 13174 10104 13230 10160
rect 13542 10512 13598 10568
rect 13910 14456 13966 14512
rect 14278 23860 14334 23896
rect 14278 23840 14280 23860
rect 14280 23840 14332 23860
rect 14332 23840 14334 23860
rect 14094 21528 14150 21584
rect 14094 19352 14150 19408
rect 14094 18808 14150 18864
rect 14370 21140 14426 21176
rect 14370 21120 14372 21140
rect 14372 21120 14424 21140
rect 14424 21120 14426 21140
rect 14370 20576 14426 20632
rect 14278 19080 14334 19136
rect 14922 24928 14978 24984
rect 14554 21936 14610 21992
rect 14646 21528 14702 21584
rect 14554 17448 14610 17504
rect 14278 17312 14334 17368
rect 14370 16360 14426 16416
rect 14186 15680 14242 15736
rect 14462 15700 14518 15736
rect 14462 15680 14464 15700
rect 14464 15680 14516 15700
rect 14516 15680 14518 15700
rect 14094 12552 14150 12608
rect 14002 11192 14058 11248
rect 14002 10532 14058 10568
rect 14002 10512 14004 10532
rect 14004 10512 14056 10532
rect 14056 10512 14058 10532
rect 13634 9832 13690 9888
rect 13174 7792 13230 7848
rect 12438 1536 12494 1592
rect 13082 6840 13138 6896
rect 13726 8608 13782 8664
rect 13542 6024 13598 6080
rect 13726 6432 13782 6488
rect 13726 5208 13782 5264
rect 13818 4392 13874 4448
rect 14370 14048 14426 14104
rect 14278 11464 14334 11520
rect 14278 10376 14334 10432
rect 14830 22208 14886 22264
rect 15014 20576 15070 20632
rect 15198 25336 15254 25392
rect 15290 24792 15346 24848
rect 15290 24520 15346 24576
rect 15198 20576 15254 20632
rect 15198 18808 15254 18864
rect 15106 15816 15162 15872
rect 14646 13504 14702 13560
rect 14830 11192 14886 11248
rect 14554 10512 14610 10568
rect 14462 10104 14518 10160
rect 14462 9832 14518 9888
rect 14094 8608 14150 8664
rect 14002 8336 14058 8392
rect 14094 8200 14150 8256
rect 13726 2896 13782 2952
rect 14094 7112 14150 7168
rect 14186 6180 14242 6216
rect 14186 6160 14188 6180
rect 14188 6160 14240 6180
rect 14240 6160 14242 6180
rect 14186 4428 14188 4448
rect 14188 4428 14240 4448
rect 14240 4428 14242 4448
rect 14186 4392 14242 4428
rect 14370 8336 14426 8392
rect 14462 7540 14518 7576
rect 14462 7520 14464 7540
rect 14464 7520 14516 7540
rect 14516 7520 14518 7540
rect 14370 5636 14426 5672
rect 14370 5616 14372 5636
rect 14372 5616 14424 5636
rect 14424 5616 14426 5636
rect 14186 3984 14242 4040
rect 14370 3188 14426 3224
rect 15290 13776 15346 13832
rect 15198 13252 15254 13288
rect 15198 13232 15200 13252
rect 15200 13232 15252 13252
rect 15252 13232 15254 13252
rect 15014 12416 15070 12472
rect 15290 12844 15346 12880
rect 15290 12824 15292 12844
rect 15292 12824 15344 12844
rect 15344 12824 15346 12844
rect 15014 10956 15016 10976
rect 15016 10956 15068 10976
rect 15068 10956 15070 10976
rect 15014 10920 15070 10956
rect 15106 10784 15162 10840
rect 15014 10376 15070 10432
rect 15290 10648 15346 10704
rect 14922 9444 14978 9480
rect 14922 9424 14924 9444
rect 14924 9424 14976 9444
rect 14976 9424 14978 9444
rect 15014 8200 15070 8256
rect 15014 7248 15070 7304
rect 15290 8336 15346 8392
rect 15474 16224 15530 16280
rect 15750 24792 15806 24848
rect 15842 22772 15898 22808
rect 15842 22752 15844 22772
rect 15844 22752 15896 22772
rect 15896 22752 15898 22772
rect 15842 22208 15898 22264
rect 15658 19896 15714 19952
rect 15658 19080 15714 19136
rect 15842 21140 15898 21176
rect 15842 21120 15844 21140
rect 15844 21120 15896 21140
rect 15896 21120 15898 21140
rect 16210 22752 16266 22808
rect 16210 22344 16266 22400
rect 16302 22208 16358 22264
rect 16210 19916 16266 19952
rect 16210 19896 16212 19916
rect 16212 19896 16264 19916
rect 16264 19896 16266 19916
rect 16118 19624 16174 19680
rect 15934 19216 15990 19272
rect 16026 18264 16082 18320
rect 16026 17584 16082 17640
rect 16026 16632 16082 16688
rect 15934 16088 15990 16144
rect 15750 14048 15806 14104
rect 15842 13504 15898 13560
rect 15750 13232 15806 13288
rect 15290 7656 15346 7712
rect 15566 11756 15622 11792
rect 15566 11736 15568 11756
rect 15568 11736 15620 11756
rect 15620 11736 15622 11756
rect 15750 11464 15806 11520
rect 16118 16224 16174 16280
rect 17038 36488 17094 36544
rect 16854 23432 16910 23488
rect 16854 21972 16856 21992
rect 16856 21972 16908 21992
rect 16908 21972 16910 21992
rect 16854 21936 16910 21972
rect 16670 20712 16726 20768
rect 16578 20440 16634 20496
rect 16486 20304 16542 20360
rect 16670 20032 16726 20088
rect 16486 19624 16542 19680
rect 16394 16768 16450 16824
rect 16302 16632 16358 16688
rect 16670 18572 16672 18592
rect 16672 18572 16724 18592
rect 16724 18572 16726 18592
rect 16670 18536 16726 18572
rect 16670 17992 16726 18048
rect 16670 17196 16726 17232
rect 16670 17176 16672 17196
rect 16672 17176 16724 17196
rect 16724 17176 16726 17196
rect 16670 16496 16726 16552
rect 16394 16360 16450 16416
rect 16210 15680 16266 15736
rect 16210 14864 16266 14920
rect 16118 14728 16174 14784
rect 16486 15852 16488 15872
rect 16488 15852 16540 15872
rect 16540 15852 16542 15872
rect 16486 15816 16542 15852
rect 16394 13776 16450 13832
rect 16210 12552 16266 12608
rect 16026 11736 16082 11792
rect 15934 9968 15990 10024
rect 15750 9580 15806 9616
rect 15750 9560 15752 9580
rect 15752 9560 15804 9580
rect 15804 9560 15806 9580
rect 15658 9424 15714 9480
rect 15566 8236 15568 8256
rect 15568 8236 15620 8256
rect 15620 8236 15622 8256
rect 15566 8200 15622 8236
rect 15382 6840 15438 6896
rect 15106 6332 15108 6352
rect 15108 6332 15160 6352
rect 15160 6332 15162 6352
rect 15106 6296 15162 6332
rect 15382 6196 15384 6216
rect 15384 6196 15436 6216
rect 15436 6196 15438 6216
rect 15382 6160 15438 6196
rect 15382 4020 15384 4040
rect 15384 4020 15436 4040
rect 15436 4020 15438 4040
rect 15382 3984 15438 4020
rect 15198 3712 15254 3768
rect 15106 3304 15162 3360
rect 14370 3168 14372 3188
rect 14372 3168 14424 3188
rect 14424 3168 14426 3188
rect 16118 9968 16174 10024
rect 16762 11192 16818 11248
rect 16670 11056 16726 11112
rect 16394 10920 16450 10976
rect 16118 7792 16174 7848
rect 15658 6296 15714 6352
rect 15842 3984 15898 4040
rect 15842 3576 15898 3632
rect 15934 3440 15990 3496
rect 16302 7828 16304 7848
rect 16304 7828 16356 7848
rect 16356 7828 16358 7848
rect 16302 7792 16358 7828
rect 16302 7112 16358 7168
rect 16762 10512 16818 10568
rect 16670 10240 16726 10296
rect 17406 21836 17408 21856
rect 17408 21836 17460 21856
rect 17460 21836 17462 21856
rect 17406 21800 17462 21836
rect 17130 19760 17186 19816
rect 16946 17176 17002 17232
rect 17222 19624 17278 19680
rect 17222 19216 17278 19272
rect 17130 18400 17186 18456
rect 17774 36488 17830 36544
rect 17866 23432 17922 23488
rect 17222 18264 17278 18320
rect 17130 17876 17186 17912
rect 17130 17856 17132 17876
rect 17132 17856 17184 17876
rect 17184 17856 17186 17876
rect 17498 17992 17554 18048
rect 17498 17620 17500 17640
rect 17500 17620 17552 17640
rect 17552 17620 17554 17640
rect 17498 17584 17554 17620
rect 17406 17312 17462 17368
rect 18050 23840 18106 23896
rect 18050 23196 18052 23216
rect 18052 23196 18104 23216
rect 18104 23196 18106 23216
rect 18050 23160 18106 23196
rect 18326 34584 18382 34640
rect 18142 22344 18198 22400
rect 18050 21020 18052 21040
rect 18052 21020 18104 21040
rect 18104 21020 18106 21040
rect 18050 20984 18106 21020
rect 18510 26016 18566 26072
rect 18510 23432 18566 23488
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19890 36080 19946 36136
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19430 35264 19486 35320
rect 19246 24792 19302 24848
rect 18694 23432 18750 23488
rect 18510 23160 18566 23216
rect 18510 22752 18566 22808
rect 18142 20848 18198 20904
rect 17774 18400 17830 18456
rect 16946 12164 17002 12200
rect 16946 12144 16948 12164
rect 16948 12144 17000 12164
rect 17000 12144 17002 12164
rect 16854 10240 16910 10296
rect 16762 9832 16818 9888
rect 16670 9696 16726 9752
rect 17038 11328 17094 11384
rect 17222 12688 17278 12744
rect 17406 15308 17408 15328
rect 17408 15308 17460 15328
rect 17460 15308 17462 15328
rect 17406 15272 17462 15308
rect 17498 12844 17554 12880
rect 17498 12824 17500 12844
rect 17500 12824 17552 12844
rect 17552 12824 17554 12844
rect 18326 21256 18382 21312
rect 18418 20712 18474 20768
rect 19338 23568 19394 23624
rect 19246 22924 19248 22944
rect 19248 22924 19300 22944
rect 19300 22924 19302 22944
rect 19246 22888 19302 22924
rect 19338 22480 19394 22536
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19890 22616 19946 22672
rect 19246 21800 19302 21856
rect 18970 20596 19026 20632
rect 18970 20576 18972 20596
rect 18972 20576 19024 20596
rect 19024 20576 19026 20596
rect 18142 19760 18198 19816
rect 18142 19216 18198 19272
rect 18050 18536 18106 18592
rect 18142 18028 18144 18048
rect 18144 18028 18196 18048
rect 18196 18028 18198 18048
rect 18142 17992 18198 18028
rect 18326 17992 18382 18048
rect 18142 17856 18198 17912
rect 18050 17720 18106 17776
rect 17682 15680 17738 15736
rect 17314 12316 17316 12336
rect 17316 12316 17368 12336
rect 17368 12316 17370 12336
rect 17314 12280 17370 12316
rect 17590 12280 17646 12336
rect 17498 12008 17554 12064
rect 17406 11736 17462 11792
rect 16946 9560 17002 9616
rect 17222 10784 17278 10840
rect 17222 9988 17278 10024
rect 17222 9968 17224 9988
rect 17224 9968 17276 9988
rect 17276 9968 17278 9988
rect 16486 9172 16542 9208
rect 16486 9152 16488 9172
rect 16488 9152 16540 9172
rect 16540 9152 16542 9172
rect 16762 9152 16818 9208
rect 17038 9444 17094 9480
rect 17038 9424 17040 9444
rect 17040 9424 17092 9444
rect 17092 9424 17094 9444
rect 16394 6024 16450 6080
rect 15842 2352 15898 2408
rect 17038 9152 17094 9208
rect 16946 8472 17002 8528
rect 16946 7828 16948 7848
rect 16948 7828 17000 7848
rect 17000 7828 17002 7848
rect 16946 7792 17002 7828
rect 16762 5888 16818 5944
rect 16578 3340 16580 3360
rect 16580 3340 16632 3360
rect 16632 3340 16634 3360
rect 16578 3304 16634 3340
rect 16854 5072 16910 5128
rect 17130 6840 17186 6896
rect 17038 3168 17094 3224
rect 18510 17720 18566 17776
rect 18878 18808 18934 18864
rect 18878 18420 18934 18456
rect 18878 18400 18880 18420
rect 18880 18400 18932 18420
rect 18932 18400 18934 18420
rect 18602 17332 18658 17368
rect 18602 17312 18604 17332
rect 18604 17312 18656 17332
rect 18656 17312 18658 17332
rect 18602 16904 18658 16960
rect 18418 16768 18474 16824
rect 18234 16360 18290 16416
rect 18234 16224 18290 16280
rect 17866 14184 17922 14240
rect 18050 14184 18106 14240
rect 18142 13368 18198 13424
rect 17866 12552 17922 12608
rect 17866 11348 17922 11384
rect 17866 11328 17868 11348
rect 17868 11328 17920 11348
rect 17920 11328 17922 11348
rect 18050 12416 18106 12472
rect 17590 9444 17646 9480
rect 17590 9424 17592 9444
rect 17592 9424 17644 9444
rect 17644 9424 17646 9444
rect 17406 8608 17462 8664
rect 17406 8084 17462 8120
rect 17406 8064 17408 8084
rect 17408 8064 17460 8084
rect 17460 8064 17462 8084
rect 17314 7248 17370 7304
rect 17222 6704 17278 6760
rect 17314 4392 17370 4448
rect 17314 4120 17370 4176
rect 17590 5752 17646 5808
rect 17590 5652 17592 5672
rect 17592 5652 17644 5672
rect 17644 5652 17646 5672
rect 17590 5616 17646 5652
rect 18142 10260 18198 10296
rect 18142 10240 18144 10260
rect 18144 10240 18196 10260
rect 18196 10240 18198 10260
rect 17866 9288 17922 9344
rect 18050 9152 18106 9208
rect 17682 4256 17738 4312
rect 17774 2624 17830 2680
rect 17314 1536 17370 1592
rect 18786 17312 18842 17368
rect 18694 16496 18750 16552
rect 18602 15156 18658 15192
rect 18602 15136 18604 15156
rect 18604 15136 18656 15156
rect 18656 15136 18658 15156
rect 18602 14864 18658 14920
rect 18694 14592 18750 14648
rect 18418 12552 18474 12608
rect 18326 12416 18382 12472
rect 18326 11872 18382 11928
rect 18602 13232 18658 13288
rect 18602 12008 18658 12064
rect 18602 11892 18658 11928
rect 18602 11872 18604 11892
rect 18604 11872 18656 11892
rect 18656 11872 18658 11892
rect 18418 11192 18474 11248
rect 18326 8880 18382 8936
rect 18970 17584 19026 17640
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19798 21256 19854 21312
rect 20350 28872 20406 28928
rect 20258 24792 20314 24848
rect 19154 18944 19210 19000
rect 18878 16224 18934 16280
rect 18878 15952 18934 16008
rect 19154 16768 19210 16824
rect 19062 16632 19118 16688
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19522 20440 19578 20496
rect 19430 20032 19486 20088
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19522 19236 19578 19272
rect 19522 19216 19524 19236
rect 19524 19216 19576 19236
rect 19576 19216 19578 19236
rect 19706 19080 19762 19136
rect 19798 18692 19854 18728
rect 19798 18672 19800 18692
rect 19800 18672 19852 18692
rect 19852 18672 19854 18692
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19706 17720 19762 17776
rect 19614 17584 19670 17640
rect 19982 17720 20038 17776
rect 19062 15816 19118 15872
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19982 17448 20038 17504
rect 19706 17176 19762 17232
rect 19798 16632 19854 16688
rect 20810 27376 20866 27432
rect 20718 25880 20774 25936
rect 20718 25200 20774 25256
rect 20442 20712 20498 20768
rect 21086 37440 21142 37496
rect 20718 20032 20774 20088
rect 20626 19624 20682 19680
rect 20534 19216 20590 19272
rect 20442 18808 20498 18864
rect 20350 18264 20406 18320
rect 20258 17176 20314 17232
rect 20442 17992 20498 18048
rect 20442 17876 20498 17912
rect 20442 17856 20444 17876
rect 20444 17856 20496 17876
rect 20496 17856 20498 17876
rect 20074 16360 20130 16416
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19982 16224 20038 16280
rect 19614 15816 19670 15872
rect 19246 15580 19248 15600
rect 19248 15580 19300 15600
rect 19300 15580 19302 15600
rect 19246 15544 19302 15580
rect 19982 15816 20038 15872
rect 20074 15544 20130 15600
rect 20258 15408 20314 15464
rect 19430 15272 19486 15328
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20166 15308 20168 15328
rect 20168 15308 20220 15328
rect 20220 15308 20222 15328
rect 20166 15272 20222 15308
rect 19982 15136 20038 15192
rect 20718 19080 20774 19136
rect 20534 16360 20590 16416
rect 20534 15952 20590 16008
rect 20534 15544 20590 15600
rect 21178 23432 21234 23488
rect 21362 22344 21418 22400
rect 20902 17876 20958 17912
rect 20902 17856 20904 17876
rect 20904 17856 20956 17876
rect 20956 17856 20958 17876
rect 21270 19488 21326 19544
rect 21638 21120 21694 21176
rect 20810 17312 20866 17368
rect 20810 15680 20866 15736
rect 20718 15564 20774 15600
rect 20718 15544 20720 15564
rect 20720 15544 20772 15564
rect 20772 15544 20774 15564
rect 19154 14592 19210 14648
rect 19522 14728 19578 14784
rect 19154 14048 19210 14104
rect 18878 13096 18934 13152
rect 19246 13504 19302 13560
rect 19430 14184 19486 14240
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 20074 14184 20130 14240
rect 19706 13796 19762 13832
rect 19706 13776 19708 13796
rect 19708 13776 19760 13796
rect 19760 13776 19762 13796
rect 19522 13640 19578 13696
rect 20350 15000 20406 15056
rect 20534 14728 20590 14784
rect 19982 13776 20038 13832
rect 20166 13796 20222 13832
rect 20166 13776 20168 13796
rect 20168 13776 20220 13796
rect 20220 13776 20222 13796
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19706 12860 19708 12880
rect 19708 12860 19760 12880
rect 19760 12860 19762 12880
rect 19706 12824 19762 12860
rect 19614 12588 19616 12608
rect 19616 12588 19668 12608
rect 19668 12588 19670 12608
rect 19614 12552 19670 12588
rect 19062 10920 19118 10976
rect 18786 9968 18842 10024
rect 18510 9696 18566 9752
rect 18602 9424 18658 9480
rect 18694 8492 18750 8528
rect 18694 8472 18696 8492
rect 18696 8472 18748 8492
rect 18748 8472 18750 8492
rect 18602 8084 18658 8120
rect 18602 8064 18604 8084
rect 18604 8064 18656 8084
rect 18656 8064 18658 8084
rect 18326 5344 18382 5400
rect 17866 1672 17922 1728
rect 18234 2624 18290 2680
rect 19706 12300 19762 12336
rect 19706 12280 19708 12300
rect 19708 12280 19760 12300
rect 19760 12280 19762 12300
rect 19430 12008 19486 12064
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19430 11736 19486 11792
rect 19614 11736 19670 11792
rect 19246 10784 19302 10840
rect 19890 11328 19946 11384
rect 20258 11600 20314 11656
rect 20074 11348 20130 11384
rect 20074 11328 20076 11348
rect 20076 11328 20128 11348
rect 20128 11328 20130 11348
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19982 10804 20038 10840
rect 19982 10784 19984 10804
rect 19984 10784 20036 10804
rect 20036 10784 20038 10804
rect 19890 10648 19946 10704
rect 20258 11076 20314 11112
rect 20258 11056 20260 11076
rect 20260 11056 20312 11076
rect 20312 11056 20314 11076
rect 19154 9152 19210 9208
rect 19062 9016 19118 9072
rect 18970 8744 19026 8800
rect 19154 8628 19210 8664
rect 19154 8608 19156 8628
rect 19156 8608 19208 8628
rect 19208 8608 19210 8628
rect 18970 8064 19026 8120
rect 18970 7656 19026 7712
rect 18694 3576 18750 3632
rect 18510 1944 18566 2000
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19430 9696 19486 9752
rect 20074 10104 20130 10160
rect 19522 9424 19578 9480
rect 19890 9016 19946 9072
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 20994 15272 21050 15328
rect 20810 15156 20866 15192
rect 20810 15136 20812 15156
rect 20812 15136 20864 15156
rect 20864 15136 20866 15156
rect 21454 18420 21510 18456
rect 21454 18400 21456 18420
rect 21456 18400 21508 18420
rect 21508 18400 21510 18420
rect 21270 15428 21326 15464
rect 21270 15408 21272 15428
rect 21272 15408 21324 15428
rect 21324 15408 21326 15428
rect 20994 14864 21050 14920
rect 20810 14592 20866 14648
rect 20810 14048 20866 14104
rect 20810 13640 20866 13696
rect 20626 12416 20682 12472
rect 20626 12144 20682 12200
rect 20810 12008 20866 12064
rect 20810 11620 20866 11656
rect 20810 11600 20812 11620
rect 20812 11600 20864 11620
rect 20864 11600 20866 11620
rect 21086 14048 21142 14104
rect 22098 26424 22154 26480
rect 22190 23024 22246 23080
rect 22006 22208 22062 22264
rect 22006 19488 22062 19544
rect 21822 18672 21878 18728
rect 21730 17856 21786 17912
rect 21638 15680 21694 15736
rect 21546 15544 21602 15600
rect 21270 14340 21326 14376
rect 21270 14320 21272 14340
rect 21272 14320 21324 14340
rect 21324 14320 21326 14340
rect 21454 13912 21510 13968
rect 20994 12144 21050 12200
rect 21178 12552 21234 12608
rect 21178 12008 21234 12064
rect 20534 10920 20590 10976
rect 20534 10140 20536 10160
rect 20536 10140 20588 10160
rect 20588 10140 20590 10160
rect 20534 10104 20590 10140
rect 19982 8608 20038 8664
rect 19522 8200 19578 8256
rect 19798 7828 19800 7848
rect 19800 7828 19852 7848
rect 19852 7828 19854 7848
rect 19798 7792 19854 7828
rect 19982 7656 20038 7712
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19430 7404 19486 7440
rect 19430 7384 19432 7404
rect 19432 7384 19484 7404
rect 19484 7384 19486 7404
rect 19338 3460 19394 3496
rect 19706 6704 19762 6760
rect 20074 6568 20130 6624
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19982 6432 20038 6488
rect 19706 5616 19762 5672
rect 20074 6296 20130 6352
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 20534 9832 20590 9888
rect 20994 11056 21050 11112
rect 20810 10920 20866 10976
rect 20902 10376 20958 10432
rect 20902 9832 20958 9888
rect 20626 8336 20682 8392
rect 20350 6296 20406 6352
rect 19338 3440 19340 3460
rect 19340 3440 19392 3460
rect 19392 3440 19394 3460
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20442 3984 20498 4040
rect 20626 6840 20682 6896
rect 20718 4392 20774 4448
rect 21178 10240 21234 10296
rect 21178 9832 21234 9888
rect 21086 7928 21142 7984
rect 21454 13252 21510 13288
rect 21454 13232 21456 13252
rect 21456 13232 21508 13252
rect 21508 13232 21510 13252
rect 21454 12008 21510 12064
rect 21454 11056 21510 11112
rect 21822 16632 21878 16688
rect 22190 20748 22192 20768
rect 22192 20748 22244 20768
rect 22244 20748 22246 20768
rect 22190 20712 22246 20748
rect 22650 20596 22706 20632
rect 22650 20576 22652 20596
rect 22652 20576 22704 20596
rect 22704 20576 22706 20596
rect 23294 29416 23350 29472
rect 23202 26016 23258 26072
rect 22098 16768 22154 16824
rect 22006 16632 22062 16688
rect 22006 15136 22062 15192
rect 21822 14728 21878 14784
rect 21822 13504 21878 13560
rect 21730 13368 21786 13424
rect 21914 13096 21970 13152
rect 21822 12960 21878 13016
rect 21730 12688 21786 12744
rect 22466 17584 22522 17640
rect 22466 17040 22522 17096
rect 22466 16768 22522 16824
rect 22466 16496 22522 16552
rect 22098 13524 22154 13560
rect 22098 13504 22100 13524
rect 22100 13504 22152 13524
rect 22152 13504 22154 13524
rect 21822 12144 21878 12200
rect 21362 8880 21418 8936
rect 21454 8744 21510 8800
rect 21454 8200 21510 8256
rect 21270 7384 21326 7440
rect 21086 5208 21142 5264
rect 20166 992 20222 1048
rect 20718 1536 20774 1592
rect 21546 4120 21602 4176
rect 21914 10412 21916 10432
rect 21916 10412 21968 10432
rect 21968 10412 21970 10432
rect 21914 10376 21970 10412
rect 22098 9172 22154 9208
rect 22098 9152 22100 9172
rect 22100 9152 22152 9172
rect 22152 9152 22154 9172
rect 22190 9016 22246 9072
rect 21914 7928 21970 7984
rect 22926 18420 22982 18456
rect 22926 18400 22928 18420
rect 22928 18400 22980 18420
rect 22980 18400 22982 18420
rect 23478 21428 23480 21448
rect 23480 21428 23532 21448
rect 23532 21428 23534 21448
rect 23478 21392 23534 21428
rect 23202 18264 23258 18320
rect 23662 20032 23718 20088
rect 23478 19624 23534 19680
rect 23386 18264 23442 18320
rect 22926 17040 22982 17096
rect 23294 17720 23350 17776
rect 23110 17176 23166 17232
rect 22834 15272 22890 15328
rect 22742 14728 22798 14784
rect 22742 14048 22798 14104
rect 22650 13504 22706 13560
rect 22558 13368 22614 13424
rect 22742 13368 22798 13424
rect 23294 16768 23350 16824
rect 23294 15000 23350 15056
rect 23202 14320 23258 14376
rect 22558 11056 22614 11112
rect 22558 9152 22614 9208
rect 22558 9036 22614 9072
rect 22558 9016 22560 9036
rect 22560 9016 22612 9036
rect 22612 9016 22614 9036
rect 22374 8064 22430 8120
rect 21914 6840 21970 6896
rect 22282 6840 22338 6896
rect 22190 5636 22246 5672
rect 22190 5616 22192 5636
rect 22192 5616 22244 5636
rect 22244 5616 22246 5636
rect 21914 2760 21970 2816
rect 22374 5208 22430 5264
rect 22098 4528 22154 4584
rect 22190 1284 22246 1320
rect 22190 1264 22192 1284
rect 22192 1264 22244 1284
rect 22244 1264 22246 1284
rect 22742 4392 22798 4448
rect 23478 15952 23534 16008
rect 23386 14068 23442 14104
rect 23386 14048 23388 14068
rect 23388 14048 23440 14068
rect 23440 14048 23442 14068
rect 23570 14184 23626 14240
rect 23846 19352 23902 19408
rect 23662 13912 23718 13968
rect 23662 13368 23718 13424
rect 23570 13232 23626 13288
rect 24214 20168 24270 20224
rect 24030 16940 24032 16960
rect 24032 16940 24084 16960
rect 24084 16940 24086 16960
rect 24030 16904 24086 16940
rect 24030 16088 24086 16144
rect 24030 14884 24086 14920
rect 24030 14864 24032 14884
rect 24032 14864 24084 14884
rect 24084 14864 24086 14884
rect 23846 13368 23902 13424
rect 23570 12960 23626 13016
rect 23754 12960 23810 13016
rect 23478 12708 23534 12744
rect 23478 12688 23480 12708
rect 23480 12688 23532 12708
rect 23532 12688 23534 12708
rect 23110 7248 23166 7304
rect 22926 6704 22982 6760
rect 23570 11500 23572 11520
rect 23572 11500 23624 11520
rect 23624 11500 23626 11520
rect 23570 11464 23626 11500
rect 23846 8608 23902 8664
rect 22926 5752 22982 5808
rect 22926 5092 22982 5128
rect 22926 5072 22928 5092
rect 22928 5072 22980 5092
rect 22980 5072 22982 5092
rect 23110 4120 23166 4176
rect 23846 7520 23902 7576
rect 24674 30368 24730 30424
rect 24582 25336 24638 25392
rect 24398 23704 24454 23760
rect 24306 17856 24362 17912
rect 24490 20476 24492 20496
rect 24492 20476 24544 20496
rect 24544 20476 24546 20496
rect 24490 20440 24546 20476
rect 24398 15680 24454 15736
rect 24766 19080 24822 19136
rect 25042 28872 25098 28928
rect 25042 19488 25098 19544
rect 24950 18964 25006 19000
rect 24950 18944 24952 18964
rect 24952 18944 25004 18964
rect 25004 18944 25006 18964
rect 24950 18808 25006 18864
rect 24858 18672 24914 18728
rect 24766 17448 24822 17504
rect 24582 16360 24638 16416
rect 25502 23160 25558 23216
rect 25502 19252 25504 19272
rect 25504 19252 25556 19272
rect 25556 19252 25558 19272
rect 25502 19216 25558 19252
rect 25502 18264 25558 18320
rect 24490 15544 24546 15600
rect 24214 15136 24270 15192
rect 24398 11464 24454 11520
rect 24398 11348 24454 11384
rect 24398 11328 24400 11348
rect 24400 11328 24452 11348
rect 24452 11328 24454 11348
rect 23846 6704 23902 6760
rect 23570 6332 23572 6352
rect 23572 6332 23624 6352
rect 23624 6332 23626 6352
rect 23570 6296 23626 6332
rect 23662 4936 23718 4992
rect 23570 4684 23626 4720
rect 23570 4664 23572 4684
rect 23572 4664 23624 4684
rect 23624 4664 23626 4684
rect 24214 9596 24216 9616
rect 24216 9596 24268 9616
rect 24268 9596 24270 9616
rect 24214 9560 24270 9596
rect 24030 4120 24086 4176
rect 24490 8880 24546 8936
rect 24674 14456 24730 14512
rect 24674 10548 24676 10568
rect 24676 10548 24728 10568
rect 24728 10548 24730 10568
rect 24674 10512 24730 10548
rect 24950 10376 25006 10432
rect 24858 9424 24914 9480
rect 25042 9288 25098 9344
rect 24858 8744 24914 8800
rect 25042 8780 25044 8800
rect 25044 8780 25096 8800
rect 25096 8780 25098 8800
rect 25042 8744 25098 8780
rect 25042 8200 25098 8256
rect 25318 16244 25374 16280
rect 25318 16224 25320 16244
rect 25320 16224 25372 16244
rect 25372 16224 25374 16244
rect 25318 15408 25374 15464
rect 25226 15136 25282 15192
rect 25318 13232 25374 13288
rect 25226 11872 25282 11928
rect 25226 10648 25282 10704
rect 25226 10376 25282 10432
rect 25226 9288 25282 9344
rect 25502 15136 25558 15192
rect 25686 12436 25742 12472
rect 25686 12416 25688 12436
rect 25688 12416 25740 12436
rect 25740 12416 25742 12436
rect 25686 10920 25742 10976
rect 25870 19352 25926 19408
rect 26054 19352 26110 19408
rect 26146 15816 26202 15872
rect 26054 15272 26110 15328
rect 26054 13232 26110 13288
rect 25962 13096 26018 13152
rect 25870 12824 25926 12880
rect 26790 24656 26846 24712
rect 26330 16224 26386 16280
rect 26330 15952 26386 16008
rect 26330 15700 26386 15736
rect 26330 15680 26332 15700
rect 26332 15680 26384 15700
rect 26384 15680 26386 15700
rect 26238 12280 26294 12336
rect 26238 11192 26294 11248
rect 25686 10104 25742 10160
rect 25502 9832 25558 9888
rect 25594 8084 25650 8120
rect 25594 8064 25596 8084
rect 25596 8064 25648 8084
rect 25648 8064 25650 8084
rect 24582 3440 24638 3496
rect 24398 1128 24454 1184
rect 24950 4120 25006 4176
rect 25134 3884 25136 3904
rect 25136 3884 25188 3904
rect 25188 3884 25190 3904
rect 25134 3848 25190 3884
rect 26238 9968 26294 10024
rect 25962 9596 25964 9616
rect 25964 9596 26016 9616
rect 26016 9596 26018 9616
rect 25962 9560 26018 9596
rect 26606 18572 26608 18592
rect 26608 18572 26660 18592
rect 26660 18572 26662 18592
rect 26606 18536 26662 18572
rect 25962 8372 25964 8392
rect 25964 8372 26016 8392
rect 26016 8372 26018 8392
rect 25962 8336 26018 8372
rect 26146 7112 26202 7168
rect 25962 2508 26018 2544
rect 25962 2488 25964 2508
rect 25964 2488 26016 2508
rect 26016 2488 26018 2508
rect 26422 1808 26478 1864
rect 27618 35264 27674 35320
rect 27526 25608 27582 25664
rect 26974 19352 27030 19408
rect 27066 16768 27122 16824
rect 26974 14728 27030 14784
rect 27250 19216 27306 19272
rect 27158 10104 27214 10160
rect 27894 25880 27950 25936
rect 27618 19780 27674 19816
rect 27618 19760 27620 19780
rect 27620 19760 27672 19780
rect 27672 19760 27674 19780
rect 27526 17176 27582 17232
rect 27434 14612 27490 14648
rect 27434 14592 27436 14612
rect 27436 14592 27488 14612
rect 27488 14592 27490 14612
rect 27710 15020 27766 15056
rect 27710 15000 27712 15020
rect 27712 15000 27764 15020
rect 27764 15000 27766 15020
rect 28262 25744 28318 25800
rect 27986 17176 28042 17232
rect 27526 14320 27582 14376
rect 27434 14184 27490 14240
rect 27434 12044 27436 12064
rect 27436 12044 27488 12064
rect 27488 12044 27490 12064
rect 27434 12008 27490 12044
rect 27894 13232 27950 13288
rect 27710 10784 27766 10840
rect 27986 11756 28042 11792
rect 27986 11736 27988 11756
rect 27988 11736 28040 11756
rect 28040 11736 28042 11756
rect 26882 6840 26938 6896
rect 26882 6432 26938 6488
rect 27158 5908 27214 5944
rect 27158 5888 27160 5908
rect 27160 5888 27212 5908
rect 27212 5888 27214 5908
rect 27342 5072 27398 5128
rect 27802 5908 27858 5944
rect 27802 5888 27804 5908
rect 27804 5888 27856 5908
rect 27856 5888 27858 5908
rect 28170 18128 28226 18184
rect 28354 20596 28410 20632
rect 28354 20576 28356 20596
rect 28356 20576 28408 20596
rect 28408 20576 28410 20596
rect 28446 19080 28502 19136
rect 28262 17876 28318 17912
rect 28262 17856 28264 17876
rect 28264 17856 28316 17876
rect 28316 17856 28318 17876
rect 28262 13640 28318 13696
rect 28998 28464 29054 28520
rect 29090 20168 29146 20224
rect 29090 19488 29146 19544
rect 28998 17040 29054 17096
rect 28630 14456 28686 14512
rect 28262 12824 28318 12880
rect 28170 12416 28226 12472
rect 27986 1944 28042 2000
rect 28538 5480 28594 5536
rect 28998 10104 29054 10160
rect 30286 29280 30342 29336
rect 29458 16768 29514 16824
rect 29274 14068 29330 14104
rect 29274 14048 29276 14068
rect 29276 14048 29328 14068
rect 29328 14048 29330 14068
rect 29274 13776 29330 13832
rect 29090 6704 29146 6760
rect 28906 4800 28962 4856
rect 29550 16668 29552 16688
rect 29552 16668 29604 16688
rect 29604 16668 29606 16688
rect 29550 16632 29606 16668
rect 30654 29416 30710 29472
rect 29734 12960 29790 13016
rect 30194 19488 30250 19544
rect 30286 19216 30342 19272
rect 29550 12300 29606 12336
rect 29550 12280 29552 12300
rect 29552 12280 29604 12300
rect 29604 12280 29606 12300
rect 29458 3712 29514 3768
rect 29918 11464 29974 11520
rect 30378 13504 30434 13560
rect 30562 22380 30564 22400
rect 30564 22380 30616 22400
rect 30616 22380 30618 22400
rect 30562 22344 30618 22380
rect 30470 13368 30526 13424
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 31114 30368 31170 30424
rect 31850 26696 31906 26752
rect 31298 22380 31300 22400
rect 31300 22380 31352 22400
rect 31352 22380 31354 22400
rect 31298 22344 31354 22380
rect 31114 14728 31170 14784
rect 30930 11600 30986 11656
rect 31390 19660 31392 19680
rect 31392 19660 31444 19680
rect 31444 19660 31446 19680
rect 31390 19624 31446 19660
rect 31666 21392 31722 21448
rect 31666 19216 31722 19272
rect 31666 18264 31722 18320
rect 31574 16224 31630 16280
rect 31666 12416 31722 12472
rect 31666 12280 31722 12336
rect 31666 9288 31722 9344
rect 30378 1400 30434 1456
rect 32126 23296 32182 23352
rect 31942 21936 31998 21992
rect 31850 9832 31906 9888
rect 32034 19488 32090 19544
rect 32586 20168 32642 20224
rect 32310 12688 32366 12744
rect 31942 7928 31998 7984
rect 31942 3576 31998 3632
rect 32862 26560 32918 26616
rect 32678 8744 32734 8800
rect 33230 11872 33286 11928
rect 33782 19624 33838 19680
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34702 34584 34758 34640
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34518 30504 34574 30560
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34518 29008 34574 29064
rect 33690 10376 33746 10432
rect 33598 9152 33654 9208
rect 33414 8472 33470 8528
rect 32954 7792 33010 7848
rect 32862 7384 32918 7440
rect 32770 6160 32826 6216
rect 33230 2916 33286 2952
rect 33230 2896 33232 2916
rect 33232 2896 33284 2916
rect 33284 2896 33286 2916
rect 33874 5208 33930 5264
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34794 27648 34850 27704
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35438 20984 35494 21040
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34794 12008 34850 12064
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35530 20440 35586 20496
rect 35438 10512 35494 10568
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34702 9016 34758 9072
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34518 8064 34574 8120
rect 34150 7520 34206 7576
rect 34058 5072 34114 5128
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34518 3068 34520 3088
rect 34520 3068 34572 3088
rect 34572 3068 34574 3088
rect 34518 3032 34574 3068
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35070 2524 35072 2544
rect 35072 2524 35124 2544
rect 35124 2524 35126 2544
rect 35070 2488 35126 2524
rect 37278 32408 37334 32464
rect 40406 37304 40462 37360
rect 41234 37848 41290 37904
rect 40774 21392 40830 21448
rect 44086 29996 44088 30016
rect 44088 29996 44140 30016
rect 44140 29996 44142 30016
rect 44086 29960 44142 29996
rect 35898 14320 35954 14376
rect 37462 6568 37518 6624
rect 38014 9968 38070 10024
rect 42062 14864 42118 14920
rect 42522 11736 42578 11792
rect 42246 11600 42302 11656
rect 39854 4256 39910 4312
rect 39394 4120 39450 4176
rect 40222 3168 40278 3224
rect 43258 10920 43314 10976
rect 43074 8880 43130 8936
rect 42890 2352 42946 2408
rect 43350 10512 43406 10568
rect 44086 9968 44142 10024
rect 40130 584 40186 640
<< metal3 >>
rect 0 39674 800 39704
rect 3969 39674 4035 39677
rect 0 39672 4035 39674
rect 0 39616 3974 39672
rect 4030 39616 4035 39672
rect 0 39614 4035 39616
rect 0 39584 800 39614
rect 3969 39611 4035 39614
rect 0 39130 800 39160
rect 2865 39130 2931 39133
rect 0 39128 2931 39130
rect 0 39072 2870 39128
rect 2926 39072 2931 39128
rect 0 39070 2931 39072
rect 0 39040 800 39070
rect 2865 39067 2931 39070
rect 0 38586 800 38616
rect 3509 38586 3575 38589
rect 0 38584 3575 38586
rect 0 38528 3514 38584
rect 3570 38528 3575 38584
rect 0 38526 3575 38528
rect 0 38496 800 38526
rect 3509 38523 3575 38526
rect 0 37906 800 37936
rect 3141 37906 3207 37909
rect 0 37904 3207 37906
rect 0 37848 3146 37904
rect 3202 37848 3207 37904
rect 0 37846 3207 37848
rect 0 37816 800 37846
rect 3141 37843 3207 37846
rect 27470 37844 27476 37908
rect 27540 37906 27546 37908
rect 41229 37906 41295 37909
rect 27540 37904 41295 37906
rect 27540 37848 41234 37904
rect 41290 37848 41295 37904
rect 27540 37846 41295 37848
rect 27540 37844 27546 37846
rect 41229 37843 41295 37846
rect 5349 37634 5415 37637
rect 22502 37634 22508 37636
rect 5349 37632 22508 37634
rect 5349 37576 5354 37632
rect 5410 37576 22508 37632
rect 5349 37574 22508 37576
rect 5349 37571 5415 37574
rect 22502 37572 22508 37574
rect 22572 37572 22578 37636
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 4705 37498 4771 37501
rect 18086 37498 18092 37500
rect 4705 37496 18092 37498
rect 4705 37440 4710 37496
rect 4766 37440 18092 37496
rect 4705 37438 18092 37440
rect 4705 37435 4771 37438
rect 18086 37436 18092 37438
rect 18156 37436 18162 37500
rect 21081 37498 21147 37501
rect 28390 37498 28396 37500
rect 21081 37496 28396 37498
rect 21081 37440 21086 37496
rect 21142 37440 28396 37496
rect 21081 37438 28396 37440
rect 21081 37435 21147 37438
rect 28390 37436 28396 37438
rect 28460 37436 28466 37500
rect 0 37362 800 37392
rect 3693 37362 3759 37365
rect 0 37360 3759 37362
rect 0 37304 3698 37360
rect 3754 37304 3759 37360
rect 0 37302 3759 37304
rect 0 37272 800 37302
rect 3693 37299 3759 37302
rect 8109 37362 8175 37365
rect 15878 37362 15884 37364
rect 8109 37360 15884 37362
rect 8109 37304 8114 37360
rect 8170 37304 15884 37360
rect 8109 37302 15884 37304
rect 8109 37299 8175 37302
rect 15878 37300 15884 37302
rect 15948 37300 15954 37364
rect 23974 37300 23980 37364
rect 24044 37362 24050 37364
rect 40401 37362 40467 37365
rect 24044 37360 40467 37362
rect 24044 37304 40406 37360
rect 40462 37304 40467 37360
rect 24044 37302 40467 37304
rect 24044 37300 24050 37302
rect 40401 37299 40467 37302
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36848
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36728 800 36758
rect 2773 36755 2839 36758
rect 17033 36548 17099 36549
rect 17769 36548 17835 36549
rect 16982 36546 16988 36548
rect 16942 36486 16988 36546
rect 17052 36544 17099 36548
rect 17718 36546 17724 36548
rect 17094 36488 17099 36544
rect 16982 36484 16988 36486
rect 17052 36484 17099 36488
rect 17678 36486 17724 36546
rect 17788 36544 17835 36548
rect 17830 36488 17835 36544
rect 17718 36484 17724 36486
rect 17788 36484 17835 36488
rect 17033 36483 17099 36484
rect 17769 36483 17835 36484
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36168
rect 4061 36138 4127 36141
rect 0 36136 4127 36138
rect 0 36080 4066 36136
rect 4122 36080 4127 36136
rect 0 36078 4127 36080
rect 0 36048 800 36078
rect 4061 36075 4127 36078
rect 19374 36076 19380 36140
rect 19444 36138 19450 36140
rect 19885 36138 19951 36141
rect 19444 36136 19951 36138
rect 19444 36080 19890 36136
rect 19946 36080 19951 36136
rect 19444 36078 19951 36080
rect 19444 36076 19450 36078
rect 19885 36075 19951 36078
rect 4981 36002 5047 36005
rect 14365 36004 14431 36005
rect 5574 36002 5580 36004
rect 4981 36000 5580 36002
rect 4981 35944 4986 36000
rect 5042 35944 5580 36000
rect 4981 35942 5580 35944
rect 4981 35939 5047 35942
rect 5574 35940 5580 35942
rect 5644 35940 5650 36004
rect 14365 36000 14412 36004
rect 14476 36002 14482 36004
rect 14365 35944 14370 36000
rect 14365 35940 14412 35944
rect 14476 35942 14522 36002
rect 14476 35940 14482 35942
rect 14365 35939 14431 35940
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35594 800 35624
rect 1393 35594 1459 35597
rect 0 35592 1459 35594
rect 0 35536 1398 35592
rect 1454 35536 1459 35592
rect 0 35534 1459 35536
rect 0 35504 800 35534
rect 1393 35531 1459 35534
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 19425 35322 19491 35325
rect 27613 35322 27679 35325
rect 19425 35320 27679 35322
rect 19425 35264 19430 35320
rect 19486 35264 27618 35320
rect 27674 35264 27679 35320
rect 19425 35262 27679 35264
rect 19425 35259 19491 35262
rect 27613 35259 27679 35262
rect 0 35050 800 35080
rect 3509 35050 3575 35053
rect 0 35048 3575 35050
rect 0 34992 3514 35048
rect 3570 34992 3575 35048
rect 0 34990 3575 34992
rect 0 34960 800 34990
rect 3509 34987 3575 34990
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 4705 34644 4771 34645
rect 4654 34642 4660 34644
rect 4614 34582 4660 34642
rect 4724 34640 4771 34644
rect 4766 34584 4771 34640
rect 4654 34580 4660 34582
rect 4724 34580 4771 34584
rect 4705 34579 4771 34580
rect 13721 34642 13787 34645
rect 14958 34642 14964 34644
rect 13721 34640 14964 34642
rect 13721 34584 13726 34640
rect 13782 34584 14964 34640
rect 13721 34582 14964 34584
rect 13721 34579 13787 34582
rect 14958 34580 14964 34582
rect 15028 34580 15034 34644
rect 17534 34580 17540 34644
rect 17604 34642 17610 34644
rect 18321 34642 18387 34645
rect 17604 34640 18387 34642
rect 17604 34584 18326 34640
rect 18382 34584 18387 34640
rect 17604 34582 18387 34584
rect 17604 34580 17610 34582
rect 18321 34579 18387 34582
rect 26734 34580 26740 34644
rect 26804 34642 26810 34644
rect 34697 34642 34763 34645
rect 26804 34640 34763 34642
rect 26804 34584 34702 34640
rect 34758 34584 34763 34640
rect 26804 34582 34763 34584
rect 26804 34580 26810 34582
rect 34697 34579 34763 34582
rect 0 34370 800 34400
rect 1393 34370 1459 34373
rect 0 34368 1459 34370
rect 0 34312 1398 34368
rect 1454 34312 1459 34368
rect 0 34310 1459 34312
rect 0 34280 800 34310
rect 1393 34307 1459 34310
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33826 800 33856
rect 3601 33826 3667 33829
rect 0 33824 3667 33826
rect 0 33768 3606 33824
rect 3662 33768 3667 33824
rect 0 33766 3667 33768
rect 0 33736 800 33766
rect 3601 33763 3667 33766
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33282 800 33312
rect 1485 33282 1551 33285
rect 0 33280 1551 33282
rect 0 33224 1490 33280
rect 1546 33224 1551 33280
rect 0 33222 1551 33224
rect 0 33192 800 33222
rect 1485 33219 1551 33222
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 19568 32672 19888 32673
rect 0 32602 800 32632
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 3417 32602 3483 32605
rect 0 32600 3483 32602
rect 0 32544 3422 32600
rect 3478 32544 3483 32600
rect 0 32542 3483 32544
rect 0 32512 800 32542
rect 3417 32539 3483 32542
rect 10869 32466 10935 32469
rect 22686 32466 22692 32468
rect 10869 32464 22692 32466
rect 10869 32408 10874 32464
rect 10930 32408 22692 32464
rect 10869 32406 22692 32408
rect 10869 32403 10935 32406
rect 22686 32404 22692 32406
rect 22756 32404 22762 32468
rect 25998 32404 26004 32468
rect 26068 32466 26074 32468
rect 37273 32466 37339 32469
rect 26068 32464 37339 32466
rect 26068 32408 37278 32464
rect 37334 32408 37339 32464
rect 26068 32406 37339 32408
rect 26068 32404 26074 32406
rect 37273 32403 37339 32406
rect 4208 32128 4528 32129
rect 0 32058 800 32088
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 1485 32058 1551 32061
rect 0 32056 1551 32058
rect 0 32000 1490 32056
rect 1546 32000 1551 32056
rect 0 31998 1551 32000
rect 0 31968 800 31998
rect 1485 31995 1551 31998
rect 19568 31584 19888 31585
rect 0 31514 800 31544
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 2865 31514 2931 31517
rect 0 31512 2931 31514
rect 0 31456 2870 31512
rect 2926 31456 2931 31512
rect 0 31454 2931 31456
rect 0 31424 800 31454
rect 2865 31451 2931 31454
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30834 800 30864
rect 1393 30834 1459 30837
rect 0 30832 1459 30834
rect 0 30776 1398 30832
rect 1454 30776 1459 30832
rect 0 30774 1459 30776
rect 0 30744 800 30774
rect 1393 30771 1459 30774
rect 13169 30562 13235 30565
rect 17902 30562 17908 30564
rect 13169 30560 17908 30562
rect 13169 30504 13174 30560
rect 13230 30504 17908 30560
rect 13169 30502 17908 30504
rect 13169 30499 13235 30502
rect 17902 30500 17908 30502
rect 17972 30500 17978 30564
rect 27286 30500 27292 30564
rect 27356 30562 27362 30564
rect 34513 30562 34579 30565
rect 27356 30560 34579 30562
rect 27356 30504 34518 30560
rect 34574 30504 34579 30560
rect 27356 30502 34579 30504
rect 27356 30500 27362 30502
rect 34513 30499 34579 30502
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 13353 30426 13419 30429
rect 14774 30426 14780 30428
rect 13353 30424 14780 30426
rect 13353 30368 13358 30424
rect 13414 30368 14780 30424
rect 13353 30366 14780 30368
rect 13353 30363 13419 30366
rect 14774 30364 14780 30366
rect 14844 30364 14850 30428
rect 24669 30426 24735 30429
rect 31109 30426 31175 30429
rect 24669 30424 31175 30426
rect 24669 30368 24674 30424
rect 24730 30368 31114 30424
rect 31170 30368 31175 30424
rect 24669 30366 31175 30368
rect 24669 30363 24735 30366
rect 31109 30363 31175 30366
rect 0 30290 800 30320
rect 3509 30290 3575 30293
rect 0 30288 3575 30290
rect 0 30232 3514 30288
rect 3570 30232 3575 30288
rect 0 30230 3575 30232
rect 0 30200 800 30230
rect 3509 30227 3575 30230
rect 44081 30018 44147 30021
rect 45200 30018 46000 30048
rect 44081 30016 46000 30018
rect 44081 29960 44086 30016
rect 44142 29960 46000 30016
rect 44081 29958 46000 29960
rect 44081 29955 44147 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 45200 29928 46000 29958
rect 34928 29887 35248 29888
rect 0 29746 800 29776
rect 1393 29746 1459 29749
rect 0 29744 1459 29746
rect 0 29688 1398 29744
rect 1454 29688 1459 29744
rect 0 29686 1459 29688
rect 0 29656 800 29686
rect 1393 29683 1459 29686
rect 23289 29474 23355 29477
rect 30649 29474 30715 29477
rect 23289 29472 30715 29474
rect 23289 29416 23294 29472
rect 23350 29416 30654 29472
rect 30710 29416 30715 29472
rect 23289 29414 30715 29416
rect 23289 29411 23355 29414
rect 30649 29411 30715 29414
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 25446 29276 25452 29340
rect 25516 29338 25522 29340
rect 30281 29338 30347 29341
rect 25516 29336 30347 29338
rect 25516 29280 30286 29336
rect 30342 29280 30347 29336
rect 25516 29278 30347 29280
rect 25516 29276 25522 29278
rect 30281 29275 30347 29278
rect 5942 29140 5948 29204
rect 6012 29202 6018 29204
rect 33174 29202 33180 29204
rect 6012 29142 33180 29202
rect 6012 29140 6018 29142
rect 33174 29140 33180 29142
rect 33244 29140 33250 29204
rect 0 29066 800 29096
rect 3877 29068 3943 29069
rect 3550 29066 3556 29068
rect 0 29006 3556 29066
rect 0 28976 800 29006
rect 3550 29004 3556 29006
rect 3620 29004 3626 29068
rect 3877 29066 3924 29068
rect 3832 29064 3924 29066
rect 3832 29008 3882 29064
rect 3832 29006 3924 29008
rect 3877 29004 3924 29006
rect 3988 29004 3994 29068
rect 5206 29004 5212 29068
rect 5276 29066 5282 29068
rect 34513 29066 34579 29069
rect 5276 29064 34579 29066
rect 5276 29008 34518 29064
rect 34574 29008 34579 29064
rect 5276 29006 34579 29008
rect 5276 29004 5282 29006
rect 3877 29003 3943 29004
rect 34513 29003 34579 29006
rect 9489 28930 9555 28933
rect 15142 28930 15148 28932
rect 9489 28928 15148 28930
rect 9489 28872 9494 28928
rect 9550 28872 15148 28928
rect 9489 28870 15148 28872
rect 9489 28867 9555 28870
rect 15142 28868 15148 28870
rect 15212 28868 15218 28932
rect 20345 28930 20411 28933
rect 25037 28930 25103 28933
rect 20345 28928 25103 28930
rect 20345 28872 20350 28928
rect 20406 28872 25042 28928
rect 25098 28872 25103 28928
rect 20345 28870 25103 28872
rect 20345 28867 20411 28870
rect 25037 28867 25103 28870
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28522 800 28552
rect 1485 28522 1551 28525
rect 0 28520 1551 28522
rect 0 28464 1490 28520
rect 1546 28464 1551 28520
rect 0 28462 1551 28464
rect 0 28432 800 28462
rect 1485 28459 1551 28462
rect 18454 28460 18460 28524
rect 18524 28522 18530 28524
rect 28993 28522 29059 28525
rect 18524 28520 29059 28522
rect 18524 28464 28998 28520
rect 29054 28464 29059 28520
rect 18524 28462 29059 28464
rect 18524 28460 18530 28462
rect 28993 28459 29059 28462
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 1342 28052 1348 28116
rect 1412 28114 1418 28116
rect 23422 28114 23428 28116
rect 1412 28054 23428 28114
rect 1412 28052 1418 28054
rect 23422 28052 23428 28054
rect 23492 28052 23498 28116
rect 0 27978 800 28008
rect 3417 27978 3483 27981
rect 0 27976 3483 27978
rect 0 27920 3422 27976
rect 3478 27920 3483 27976
rect 0 27918 3483 27920
rect 0 27888 800 27918
rect 3417 27915 3483 27918
rect 6862 27916 6868 27980
rect 6932 27978 6938 27980
rect 20478 27978 20484 27980
rect 6932 27918 20484 27978
rect 6932 27916 6938 27918
rect 20478 27916 20484 27918
rect 20548 27916 20554 27980
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 10409 27706 10475 27709
rect 34789 27706 34855 27709
rect 10409 27704 34855 27706
rect 10409 27648 10414 27704
rect 10470 27648 34794 27704
rect 34850 27648 34855 27704
rect 10409 27646 34855 27648
rect 10409 27643 10475 27646
rect 34789 27643 34855 27646
rect 933 27434 999 27437
rect 20805 27434 20871 27437
rect 933 27432 20871 27434
rect 933 27376 938 27432
rect 994 27376 20810 27432
rect 20866 27376 20871 27432
rect 933 27374 20871 27376
rect 933 27371 999 27374
rect 20805 27371 20871 27374
rect 0 27298 800 27328
rect 1393 27298 1459 27301
rect 0 27296 1459 27298
rect 0 27240 1398 27296
rect 1454 27240 1459 27296
rect 0 27238 1459 27240
rect 0 27208 800 27238
rect 1393 27235 1459 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 7373 27162 7439 27165
rect 7598 27162 7604 27164
rect 7373 27160 7604 27162
rect 7373 27104 7378 27160
rect 7434 27104 7604 27160
rect 7373 27102 7604 27104
rect 7373 27099 7439 27102
rect 7598 27100 7604 27102
rect 7668 27100 7674 27164
rect 12709 27026 12775 27029
rect 16062 27026 16068 27028
rect 12709 27024 16068 27026
rect 12709 26968 12714 27024
rect 12770 26968 16068 27024
rect 12709 26966 16068 26968
rect 12709 26963 12775 26966
rect 16062 26964 16068 26966
rect 16132 26964 16138 27028
rect 6913 26890 6979 26893
rect 7046 26890 7052 26892
rect 6913 26888 7052 26890
rect 6913 26832 6918 26888
rect 6974 26832 7052 26888
rect 6913 26830 7052 26832
rect 6913 26827 6979 26830
rect 7046 26828 7052 26830
rect 7116 26828 7122 26892
rect 24894 26890 24900 26892
rect 9446 26830 24900 26890
rect 0 26754 800 26784
rect 4061 26754 4127 26757
rect 0 26752 4127 26754
rect 0 26696 4066 26752
rect 4122 26696 4127 26752
rect 0 26694 4127 26696
rect 0 26664 800 26694
rect 4061 26691 4127 26694
rect 7230 26692 7236 26756
rect 7300 26754 7306 26756
rect 8569 26754 8635 26757
rect 9446 26754 9506 26830
rect 24894 26828 24900 26830
rect 24964 26828 24970 26892
rect 7300 26752 9506 26754
rect 7300 26696 8574 26752
rect 8630 26696 9506 26752
rect 7300 26694 9506 26696
rect 7300 26692 7306 26694
rect 8569 26691 8635 26694
rect 11830 26692 11836 26756
rect 11900 26754 11906 26756
rect 31845 26754 31911 26757
rect 11900 26752 31911 26754
rect 11900 26696 31850 26752
rect 31906 26696 31911 26752
rect 11900 26694 31911 26696
rect 11900 26692 11906 26694
rect 31845 26691 31911 26694
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 13302 26556 13308 26620
rect 13372 26618 13378 26620
rect 32857 26618 32923 26621
rect 13372 26616 32923 26618
rect 13372 26560 32862 26616
rect 32918 26560 32923 26616
rect 13372 26558 32923 26560
rect 13372 26556 13378 26558
rect 32857 26555 32923 26558
rect 9489 26484 9555 26485
rect 9438 26482 9444 26484
rect 9398 26422 9444 26482
rect 9508 26480 9555 26484
rect 9550 26424 9555 26480
rect 9438 26420 9444 26422
rect 9508 26420 9555 26424
rect 9489 26419 9555 26420
rect 12617 26482 12683 26485
rect 12750 26482 12756 26484
rect 12617 26480 12756 26482
rect 12617 26424 12622 26480
rect 12678 26424 12756 26480
rect 12617 26422 12756 26424
rect 12617 26419 12683 26422
rect 12750 26420 12756 26422
rect 12820 26420 12826 26484
rect 14038 26420 14044 26484
rect 14108 26482 14114 26484
rect 22093 26482 22159 26485
rect 14108 26480 22159 26482
rect 14108 26424 22098 26480
rect 22154 26424 22159 26480
rect 14108 26422 22159 26424
rect 14108 26420 14114 26422
rect 22093 26419 22159 26422
rect 1158 26284 1164 26348
rect 1228 26346 1234 26348
rect 13077 26346 13143 26349
rect 1228 26344 13143 26346
rect 1228 26288 13082 26344
rect 13138 26288 13143 26344
rect 1228 26286 13143 26288
rect 1228 26284 1234 26286
rect 13077 26283 13143 26286
rect 13721 26346 13787 26349
rect 21030 26346 21036 26348
rect 13721 26344 21036 26346
rect 13721 26288 13726 26344
rect 13782 26288 21036 26344
rect 13721 26286 21036 26288
rect 13721 26283 13787 26286
rect 21030 26284 21036 26286
rect 21100 26284 21106 26348
rect 0 26210 800 26240
rect 1393 26210 1459 26213
rect 6913 26212 6979 26213
rect 0 26208 1459 26210
rect 0 26152 1398 26208
rect 1454 26152 1459 26208
rect 0 26150 1459 26152
rect 0 26120 800 26150
rect 1393 26147 1459 26150
rect 6862 26148 6868 26212
rect 6932 26210 6979 26212
rect 6932 26208 7024 26210
rect 6974 26152 7024 26208
rect 6932 26150 7024 26152
rect 6932 26148 6979 26150
rect 6913 26147 6979 26148
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 18505 26074 18571 26077
rect 23197 26074 23263 26077
rect 2730 26072 18571 26074
rect 2730 26016 18510 26072
rect 18566 26016 18571 26072
rect 2730 26014 18571 26016
rect 0 25530 800 25560
rect 2730 25530 2790 26014
rect 18505 26011 18571 26014
rect 20532 26072 23263 26074
rect 20532 26016 23202 26072
rect 23258 26016 23263 26072
rect 20532 26014 23263 26016
rect 12709 25938 12775 25941
rect 20532 25938 20592 26014
rect 23197 26011 23263 26014
rect 12709 25936 20592 25938
rect 12709 25880 12714 25936
rect 12770 25880 20592 25936
rect 12709 25878 20592 25880
rect 20713 25938 20779 25941
rect 27889 25938 27955 25941
rect 20713 25936 27955 25938
rect 20713 25880 20718 25936
rect 20774 25880 27894 25936
rect 27950 25880 27955 25936
rect 20713 25878 27955 25880
rect 12709 25875 12775 25878
rect 20713 25875 20779 25878
rect 27889 25875 27955 25878
rect 28257 25802 28323 25805
rect 12390 25800 28323 25802
rect 12390 25744 28262 25800
rect 28318 25744 28323 25800
rect 12390 25742 28323 25744
rect 11094 25604 11100 25668
rect 11164 25666 11170 25668
rect 11513 25666 11579 25669
rect 12390 25666 12450 25742
rect 28257 25739 28323 25742
rect 11164 25664 12450 25666
rect 11164 25608 11518 25664
rect 11574 25608 12450 25664
rect 11164 25606 12450 25608
rect 12525 25666 12591 25669
rect 27521 25666 27587 25669
rect 12525 25664 27587 25666
rect 12525 25608 12530 25664
rect 12586 25608 27526 25664
rect 27582 25608 27587 25664
rect 12525 25606 27587 25608
rect 11164 25604 11170 25606
rect 11513 25603 11579 25606
rect 12525 25603 12591 25606
rect 27521 25603 27587 25606
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25470 2790 25530
rect 0 25440 800 25470
rect 9070 25468 9076 25532
rect 9140 25530 9146 25532
rect 29310 25530 29316 25532
rect 9140 25470 29316 25530
rect 9140 25468 9146 25470
rect 29310 25468 29316 25470
rect 29380 25468 29386 25532
rect 15193 25394 15259 25397
rect 24577 25394 24643 25397
rect 15193 25392 24643 25394
rect 15193 25336 15198 25392
rect 15254 25336 24582 25392
rect 24638 25336 24643 25392
rect 15193 25334 24643 25336
rect 15193 25331 15259 25334
rect 24577 25331 24643 25334
rect 12525 25258 12591 25261
rect 13077 25258 13143 25261
rect 20713 25258 20779 25261
rect 12525 25256 20779 25258
rect 12525 25200 12530 25256
rect 12586 25200 13082 25256
rect 13138 25200 20718 25256
rect 20774 25200 20779 25256
rect 12525 25198 20779 25200
rect 12525 25195 12591 25198
rect 13077 25195 13143 25198
rect 20713 25195 20779 25198
rect 10358 25060 10364 25124
rect 10428 25122 10434 25124
rect 11421 25122 11487 25125
rect 10428 25120 11487 25122
rect 10428 25064 11426 25120
rect 11482 25064 11487 25120
rect 10428 25062 11487 25064
rect 10428 25060 10434 25062
rect 11421 25059 11487 25062
rect 19568 25056 19888 25057
rect 0 24986 800 25016
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 1393 24986 1459 24989
rect 0 24984 1459 24986
rect 0 24928 1398 24984
rect 1454 24928 1459 24984
rect 0 24926 1459 24928
rect 0 24896 800 24926
rect 1393 24923 1459 24926
rect 11513 24986 11579 24989
rect 14917 24986 14983 24989
rect 11513 24984 14983 24986
rect 11513 24928 11518 24984
rect 11574 24928 14922 24984
rect 14978 24928 14983 24984
rect 11513 24926 14983 24928
rect 11513 24923 11579 24926
rect 14917 24923 14983 24926
rect 20118 24926 20914 24986
rect 8661 24852 8727 24853
rect 8661 24850 8708 24852
rect 8616 24848 8708 24850
rect 8616 24792 8666 24848
rect 8616 24790 8708 24792
rect 8661 24788 8708 24790
rect 8772 24788 8778 24852
rect 10593 24850 10659 24853
rect 15285 24850 15351 24853
rect 15745 24852 15811 24853
rect 15694 24850 15700 24852
rect 10593 24848 15351 24850
rect 10593 24792 10598 24848
rect 10654 24792 15290 24848
rect 15346 24792 15351 24848
rect 10593 24790 15351 24792
rect 15654 24790 15700 24850
rect 15764 24848 15811 24852
rect 15806 24792 15811 24848
rect 8661 24787 8727 24788
rect 10593 24787 10659 24790
rect 15285 24787 15351 24790
rect 15694 24788 15700 24790
rect 15764 24788 15811 24792
rect 15745 24787 15811 24788
rect 19241 24850 19307 24853
rect 20118 24850 20178 24926
rect 19241 24848 20178 24850
rect 19241 24792 19246 24848
rect 19302 24792 20178 24848
rect 19241 24790 20178 24792
rect 20253 24850 20319 24853
rect 20662 24850 20668 24852
rect 20253 24848 20668 24850
rect 20253 24792 20258 24848
rect 20314 24792 20668 24848
rect 20253 24790 20668 24792
rect 19241 24787 19307 24790
rect 20253 24787 20319 24790
rect 20662 24788 20668 24790
rect 20732 24788 20738 24852
rect 20854 24850 20914 24926
rect 32254 24850 32260 24852
rect 20854 24790 32260 24850
rect 32254 24788 32260 24790
rect 32324 24788 32330 24852
rect 4153 24714 4219 24717
rect 10961 24714 11027 24717
rect 26785 24714 26851 24717
rect 4153 24712 11027 24714
rect 4153 24656 4158 24712
rect 4214 24656 10966 24712
rect 11022 24656 11027 24712
rect 4153 24654 11027 24656
rect 4153 24651 4219 24654
rect 10961 24651 11027 24654
rect 12390 24712 26851 24714
rect 12390 24656 26790 24712
rect 26846 24656 26851 24712
rect 12390 24654 26851 24656
rect 1710 24516 1716 24580
rect 1780 24578 1786 24580
rect 2405 24578 2471 24581
rect 1780 24576 2471 24578
rect 1780 24520 2410 24576
rect 2466 24520 2471 24576
rect 1780 24518 2471 24520
rect 1780 24516 1786 24518
rect 2405 24515 2471 24518
rect 5390 24516 5396 24580
rect 5460 24578 5466 24580
rect 9949 24578 10015 24581
rect 12390 24578 12450 24654
rect 26785 24651 26851 24654
rect 5460 24576 12450 24578
rect 5460 24520 9954 24576
rect 10010 24520 12450 24576
rect 5460 24518 12450 24520
rect 15285 24578 15351 24581
rect 20846 24578 20852 24580
rect 15285 24576 20852 24578
rect 15285 24520 15290 24576
rect 15346 24520 20852 24576
rect 15285 24518 20852 24520
rect 5460 24516 5466 24518
rect 9949 24515 10015 24518
rect 15285 24515 15351 24518
rect 20846 24516 20852 24518
rect 20916 24516 20922 24580
rect 4208 24512 4528 24513
rect 0 24442 800 24472
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 4061 24442 4127 24445
rect 0 24440 4127 24442
rect 0 24384 4066 24440
rect 4122 24384 4127 24440
rect 0 24382 4127 24384
rect 0 24352 800 24382
rect 4061 24379 4127 24382
rect 10910 24380 10916 24444
rect 10980 24442 10986 24444
rect 21766 24442 21772 24444
rect 10980 24382 21772 24442
rect 10980 24380 10986 24382
rect 21766 24380 21772 24382
rect 21836 24380 21842 24444
rect 10041 24306 10107 24309
rect 13629 24306 13695 24309
rect 10041 24304 13695 24306
rect 10041 24248 10046 24304
rect 10102 24248 13634 24304
rect 13690 24248 13695 24304
rect 10041 24246 13695 24248
rect 10041 24243 10107 24246
rect 13629 24243 13695 24246
rect 9213 24170 9279 24173
rect 20294 24170 20300 24172
rect 9213 24168 20300 24170
rect 9213 24112 9218 24168
rect 9274 24112 20300 24168
rect 9213 24110 20300 24112
rect 9213 24107 9279 24110
rect 20294 24108 20300 24110
rect 20364 24108 20370 24172
rect 2262 23972 2268 24036
rect 2332 24034 2338 24036
rect 2405 24034 2471 24037
rect 8293 24034 8359 24037
rect 10133 24036 10199 24037
rect 10133 24034 10180 24036
rect 2332 24032 8359 24034
rect 2332 23976 2410 24032
rect 2466 23976 8298 24032
rect 8354 23976 8359 24032
rect 2332 23974 8359 23976
rect 10088 24032 10180 24034
rect 10088 23976 10138 24032
rect 10088 23974 10180 23976
rect 2332 23972 2338 23974
rect 2405 23971 2471 23974
rect 8293 23971 8359 23974
rect 10133 23972 10180 23974
rect 10244 23972 10250 24036
rect 10133 23971 10199 23972
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 2865 23900 2931 23901
rect 2814 23836 2820 23900
rect 2884 23898 2931 23900
rect 4981 23898 5047 23901
rect 5758 23898 5764 23900
rect 2884 23896 2976 23898
rect 2926 23840 2976 23896
rect 2884 23838 2976 23840
rect 4981 23896 5764 23898
rect 4981 23840 4986 23896
rect 5042 23840 5764 23896
rect 4981 23838 5764 23840
rect 2884 23836 2931 23838
rect 2865 23835 2931 23836
rect 4981 23835 5047 23838
rect 5758 23836 5764 23838
rect 5828 23836 5834 23900
rect 10409 23898 10475 23901
rect 10542 23898 10548 23900
rect 10409 23896 10548 23898
rect 10409 23840 10414 23896
rect 10470 23840 10548 23896
rect 10409 23838 10548 23840
rect 10409 23835 10475 23838
rect 10542 23836 10548 23838
rect 10612 23836 10618 23900
rect 14273 23898 14339 23901
rect 18045 23898 18111 23901
rect 14273 23896 18111 23898
rect 14273 23840 14278 23896
rect 14334 23840 18050 23896
rect 18106 23840 18111 23896
rect 14273 23838 18111 23840
rect 14273 23835 14339 23838
rect 18045 23835 18111 23838
rect 0 23762 800 23792
rect 1485 23762 1551 23765
rect 0 23760 1551 23762
rect 0 23704 1490 23760
rect 1546 23704 1551 23760
rect 0 23702 1551 23704
rect 0 23672 800 23702
rect 1485 23699 1551 23702
rect 10041 23762 10107 23765
rect 17166 23762 17172 23764
rect 10041 23760 17172 23762
rect 10041 23704 10046 23760
rect 10102 23704 17172 23760
rect 10041 23702 17172 23704
rect 10041 23699 10107 23702
rect 17166 23700 17172 23702
rect 17236 23700 17242 23764
rect 24393 23762 24459 23765
rect 17358 23760 24459 23762
rect 17358 23704 24398 23760
rect 24454 23704 24459 23760
rect 17358 23702 24459 23704
rect 5625 23626 5691 23629
rect 982 23624 5691 23626
rect 982 23568 5630 23624
rect 5686 23568 5691 23624
rect 982 23566 5691 23568
rect 841 23490 907 23493
rect 982 23490 1042 23566
rect 5625 23563 5691 23566
rect 6637 23628 6703 23629
rect 6637 23624 6684 23628
rect 6748 23626 6754 23628
rect 6637 23568 6642 23624
rect 6637 23564 6684 23568
rect 6748 23566 6794 23626
rect 6748 23564 6754 23566
rect 7782 23564 7788 23628
rect 7852 23626 7858 23628
rect 12893 23626 12959 23629
rect 7852 23624 12959 23626
rect 7852 23568 12898 23624
rect 12954 23568 12959 23624
rect 7852 23566 12959 23568
rect 7852 23564 7858 23566
rect 6637 23563 6703 23564
rect 12893 23563 12959 23566
rect 13537 23626 13603 23629
rect 17358 23626 17418 23702
rect 24393 23699 24459 23702
rect 13537 23624 17418 23626
rect 13537 23568 13542 23624
rect 13598 23568 17418 23624
rect 13537 23566 17418 23568
rect 19333 23626 19399 23629
rect 25078 23626 25084 23628
rect 19333 23624 25084 23626
rect 19333 23568 19338 23624
rect 19394 23568 25084 23624
rect 19333 23566 25084 23568
rect 13537 23563 13603 23566
rect 19333 23563 19399 23566
rect 25078 23564 25084 23566
rect 25148 23564 25154 23628
rect 841 23488 1042 23490
rect 841 23432 846 23488
rect 902 23432 1042 23488
rect 841 23430 1042 23432
rect 841 23427 907 23430
rect 1526 23428 1532 23492
rect 1596 23490 1602 23492
rect 2037 23490 2103 23493
rect 1596 23488 2103 23490
rect 1596 23432 2042 23488
rect 2098 23432 2103 23488
rect 1596 23430 2103 23432
rect 1596 23428 1602 23430
rect 2037 23427 2103 23430
rect 2957 23490 3023 23493
rect 4061 23490 4127 23493
rect 2957 23488 4127 23490
rect 2957 23432 2962 23488
rect 3018 23432 4066 23488
rect 4122 23432 4127 23488
rect 2957 23430 4127 23432
rect 2957 23427 3023 23430
rect 4061 23427 4127 23430
rect 4705 23490 4771 23493
rect 4838 23490 4844 23492
rect 4705 23488 4844 23490
rect 4705 23432 4710 23488
rect 4766 23432 4844 23488
rect 4705 23430 4844 23432
rect 4705 23427 4771 23430
rect 4838 23428 4844 23430
rect 4908 23428 4914 23492
rect 5165 23490 5231 23493
rect 6545 23490 6611 23493
rect 5165 23488 6611 23490
rect 5165 23432 5170 23488
rect 5226 23432 6550 23488
rect 6606 23432 6611 23488
rect 5165 23430 6611 23432
rect 5165 23427 5231 23430
rect 6545 23427 6611 23430
rect 7598 23428 7604 23492
rect 7668 23490 7674 23492
rect 7925 23490 7991 23493
rect 7668 23488 7991 23490
rect 7668 23432 7930 23488
rect 7986 23432 7991 23488
rect 7668 23430 7991 23432
rect 7668 23428 7674 23430
rect 7925 23427 7991 23430
rect 9254 23428 9260 23492
rect 9324 23490 9330 23492
rect 10501 23490 10567 23493
rect 9324 23488 10567 23490
rect 9324 23432 10506 23488
rect 10562 23432 10567 23488
rect 9324 23430 10567 23432
rect 9324 23428 9330 23430
rect 10501 23427 10567 23430
rect 12341 23490 12407 23493
rect 16849 23492 16915 23493
rect 12566 23490 12572 23492
rect 12341 23488 12572 23490
rect 12341 23432 12346 23488
rect 12402 23432 12572 23488
rect 12341 23430 12572 23432
rect 12341 23427 12407 23430
rect 12566 23428 12572 23430
rect 12636 23428 12642 23492
rect 16798 23428 16804 23492
rect 16868 23490 16915 23492
rect 16868 23488 16960 23490
rect 16910 23432 16960 23488
rect 16868 23430 16960 23432
rect 16868 23428 16915 23430
rect 17534 23428 17540 23492
rect 17604 23490 17610 23492
rect 17861 23490 17927 23493
rect 17604 23488 17927 23490
rect 17604 23432 17866 23488
rect 17922 23432 17927 23488
rect 17604 23430 17927 23432
rect 17604 23428 17610 23430
rect 16849 23427 16915 23428
rect 17861 23427 17927 23430
rect 18505 23490 18571 23493
rect 18689 23490 18755 23493
rect 21173 23490 21239 23493
rect 18505 23488 21239 23490
rect 18505 23432 18510 23488
rect 18566 23432 18694 23488
rect 18750 23432 21178 23488
rect 21234 23432 21239 23488
rect 18505 23430 21239 23432
rect 18505 23427 18571 23430
rect 18689 23427 18755 23430
rect 21173 23427 21239 23430
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 11605 23354 11671 23357
rect 12157 23354 12223 23357
rect 32121 23354 32187 23357
rect 11605 23352 32187 23354
rect 11605 23296 11610 23352
rect 11666 23296 12162 23352
rect 12218 23296 32126 23352
rect 32182 23296 32187 23352
rect 11605 23294 32187 23296
rect 11605 23291 11671 23294
rect 12157 23291 12223 23294
rect 32121 23291 32187 23294
rect 0 23218 800 23248
rect 0 23158 2790 23218
rect 0 23128 800 23158
rect 2730 23082 2790 23158
rect 3918 23156 3924 23220
rect 3988 23218 3994 23220
rect 4889 23218 4955 23221
rect 3988 23216 4955 23218
rect 3988 23160 4894 23216
rect 4950 23160 4955 23216
rect 3988 23158 4955 23160
rect 3988 23156 3994 23158
rect 4889 23155 4955 23158
rect 5533 23218 5599 23221
rect 8753 23218 8819 23221
rect 18045 23220 18111 23221
rect 18045 23218 18092 23220
rect 5533 23216 8819 23218
rect 5533 23160 5538 23216
rect 5594 23160 8758 23216
rect 8814 23160 8819 23216
rect 5533 23158 8819 23160
rect 18000 23216 18092 23218
rect 18000 23160 18050 23216
rect 18000 23158 18092 23160
rect 5533 23155 5599 23158
rect 8753 23155 8819 23158
rect 18045 23156 18092 23158
rect 18156 23156 18162 23220
rect 18505 23218 18571 23221
rect 25497 23218 25563 23221
rect 18505 23216 25563 23218
rect 18505 23160 18510 23216
rect 18566 23160 25502 23216
rect 25558 23160 25563 23216
rect 18505 23158 25563 23160
rect 18045 23155 18111 23156
rect 18505 23155 18571 23158
rect 25497 23155 25563 23158
rect 10726 23082 10732 23084
rect 2730 23022 10732 23082
rect 10726 23020 10732 23022
rect 10796 23020 10802 23084
rect 13118 23020 13124 23084
rect 13188 23082 13194 23084
rect 22185 23082 22251 23085
rect 13188 23080 22251 23082
rect 13188 23024 22190 23080
rect 22246 23024 22251 23080
rect 13188 23022 22251 23024
rect 13188 23020 13194 23022
rect 22185 23019 22251 23022
rect 3969 22948 4035 22949
rect 3918 22884 3924 22948
rect 3988 22946 4035 22948
rect 9029 22946 9095 22949
rect 9438 22946 9444 22948
rect 3988 22944 4080 22946
rect 4030 22888 4080 22944
rect 3988 22886 4080 22888
rect 9029 22944 9444 22946
rect 9029 22888 9034 22944
rect 9090 22888 9444 22944
rect 9029 22886 9444 22888
rect 3988 22884 4035 22886
rect 3969 22883 4035 22884
rect 9029 22883 9095 22886
rect 9438 22884 9444 22886
rect 9508 22884 9514 22948
rect 10225 22946 10291 22949
rect 10358 22946 10364 22948
rect 10225 22944 10364 22946
rect 10225 22888 10230 22944
rect 10286 22888 10364 22944
rect 10225 22886 10364 22888
rect 10225 22883 10291 22886
rect 10358 22884 10364 22886
rect 10428 22884 10434 22948
rect 12341 22946 12407 22949
rect 12525 22946 12591 22949
rect 12341 22944 12591 22946
rect 12341 22888 12346 22944
rect 12402 22888 12530 22944
rect 12586 22888 12591 22944
rect 12341 22886 12591 22888
rect 12341 22883 12407 22886
rect 12525 22883 12591 22886
rect 13486 22884 13492 22948
rect 13556 22946 13562 22948
rect 19241 22946 19307 22949
rect 13556 22944 19307 22946
rect 13556 22888 19246 22944
rect 19302 22888 19307 22944
rect 13556 22886 19307 22888
rect 13556 22884 13562 22886
rect 19241 22883 19307 22886
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 1485 22810 1551 22813
rect 6177 22810 6243 22813
rect 1485 22808 6243 22810
rect 1485 22752 1490 22808
rect 1546 22752 6182 22808
rect 6238 22752 6243 22808
rect 1485 22750 6243 22752
rect 1485 22747 1551 22750
rect 6177 22747 6243 22750
rect 7414 22748 7420 22812
rect 7484 22810 7490 22812
rect 13445 22810 13511 22813
rect 15837 22812 15903 22813
rect 15837 22810 15884 22812
rect 7484 22808 13511 22810
rect 7484 22752 13450 22808
rect 13506 22752 13511 22808
rect 7484 22750 13511 22752
rect 15792 22808 15884 22810
rect 15792 22752 15842 22808
rect 15792 22750 15884 22752
rect 7484 22748 7490 22750
rect 13445 22747 13511 22750
rect 15837 22748 15884 22750
rect 15948 22748 15954 22812
rect 16205 22810 16271 22813
rect 18505 22810 18571 22813
rect 16205 22808 18571 22810
rect 16205 22752 16210 22808
rect 16266 22752 18510 22808
rect 18566 22752 18571 22808
rect 16205 22750 18571 22752
rect 15837 22747 15903 22748
rect 16205 22747 16271 22750
rect 18505 22747 18571 22750
rect 0 22674 800 22704
rect 1393 22674 1459 22677
rect 0 22672 1459 22674
rect 0 22616 1398 22672
rect 1454 22616 1459 22672
rect 0 22614 1459 22616
rect 0 22584 800 22614
rect 1393 22611 1459 22614
rect 9070 22612 9076 22676
rect 9140 22674 9146 22676
rect 10409 22674 10475 22677
rect 9140 22672 10475 22674
rect 9140 22616 10414 22672
rect 10470 22616 10475 22672
rect 9140 22614 10475 22616
rect 9140 22612 9146 22614
rect 10409 22611 10475 22614
rect 10777 22674 10843 22677
rect 11329 22676 11395 22677
rect 11094 22674 11100 22676
rect 10777 22672 11100 22674
rect 10777 22616 10782 22672
rect 10838 22616 11100 22672
rect 10777 22614 11100 22616
rect 10777 22611 10843 22614
rect 11094 22612 11100 22614
rect 11164 22612 11170 22676
rect 11278 22674 11284 22676
rect 11238 22614 11284 22674
rect 11348 22672 11395 22676
rect 19885 22674 19951 22677
rect 11390 22616 11395 22672
rect 11278 22612 11284 22614
rect 11348 22612 11395 22616
rect 11329 22611 11395 22612
rect 12390 22672 19951 22674
rect 12390 22616 19890 22672
rect 19946 22616 19951 22672
rect 12390 22614 19951 22616
rect 6269 22538 6335 22541
rect 9673 22538 9739 22541
rect 6269 22536 9739 22538
rect 6269 22480 6274 22536
rect 6330 22480 9678 22536
rect 9734 22480 9739 22536
rect 6269 22478 9739 22480
rect 6269 22475 6335 22478
rect 9673 22475 9739 22478
rect 10317 22540 10383 22541
rect 10317 22536 10364 22540
rect 10428 22538 10434 22540
rect 10317 22480 10322 22536
rect 10317 22476 10364 22480
rect 10428 22478 10474 22538
rect 10428 22476 10434 22478
rect 10317 22475 10383 22476
rect 8886 22340 8892 22404
rect 8956 22402 8962 22404
rect 9254 22402 9260 22404
rect 8956 22342 9260 22402
rect 8956 22340 8962 22342
rect 9254 22340 9260 22342
rect 9324 22340 9330 22404
rect 9438 22340 9444 22404
rect 9508 22402 9514 22404
rect 12390 22402 12450 22614
rect 19885 22611 19951 22614
rect 13169 22538 13235 22541
rect 13905 22538 13971 22541
rect 13169 22536 13971 22538
rect 13169 22480 13174 22536
rect 13230 22480 13910 22536
rect 13966 22480 13971 22536
rect 13169 22478 13971 22480
rect 13169 22475 13235 22478
rect 13905 22475 13971 22478
rect 17350 22476 17356 22540
rect 17420 22538 17426 22540
rect 19333 22538 19399 22541
rect 17420 22536 19399 22538
rect 17420 22480 19338 22536
rect 19394 22480 19399 22536
rect 17420 22478 19399 22480
rect 17420 22476 17426 22478
rect 19333 22475 19399 22478
rect 9508 22342 12450 22402
rect 13077 22402 13143 22405
rect 16205 22402 16271 22405
rect 13077 22400 16271 22402
rect 13077 22344 13082 22400
rect 13138 22344 16210 22400
rect 16266 22344 16271 22400
rect 13077 22342 16271 22344
rect 9508 22340 9514 22342
rect 13077 22339 13143 22342
rect 16205 22339 16271 22342
rect 18137 22402 18203 22405
rect 18270 22402 18276 22404
rect 18137 22400 18276 22402
rect 18137 22344 18142 22400
rect 18198 22344 18276 22400
rect 18137 22342 18276 22344
rect 18137 22339 18203 22342
rect 18270 22340 18276 22342
rect 18340 22340 18346 22404
rect 21357 22402 21423 22405
rect 30414 22402 30420 22404
rect 21357 22400 30420 22402
rect 21357 22344 21362 22400
rect 21418 22344 30420 22400
rect 21357 22342 30420 22344
rect 21357 22339 21423 22342
rect 30414 22340 30420 22342
rect 30484 22340 30490 22404
rect 30557 22402 30623 22405
rect 30782 22402 30788 22404
rect 30557 22400 30788 22402
rect 30557 22344 30562 22400
rect 30618 22344 30788 22400
rect 30557 22342 30788 22344
rect 30557 22339 30623 22342
rect 30782 22340 30788 22342
rect 30852 22340 30858 22404
rect 31293 22402 31359 22405
rect 31518 22402 31524 22404
rect 31293 22400 31524 22402
rect 31293 22344 31298 22400
rect 31354 22344 31524 22400
rect 31293 22342 31524 22344
rect 31293 22339 31359 22342
rect 31518 22340 31524 22342
rect 31588 22340 31594 22404
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 5165 22266 5231 22269
rect 10133 22266 10199 22269
rect 14825 22266 14891 22269
rect 5165 22264 7482 22266
rect 5165 22208 5170 22264
rect 5226 22208 7482 22264
rect 5165 22206 7482 22208
rect 5165 22203 5231 22206
rect 3049 22130 3115 22133
rect 7189 22130 7255 22133
rect 3049 22128 7255 22130
rect 3049 22072 3054 22128
rect 3110 22072 7194 22128
rect 7250 22072 7255 22128
rect 3049 22070 7255 22072
rect 7422 22130 7482 22206
rect 10133 22264 14891 22266
rect 10133 22208 10138 22264
rect 10194 22208 14830 22264
rect 14886 22208 14891 22264
rect 10133 22206 14891 22208
rect 10133 22203 10199 22206
rect 14825 22203 14891 22206
rect 15837 22266 15903 22269
rect 16297 22266 16363 22269
rect 22001 22266 22067 22269
rect 15837 22264 22067 22266
rect 15837 22208 15842 22264
rect 15898 22208 16302 22264
rect 16358 22208 22006 22264
rect 22062 22208 22067 22264
rect 15837 22206 22067 22208
rect 15837 22203 15903 22206
rect 16297 22203 16363 22206
rect 22001 22203 22067 22206
rect 10225 22130 10291 22133
rect 7422 22128 10291 22130
rect 7422 22072 10230 22128
rect 10286 22072 10291 22128
rect 7422 22070 10291 22072
rect 3049 22067 3115 22070
rect 7189 22067 7255 22070
rect 10225 22067 10291 22070
rect 10777 22130 10843 22133
rect 11053 22130 11119 22133
rect 12433 22130 12499 22133
rect 27654 22130 27660 22132
rect 10777 22128 11119 22130
rect 10777 22072 10782 22128
rect 10838 22072 11058 22128
rect 11114 22072 11119 22128
rect 10777 22070 11119 22072
rect 10777 22067 10843 22070
rect 11053 22067 11119 22070
rect 12022 22128 27660 22130
rect 12022 22072 12438 22128
rect 12494 22072 27660 22128
rect 12022 22070 27660 22072
rect 0 21994 800 22024
rect 0 21934 6930 21994
rect 0 21904 800 21934
rect 3601 21860 3667 21861
rect 3550 21858 3556 21860
rect 3510 21798 3556 21858
rect 3620 21856 3667 21860
rect 3662 21800 3667 21856
rect 3550 21796 3556 21798
rect 3620 21796 3667 21800
rect 6494 21796 6500 21860
rect 6564 21858 6570 21860
rect 6637 21858 6703 21861
rect 6564 21856 6703 21858
rect 6564 21800 6642 21856
rect 6698 21800 6703 21856
rect 6564 21798 6703 21800
rect 6870 21858 6930 21934
rect 7046 21932 7052 21996
rect 7116 21994 7122 21996
rect 7925 21994 7991 21997
rect 7116 21992 7991 21994
rect 7116 21936 7930 21992
rect 7986 21936 7991 21992
rect 7116 21934 7991 21936
rect 7116 21932 7122 21934
rect 7925 21931 7991 21934
rect 10174 21932 10180 21996
rect 10244 21994 10250 21996
rect 10317 21994 10383 21997
rect 10244 21992 10383 21994
rect 10244 21936 10322 21992
rect 10378 21936 10383 21992
rect 10244 21934 10383 21936
rect 10244 21932 10250 21934
rect 10317 21931 10383 21934
rect 10726 21932 10732 21996
rect 10796 21994 10802 21996
rect 12022 21994 12082 22070
rect 12433 22067 12499 22070
rect 27654 22068 27660 22070
rect 27724 22068 27730 22132
rect 10796 21934 12082 21994
rect 12893 21994 12959 21997
rect 14549 21994 14615 21997
rect 12893 21992 14615 21994
rect 12893 21936 12898 21992
rect 12954 21936 14554 21992
rect 14610 21936 14615 21992
rect 12893 21934 14615 21936
rect 10796 21932 10802 21934
rect 12893 21931 12959 21934
rect 14549 21931 14615 21934
rect 16849 21994 16915 21997
rect 16982 21994 16988 21996
rect 16849 21992 16988 21994
rect 16849 21936 16854 21992
rect 16910 21936 16988 21992
rect 16849 21934 16988 21936
rect 16849 21931 16915 21934
rect 16982 21932 16988 21934
rect 17052 21932 17058 21996
rect 31937 21994 32003 21997
rect 17174 21992 32003 21994
rect 17174 21936 31942 21992
rect 31998 21936 32003 21992
rect 17174 21934 32003 21936
rect 9029 21858 9095 21861
rect 6870 21856 9095 21858
rect 6870 21800 9034 21856
rect 9090 21800 9095 21856
rect 6870 21798 9095 21800
rect 6564 21796 6570 21798
rect 3601 21795 3667 21796
rect 6637 21795 6703 21798
rect 9029 21795 9095 21798
rect 11881 21858 11947 21861
rect 17174 21858 17234 21934
rect 31937 21931 32003 21934
rect 11881 21856 17234 21858
rect 11881 21800 11886 21856
rect 11942 21800 17234 21856
rect 11881 21798 17234 21800
rect 17401 21858 17467 21861
rect 17718 21858 17724 21860
rect 17401 21856 17724 21858
rect 17401 21800 17406 21856
rect 17462 21800 17724 21856
rect 17401 21798 17724 21800
rect 11881 21795 11947 21798
rect 17401 21795 17467 21798
rect 17718 21796 17724 21798
rect 17788 21796 17794 21860
rect 18638 21796 18644 21860
rect 18708 21858 18714 21860
rect 19241 21858 19307 21861
rect 18708 21856 19307 21858
rect 18708 21800 19246 21856
rect 19302 21800 19307 21856
rect 18708 21798 19307 21800
rect 18708 21796 18714 21798
rect 19241 21795 19307 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 1945 21722 2011 21725
rect 5349 21722 5415 21725
rect 1945 21720 5415 21722
rect 1945 21664 1950 21720
rect 2006 21664 5354 21720
rect 5410 21664 5415 21720
rect 1945 21662 5415 21664
rect 1945 21659 2011 21662
rect 5349 21659 5415 21662
rect 13169 21722 13235 21725
rect 13302 21722 13308 21724
rect 13169 21720 13308 21722
rect 13169 21664 13174 21720
rect 13230 21664 13308 21720
rect 13169 21662 13308 21664
rect 13169 21659 13235 21662
rect 13302 21660 13308 21662
rect 13372 21660 13378 21724
rect 13445 21722 13511 21725
rect 13445 21720 15026 21722
rect 13445 21664 13450 21720
rect 13506 21664 15026 21720
rect 13445 21662 15026 21664
rect 13445 21659 13511 21662
rect 4797 21586 4863 21589
rect 5022 21586 5028 21588
rect 4797 21584 5028 21586
rect 4797 21528 4802 21584
rect 4858 21528 5028 21584
rect 4797 21526 5028 21528
rect 4797 21523 4863 21526
rect 5022 21524 5028 21526
rect 5092 21524 5098 21588
rect 11697 21586 11763 21589
rect 14089 21586 14155 21589
rect 11697 21584 14155 21586
rect 11697 21528 11702 21584
rect 11758 21528 14094 21584
rect 14150 21528 14155 21584
rect 11697 21526 14155 21528
rect 11697 21523 11763 21526
rect 14089 21523 14155 21526
rect 14641 21586 14707 21589
rect 14774 21586 14780 21588
rect 14641 21584 14780 21586
rect 14641 21528 14646 21584
rect 14702 21528 14780 21584
rect 14641 21526 14780 21528
rect 14641 21523 14707 21526
rect 14774 21524 14780 21526
rect 14844 21524 14850 21588
rect 14966 21586 15026 21662
rect 31886 21586 31892 21588
rect 14966 21526 31892 21586
rect 31886 21524 31892 21526
rect 31956 21524 31962 21588
rect 0 21450 800 21480
rect 2865 21450 2931 21453
rect 0 21448 2931 21450
rect 0 21392 2870 21448
rect 2926 21392 2931 21448
rect 0 21390 2931 21392
rect 0 21360 800 21390
rect 2865 21387 2931 21390
rect 5441 21450 5507 21453
rect 10777 21450 10843 21453
rect 5441 21448 10843 21450
rect 5441 21392 5446 21448
rect 5502 21392 10782 21448
rect 10838 21392 10843 21448
rect 5441 21390 10843 21392
rect 5441 21387 5507 21390
rect 10777 21387 10843 21390
rect 13169 21450 13235 21453
rect 15878 21450 15884 21452
rect 13169 21448 15884 21450
rect 13169 21392 13174 21448
rect 13230 21392 15884 21448
rect 13169 21390 15884 21392
rect 13169 21387 13235 21390
rect 15878 21388 15884 21390
rect 15948 21388 15954 21452
rect 16246 21388 16252 21452
rect 16316 21450 16322 21452
rect 23473 21450 23539 21453
rect 24526 21450 24532 21452
rect 16316 21390 22110 21450
rect 16316 21388 16322 21390
rect 12750 21252 12756 21316
rect 12820 21314 12826 21316
rect 13169 21314 13235 21317
rect 18321 21314 18387 21317
rect 12820 21312 13235 21314
rect 12820 21256 13174 21312
rect 13230 21256 13235 21312
rect 12820 21254 13235 21256
rect 12820 21252 12826 21254
rect 13169 21251 13235 21254
rect 15702 21312 18387 21314
rect 15702 21256 18326 21312
rect 18382 21256 18387 21312
rect 15702 21254 18387 21256
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 565 21178 631 21181
rect 3877 21178 3943 21181
rect 565 21176 3943 21178
rect 565 21120 570 21176
rect 626 21120 3882 21176
rect 3938 21120 3943 21176
rect 565 21118 3943 21120
rect 565 21115 631 21118
rect 3877 21115 3943 21118
rect 9765 21178 9831 21181
rect 14365 21178 14431 21181
rect 9765 21176 14431 21178
rect 9765 21120 9770 21176
rect 9826 21120 14370 21176
rect 14426 21120 14431 21176
rect 9765 21118 14431 21120
rect 9765 21115 9831 21118
rect 14365 21115 14431 21118
rect 2589 21042 2655 21045
rect 3877 21042 3943 21045
rect 2589 21040 3943 21042
rect 2589 20984 2594 21040
rect 2650 20984 3882 21040
rect 3938 20984 3943 21040
rect 2589 20982 3943 20984
rect 2589 20979 2655 20982
rect 3877 20979 3943 20982
rect 4245 21042 4311 21045
rect 4654 21042 4660 21044
rect 4245 21040 4660 21042
rect 4245 20984 4250 21040
rect 4306 20984 4660 21040
rect 4245 20982 4660 20984
rect 4245 20979 4311 20982
rect 4654 20980 4660 20982
rect 4724 20980 4730 21044
rect 12014 20980 12020 21044
rect 12084 21042 12090 21044
rect 15702 21042 15762 21254
rect 18321 21251 18387 21254
rect 19793 21314 19859 21317
rect 22050 21314 22110 21390
rect 23473 21448 24532 21450
rect 23473 21392 23478 21448
rect 23534 21392 24532 21448
rect 23473 21390 24532 21392
rect 23473 21387 23539 21390
rect 24526 21388 24532 21390
rect 24596 21388 24602 21452
rect 31661 21450 31727 21453
rect 40769 21450 40835 21453
rect 31661 21448 40835 21450
rect 31661 21392 31666 21448
rect 31722 21392 40774 21448
rect 40830 21392 40835 21448
rect 31661 21390 40835 21392
rect 31661 21387 31727 21390
rect 40769 21387 40835 21390
rect 19793 21312 21834 21314
rect 19793 21256 19798 21312
rect 19854 21256 21834 21312
rect 19793 21254 21834 21256
rect 22050 21254 31770 21314
rect 19793 21251 19859 21254
rect 15837 21178 15903 21181
rect 21633 21178 21699 21181
rect 15837 21176 21699 21178
rect 15837 21120 15842 21176
rect 15898 21120 21638 21176
rect 21694 21120 21699 21176
rect 15837 21118 21699 21120
rect 21774 21178 21834 21254
rect 27102 21178 27108 21180
rect 21774 21118 27108 21178
rect 15837 21115 15903 21118
rect 21633 21115 21699 21118
rect 27102 21116 27108 21118
rect 27172 21116 27178 21180
rect 12084 20982 15762 21042
rect 12084 20980 12090 20982
rect 15878 20980 15884 21044
rect 15948 21042 15954 21044
rect 16246 21042 16252 21044
rect 15948 20982 16252 21042
rect 15948 20980 15954 20982
rect 16246 20980 16252 20982
rect 16316 20980 16322 21044
rect 18045 21042 18111 21045
rect 24158 21042 24164 21044
rect 18045 21040 24164 21042
rect 18045 20984 18050 21040
rect 18106 20984 24164 21040
rect 18045 20982 24164 20984
rect 18045 20979 18111 20982
rect 24158 20980 24164 20982
rect 24228 20980 24234 21044
rect 31710 21042 31770 21254
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 35433 21042 35499 21045
rect 31710 21040 35499 21042
rect 31710 20984 35438 21040
rect 35494 20984 35499 21040
rect 31710 20982 35499 20984
rect 35433 20979 35499 20982
rect 0 20906 800 20936
rect 2865 20906 2931 20909
rect 0 20904 2931 20906
rect 0 20848 2870 20904
rect 2926 20848 2931 20904
rect 0 20846 2931 20848
rect 0 20816 800 20846
rect 2865 20843 2931 20846
rect 3918 20844 3924 20908
rect 3988 20906 3994 20908
rect 4337 20906 4403 20909
rect 3988 20904 4403 20906
rect 3988 20848 4342 20904
rect 4398 20848 4403 20904
rect 3988 20846 4403 20848
rect 3988 20844 3994 20846
rect 4337 20843 4403 20846
rect 5441 20906 5507 20909
rect 12750 20906 12756 20908
rect 5441 20904 12756 20906
rect 5441 20848 5446 20904
rect 5502 20848 12756 20904
rect 5441 20846 12756 20848
rect 5441 20843 5507 20846
rect 12750 20844 12756 20846
rect 12820 20844 12826 20908
rect 16982 20906 16988 20908
rect 12942 20846 16988 20906
rect 974 20708 980 20772
rect 1044 20770 1050 20772
rect 5533 20770 5599 20773
rect 1044 20768 5599 20770
rect 1044 20712 5538 20768
rect 5594 20712 5599 20768
rect 1044 20710 5599 20712
rect 1044 20708 1050 20710
rect 5533 20707 5599 20710
rect 6821 20770 6887 20773
rect 7005 20770 7071 20773
rect 6821 20768 7071 20770
rect 6821 20712 6826 20768
rect 6882 20712 7010 20768
rect 7066 20712 7071 20768
rect 6821 20710 7071 20712
rect 6821 20707 6887 20710
rect 7005 20707 7071 20710
rect 12065 20770 12131 20773
rect 12198 20770 12204 20772
rect 12065 20768 12204 20770
rect 12065 20712 12070 20768
rect 12126 20712 12204 20768
rect 12065 20710 12204 20712
rect 12065 20707 12131 20710
rect 12198 20708 12204 20710
rect 12268 20708 12274 20772
rect 12525 20770 12591 20773
rect 12942 20770 13002 20846
rect 16982 20844 16988 20846
rect 17052 20844 17058 20908
rect 18137 20906 18203 20909
rect 21398 20906 21404 20908
rect 18137 20904 21404 20906
rect 18137 20848 18142 20904
rect 18198 20848 21404 20904
rect 18137 20846 21404 20848
rect 18137 20843 18203 20846
rect 21398 20844 21404 20846
rect 21468 20844 21474 20908
rect 12525 20768 13002 20770
rect 12525 20712 12530 20768
rect 12586 20712 13002 20768
rect 12525 20710 13002 20712
rect 12525 20707 12591 20710
rect 16246 20708 16252 20772
rect 16316 20770 16322 20772
rect 16665 20770 16731 20773
rect 18413 20772 18479 20773
rect 18413 20770 18460 20772
rect 16316 20768 16731 20770
rect 16316 20712 16670 20768
rect 16726 20712 16731 20768
rect 16316 20710 16731 20712
rect 18368 20768 18460 20770
rect 18368 20712 18418 20768
rect 18368 20710 18460 20712
rect 16316 20708 16322 20710
rect 16665 20707 16731 20710
rect 18413 20708 18460 20710
rect 18524 20708 18530 20772
rect 20294 20708 20300 20772
rect 20364 20770 20370 20772
rect 20437 20770 20503 20773
rect 22185 20772 22251 20773
rect 20364 20768 20503 20770
rect 20364 20712 20442 20768
rect 20498 20712 20503 20768
rect 20364 20710 20503 20712
rect 20364 20708 20370 20710
rect 18413 20707 18479 20708
rect 20437 20707 20503 20710
rect 22134 20708 22140 20772
rect 22204 20770 22251 20772
rect 22204 20768 22296 20770
rect 22246 20712 22296 20768
rect 22204 20710 22296 20712
rect 22204 20708 22251 20710
rect 22185 20707 22251 20708
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 657 20634 723 20637
rect 5533 20636 5599 20637
rect 657 20632 2790 20634
rect 657 20576 662 20632
rect 718 20576 2790 20632
rect 657 20574 2790 20576
rect 657 20571 723 20574
rect 2730 20498 2790 20574
rect 5533 20632 5580 20636
rect 5644 20634 5650 20636
rect 8109 20634 8175 20637
rect 14365 20636 14431 20637
rect 15009 20636 15075 20637
rect 15193 20636 15259 20637
rect 10174 20634 10180 20636
rect 5533 20576 5538 20632
rect 5533 20572 5580 20576
rect 5644 20574 5690 20634
rect 8109 20632 10180 20634
rect 8109 20576 8114 20632
rect 8170 20576 10180 20632
rect 8109 20574 10180 20576
rect 5644 20572 5650 20574
rect 5533 20571 5599 20572
rect 8109 20571 8175 20574
rect 10174 20572 10180 20574
rect 10244 20572 10250 20636
rect 14365 20632 14412 20636
rect 14476 20634 14482 20636
rect 14958 20634 14964 20636
rect 14365 20576 14370 20632
rect 14365 20572 14412 20576
rect 14476 20574 14522 20634
rect 14918 20574 14964 20634
rect 15028 20632 15075 20636
rect 15070 20576 15075 20632
rect 14476 20572 14482 20574
rect 14958 20572 14964 20574
rect 15028 20572 15075 20576
rect 15142 20572 15148 20636
rect 15212 20634 15259 20636
rect 15212 20632 15304 20634
rect 15254 20576 15304 20632
rect 15212 20574 15304 20576
rect 15212 20572 15259 20574
rect 16430 20572 16436 20636
rect 16500 20634 16506 20636
rect 18965 20634 19031 20637
rect 16500 20632 19031 20634
rect 16500 20576 18970 20632
rect 19026 20576 19031 20632
rect 16500 20574 19031 20576
rect 16500 20572 16506 20574
rect 14365 20571 14431 20572
rect 15009 20571 15075 20572
rect 15193 20571 15259 20572
rect 18965 20571 19031 20574
rect 22645 20636 22711 20637
rect 28349 20636 28415 20637
rect 22645 20632 22692 20636
rect 22756 20634 22762 20636
rect 28349 20634 28396 20636
rect 22645 20576 22650 20632
rect 22645 20572 22692 20576
rect 22756 20574 22802 20634
rect 28304 20632 28396 20634
rect 28304 20576 28354 20632
rect 28304 20574 28396 20576
rect 22756 20572 22762 20574
rect 28349 20572 28396 20574
rect 28460 20572 28466 20636
rect 22645 20571 22711 20572
rect 28349 20571 28415 20572
rect 5809 20498 5875 20501
rect 2730 20496 5875 20498
rect 2730 20440 5814 20496
rect 5870 20440 5875 20496
rect 2730 20438 5875 20440
rect 5809 20435 5875 20438
rect 8702 20436 8708 20500
rect 8772 20498 8778 20500
rect 8937 20498 9003 20501
rect 8772 20496 9003 20498
rect 8772 20440 8942 20496
rect 8998 20440 9003 20496
rect 8772 20438 9003 20440
rect 8772 20436 8778 20438
rect 8937 20435 9003 20438
rect 10777 20498 10843 20501
rect 16573 20498 16639 20501
rect 19517 20498 19583 20501
rect 10777 20496 16314 20498
rect 10777 20440 10782 20496
rect 10838 20440 16314 20496
rect 10777 20438 16314 20440
rect 10777 20435 10843 20438
rect 0 20362 800 20392
rect 2773 20362 2839 20365
rect 0 20360 2839 20362
rect 0 20304 2778 20360
rect 2834 20304 2839 20360
rect 0 20302 2839 20304
rect 0 20272 800 20302
rect 2773 20299 2839 20302
rect 4521 20362 4587 20365
rect 6637 20364 6703 20365
rect 4838 20362 4844 20364
rect 4521 20360 4844 20362
rect 4521 20304 4526 20360
rect 4582 20304 4844 20360
rect 4521 20302 4844 20304
rect 4521 20299 4587 20302
rect 4838 20300 4844 20302
rect 4908 20300 4914 20364
rect 6637 20362 6684 20364
rect 6556 20360 6684 20362
rect 6748 20362 6754 20364
rect 7649 20362 7715 20365
rect 6748 20360 7715 20362
rect 6556 20304 6642 20360
rect 6748 20304 7654 20360
rect 7710 20304 7715 20360
rect 6556 20302 6684 20304
rect 6637 20300 6684 20302
rect 6748 20302 7715 20304
rect 6748 20300 6754 20302
rect 6637 20299 6703 20300
rect 7649 20299 7715 20302
rect 9254 20300 9260 20364
rect 9324 20362 9330 20364
rect 12566 20362 12572 20364
rect 9324 20302 12572 20362
rect 9324 20300 9330 20302
rect 12566 20300 12572 20302
rect 12636 20300 12642 20364
rect 3693 20226 3759 20229
rect 3558 20224 3759 20226
rect 3558 20168 3698 20224
rect 3754 20168 3759 20224
rect 3558 20166 3759 20168
rect 3233 19818 3299 19821
rect 3558 19818 3618 20166
rect 3693 20163 3759 20166
rect 4613 20226 4679 20229
rect 11830 20226 11836 20228
rect 4613 20224 11836 20226
rect 4613 20168 4618 20224
rect 4674 20168 11836 20224
rect 4613 20166 11836 20168
rect 4613 20163 4679 20166
rect 11830 20164 11836 20166
rect 11900 20164 11906 20228
rect 16254 20226 16314 20438
rect 16573 20496 19583 20498
rect 16573 20440 16578 20496
rect 16634 20440 19522 20496
rect 19578 20440 19583 20496
rect 16573 20438 19583 20440
rect 16573 20435 16639 20438
rect 19517 20435 19583 20438
rect 24485 20498 24551 20501
rect 35525 20498 35591 20501
rect 24485 20496 35591 20498
rect 24485 20440 24490 20496
rect 24546 20440 35530 20496
rect 35586 20440 35591 20496
rect 24485 20438 35591 20440
rect 24485 20435 24551 20438
rect 35525 20435 35591 20438
rect 16481 20362 16547 20365
rect 16481 20360 31770 20362
rect 16481 20304 16486 20360
rect 16542 20304 31770 20360
rect 16481 20302 31770 20304
rect 16481 20299 16547 20302
rect 24209 20226 24275 20229
rect 29085 20228 29151 20229
rect 29085 20226 29132 20228
rect 16254 20224 24275 20226
rect 16254 20168 24214 20224
rect 24270 20168 24275 20224
rect 16254 20166 24275 20168
rect 29040 20224 29132 20226
rect 29040 20168 29090 20224
rect 29040 20166 29132 20168
rect 24209 20163 24275 20166
rect 29085 20164 29132 20166
rect 29196 20164 29202 20228
rect 31710 20226 31770 20302
rect 32581 20226 32647 20229
rect 31710 20224 32647 20226
rect 31710 20168 32586 20224
rect 32642 20168 32647 20224
rect 31710 20166 32647 20168
rect 29085 20163 29151 20164
rect 32581 20163 32647 20166
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 3693 20092 3759 20093
rect 3693 20088 3740 20092
rect 3804 20090 3810 20092
rect 6545 20090 6611 20093
rect 8385 20090 8451 20093
rect 3693 20032 3698 20088
rect 3693 20028 3740 20032
rect 3804 20030 3850 20090
rect 6545 20088 8451 20090
rect 6545 20032 6550 20088
rect 6606 20032 8390 20088
rect 8446 20032 8451 20088
rect 6545 20030 8451 20032
rect 3804 20028 3810 20030
rect 3693 20027 3759 20028
rect 6545 20027 6611 20030
rect 8385 20027 8451 20030
rect 13302 20028 13308 20092
rect 13372 20090 13378 20092
rect 16665 20090 16731 20093
rect 13372 20088 16731 20090
rect 13372 20032 16670 20088
rect 16726 20032 16731 20088
rect 13372 20030 16731 20032
rect 13372 20028 13378 20030
rect 16665 20027 16731 20030
rect 19425 20090 19491 20093
rect 20713 20090 20779 20093
rect 23657 20090 23723 20093
rect 19425 20088 23723 20090
rect 19425 20032 19430 20088
rect 19486 20032 20718 20088
rect 20774 20032 23662 20088
rect 23718 20032 23723 20088
rect 19425 20030 23723 20032
rect 19425 20027 19491 20030
rect 20713 20027 20779 20030
rect 23657 20027 23723 20030
rect 4245 19954 4311 19957
rect 8569 19954 8635 19957
rect 4245 19952 8635 19954
rect 4245 19896 4250 19952
rect 4306 19896 8574 19952
rect 8630 19896 8635 19952
rect 4245 19894 8635 19896
rect 4245 19891 4311 19894
rect 8569 19891 8635 19894
rect 13537 19954 13603 19957
rect 15653 19954 15719 19957
rect 13537 19952 15719 19954
rect 13537 19896 13542 19952
rect 13598 19896 15658 19952
rect 15714 19896 15719 19952
rect 13537 19894 15719 19896
rect 13537 19891 13603 19894
rect 15653 19891 15719 19894
rect 16205 19954 16271 19957
rect 25262 19954 25268 19956
rect 16205 19952 25268 19954
rect 16205 19896 16210 19952
rect 16266 19896 25268 19952
rect 16205 19894 25268 19896
rect 16205 19891 16271 19894
rect 25262 19892 25268 19894
rect 25332 19892 25338 19956
rect 7189 19818 7255 19821
rect 10685 19818 10751 19821
rect 3233 19816 7255 19818
rect 3233 19760 3238 19816
rect 3294 19760 7194 19816
rect 7250 19760 7255 19816
rect 3233 19758 7255 19760
rect 3233 19755 3299 19758
rect 7189 19755 7255 19758
rect 7422 19816 10751 19818
rect 7422 19760 10690 19816
rect 10746 19760 10751 19816
rect 7422 19758 10751 19760
rect 0 19682 800 19712
rect 3325 19682 3391 19685
rect 5349 19682 5415 19685
rect 0 19622 2790 19682
rect 0 19592 800 19622
rect 2730 19546 2790 19622
rect 3325 19680 5415 19682
rect 3325 19624 3330 19680
rect 3386 19624 5354 19680
rect 5410 19624 5415 19680
rect 3325 19622 5415 19624
rect 3325 19619 3391 19622
rect 5349 19619 5415 19622
rect 5574 19620 5580 19684
rect 5644 19682 5650 19684
rect 7422 19682 7482 19758
rect 10685 19755 10751 19758
rect 13537 19818 13603 19821
rect 13670 19818 13676 19820
rect 13537 19816 13676 19818
rect 13537 19760 13542 19816
rect 13598 19760 13676 19816
rect 13537 19758 13676 19760
rect 13537 19755 13603 19758
rect 13670 19756 13676 19758
rect 13740 19756 13746 19820
rect 14958 19756 14964 19820
rect 15028 19818 15034 19820
rect 17125 19818 17191 19821
rect 15028 19816 17191 19818
rect 15028 19760 17130 19816
rect 17186 19760 17191 19816
rect 15028 19758 17191 19760
rect 15028 19756 15034 19758
rect 17125 19755 17191 19758
rect 18137 19818 18203 19821
rect 25814 19818 25820 19820
rect 18137 19816 25820 19818
rect 18137 19760 18142 19816
rect 18198 19760 25820 19816
rect 18137 19758 25820 19760
rect 18137 19755 18203 19758
rect 25814 19756 25820 19758
rect 25884 19756 25890 19820
rect 27613 19818 27679 19821
rect 32070 19818 32076 19820
rect 27613 19816 32076 19818
rect 27613 19760 27618 19816
rect 27674 19760 32076 19816
rect 27613 19758 32076 19760
rect 27613 19755 27679 19758
rect 32070 19756 32076 19758
rect 32140 19756 32146 19820
rect 5644 19622 7482 19682
rect 5644 19620 5650 19622
rect 8150 19620 8156 19684
rect 8220 19682 8226 19684
rect 8661 19682 8727 19685
rect 8220 19680 8727 19682
rect 8220 19624 8666 19680
rect 8722 19624 8727 19680
rect 8220 19622 8727 19624
rect 8220 19620 8226 19622
rect 8661 19619 8727 19622
rect 9673 19682 9739 19685
rect 12801 19682 12867 19685
rect 9673 19680 12867 19682
rect 9673 19624 9678 19680
rect 9734 19624 12806 19680
rect 12862 19624 12867 19680
rect 9673 19622 12867 19624
rect 9673 19619 9739 19622
rect 12801 19619 12867 19622
rect 12985 19682 13051 19685
rect 16113 19682 16179 19685
rect 16481 19682 16547 19685
rect 12985 19680 16547 19682
rect 12985 19624 12990 19680
rect 13046 19624 16118 19680
rect 16174 19624 16486 19680
rect 16542 19624 16547 19680
rect 12985 19622 16547 19624
rect 12985 19619 13051 19622
rect 16113 19619 16179 19622
rect 16481 19619 16547 19622
rect 16614 19620 16620 19684
rect 16684 19682 16690 19684
rect 17217 19682 17283 19685
rect 16684 19680 17283 19682
rect 16684 19624 17222 19680
rect 17278 19624 17283 19680
rect 16684 19622 17283 19624
rect 16684 19620 16690 19622
rect 17217 19619 17283 19622
rect 20621 19682 20687 19685
rect 22318 19682 22324 19684
rect 20621 19680 22324 19682
rect 20621 19624 20626 19680
rect 20682 19624 22324 19680
rect 20621 19622 22324 19624
rect 20621 19619 20687 19622
rect 22318 19620 22324 19622
rect 22388 19620 22394 19684
rect 23473 19682 23539 19685
rect 31385 19684 31451 19685
rect 28942 19682 28948 19684
rect 23473 19680 28948 19682
rect 23473 19624 23478 19680
rect 23534 19624 28948 19680
rect 23473 19622 28948 19624
rect 23473 19619 23539 19622
rect 28942 19620 28948 19622
rect 29012 19620 29018 19684
rect 31334 19620 31340 19684
rect 31404 19682 31451 19684
rect 33777 19682 33843 19685
rect 33910 19682 33916 19684
rect 31404 19680 31496 19682
rect 31446 19624 31496 19680
rect 31404 19622 31496 19624
rect 33777 19680 33916 19682
rect 33777 19624 33782 19680
rect 33838 19624 33916 19680
rect 33777 19622 33916 19624
rect 31404 19620 31451 19622
rect 31385 19619 31451 19620
rect 33777 19619 33843 19622
rect 33910 19620 33916 19622
rect 33980 19620 33986 19684
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 9397 19546 9463 19549
rect 10317 19548 10383 19549
rect 9622 19546 9628 19548
rect 2730 19486 8770 19546
rect 3182 19348 3188 19412
rect 3252 19410 3258 19412
rect 4521 19410 4587 19413
rect 3252 19408 4587 19410
rect 3252 19352 4526 19408
rect 4582 19352 4587 19408
rect 3252 19350 4587 19352
rect 3252 19348 3258 19350
rect 4521 19347 4587 19350
rect 4705 19410 4771 19413
rect 5022 19410 5028 19412
rect 4705 19408 5028 19410
rect 4705 19352 4710 19408
rect 4766 19352 5028 19408
rect 4705 19350 5028 19352
rect 4705 19347 4771 19350
rect 5022 19348 5028 19350
rect 5092 19348 5098 19412
rect 5349 19410 5415 19413
rect 5758 19410 5764 19412
rect 5349 19408 5764 19410
rect 5349 19352 5354 19408
rect 5410 19352 5764 19408
rect 5349 19350 5764 19352
rect 5349 19347 5415 19350
rect 5758 19348 5764 19350
rect 5828 19348 5834 19412
rect 6085 19410 6151 19413
rect 6678 19410 6684 19412
rect 6085 19408 6684 19410
rect 6085 19352 6090 19408
rect 6146 19352 6684 19408
rect 6085 19350 6684 19352
rect 6085 19347 6151 19350
rect 6678 19348 6684 19350
rect 6748 19348 6754 19412
rect 8710 19410 8770 19486
rect 9397 19544 9628 19546
rect 9397 19488 9402 19544
rect 9458 19488 9628 19544
rect 9397 19486 9628 19488
rect 9397 19483 9463 19486
rect 9622 19484 9628 19486
rect 9692 19484 9698 19548
rect 10317 19544 10364 19548
rect 10428 19546 10434 19548
rect 10685 19546 10751 19549
rect 21265 19548 21331 19549
rect 22001 19548 22067 19549
rect 21214 19546 21220 19548
rect 10317 19488 10322 19544
rect 10317 19484 10364 19488
rect 10428 19486 10474 19546
rect 10685 19544 17234 19546
rect 10685 19488 10690 19544
rect 10746 19488 17234 19544
rect 10685 19486 17234 19488
rect 21174 19486 21220 19546
rect 21284 19544 21331 19548
rect 21950 19546 21956 19548
rect 21326 19488 21331 19544
rect 10428 19484 10434 19486
rect 10317 19483 10383 19484
rect 10685 19483 10751 19486
rect 10685 19410 10751 19413
rect 13353 19410 13419 19413
rect 8710 19408 13419 19410
rect 8710 19352 10690 19408
rect 10746 19352 13358 19408
rect 13414 19352 13419 19408
rect 8710 19350 13419 19352
rect 10685 19347 10751 19350
rect 13353 19347 13419 19350
rect 13629 19410 13695 19413
rect 13854 19410 13860 19412
rect 13629 19408 13860 19410
rect 13629 19352 13634 19408
rect 13690 19352 13860 19408
rect 13629 19350 13860 19352
rect 13629 19347 13695 19350
rect 13854 19348 13860 19350
rect 13924 19348 13930 19412
rect 14089 19410 14155 19413
rect 14590 19410 14596 19412
rect 14089 19408 14596 19410
rect 14089 19352 14094 19408
rect 14150 19352 14596 19408
rect 14089 19350 14596 19352
rect 14089 19347 14155 19350
rect 14590 19348 14596 19350
rect 14660 19348 14666 19412
rect 17174 19410 17234 19486
rect 21214 19484 21220 19486
rect 21284 19484 21331 19488
rect 21910 19486 21956 19546
rect 22020 19544 22067 19548
rect 22062 19488 22067 19544
rect 21950 19484 21956 19486
rect 22020 19484 22067 19488
rect 21265 19483 21331 19484
rect 22001 19483 22067 19484
rect 25037 19546 25103 19549
rect 29085 19546 29151 19549
rect 25037 19544 29151 19546
rect 25037 19488 25042 19544
rect 25098 19488 29090 19544
rect 29146 19488 29151 19544
rect 25037 19486 29151 19488
rect 25037 19483 25103 19486
rect 29085 19483 29151 19486
rect 30189 19548 30255 19549
rect 30189 19544 30236 19548
rect 30300 19546 30306 19548
rect 32029 19546 32095 19549
rect 30189 19488 30194 19544
rect 30189 19484 30236 19488
rect 30300 19486 30346 19546
rect 31710 19544 32095 19546
rect 31710 19488 32034 19544
rect 32090 19488 32095 19544
rect 31710 19486 32095 19488
rect 30300 19484 30306 19486
rect 30189 19483 30255 19484
rect 23841 19410 23907 19413
rect 17174 19408 23907 19410
rect 17174 19352 23846 19408
rect 23902 19352 23907 19408
rect 17174 19350 23907 19352
rect 23841 19347 23907 19350
rect 25078 19348 25084 19412
rect 25148 19410 25154 19412
rect 25865 19410 25931 19413
rect 26049 19412 26115 19413
rect 25148 19408 25931 19410
rect 25148 19352 25870 19408
rect 25926 19352 25931 19408
rect 25148 19350 25931 19352
rect 25148 19348 25154 19350
rect 25865 19347 25931 19350
rect 25998 19348 26004 19412
rect 26068 19410 26115 19412
rect 26969 19410 27035 19413
rect 27838 19410 27844 19412
rect 26068 19408 26160 19410
rect 26110 19352 26160 19408
rect 26068 19350 26160 19352
rect 26969 19408 27844 19410
rect 26969 19352 26974 19408
rect 27030 19352 27844 19408
rect 26969 19350 27844 19352
rect 26068 19348 26115 19350
rect 26049 19347 26115 19348
rect 26969 19347 27035 19350
rect 27838 19348 27844 19350
rect 27908 19348 27914 19412
rect 28574 19348 28580 19412
rect 28644 19410 28650 19412
rect 31710 19410 31770 19486
rect 32029 19483 32095 19486
rect 28644 19350 31770 19410
rect 28644 19348 28650 19350
rect 2037 19274 2103 19277
rect 2262 19274 2268 19276
rect 2037 19272 2268 19274
rect 2037 19216 2042 19272
rect 2098 19216 2268 19272
rect 2037 19214 2268 19216
rect 2037 19211 2103 19214
rect 2262 19212 2268 19214
rect 2332 19212 2338 19276
rect 3417 19274 3483 19277
rect 13445 19274 13511 19277
rect 3417 19272 13511 19274
rect 3417 19216 3422 19272
rect 3478 19216 13450 19272
rect 13506 19216 13511 19272
rect 3417 19214 13511 19216
rect 3417 19211 3483 19214
rect 13445 19211 13511 19214
rect 15929 19274 15995 19277
rect 16062 19274 16068 19276
rect 15929 19272 16068 19274
rect 15929 19216 15934 19272
rect 15990 19216 16068 19272
rect 15929 19214 16068 19216
rect 15929 19211 15995 19214
rect 16062 19212 16068 19214
rect 16132 19212 16138 19276
rect 16798 19212 16804 19276
rect 16868 19274 16874 19276
rect 17217 19274 17283 19277
rect 18137 19276 18203 19277
rect 18086 19274 18092 19276
rect 16868 19272 17283 19274
rect 16868 19216 17222 19272
rect 17278 19216 17283 19272
rect 16868 19214 17283 19216
rect 18046 19214 18092 19274
rect 18156 19272 18203 19276
rect 18198 19216 18203 19272
rect 16868 19212 16874 19214
rect 17217 19211 17283 19214
rect 18086 19212 18092 19214
rect 18156 19212 18203 19216
rect 19374 19212 19380 19276
rect 19444 19274 19450 19276
rect 19517 19274 19583 19277
rect 19444 19272 19583 19274
rect 19444 19216 19522 19272
rect 19578 19216 19583 19272
rect 19444 19214 19583 19216
rect 19444 19212 19450 19214
rect 18137 19211 18203 19212
rect 19517 19211 19583 19214
rect 20529 19274 20595 19277
rect 25497 19276 25563 19277
rect 22134 19274 22140 19276
rect 20529 19272 22140 19274
rect 20529 19216 20534 19272
rect 20590 19216 22140 19272
rect 20529 19214 22140 19216
rect 20529 19211 20595 19214
rect 22134 19212 22140 19214
rect 22204 19212 22210 19276
rect 25446 19212 25452 19276
rect 25516 19274 25563 19276
rect 27245 19276 27311 19277
rect 27245 19274 27292 19276
rect 25516 19272 25608 19274
rect 25558 19216 25608 19272
rect 25516 19214 25608 19216
rect 27200 19272 27292 19274
rect 27200 19216 27250 19272
rect 27200 19214 27292 19216
rect 25516 19212 25563 19214
rect 25497 19211 25563 19212
rect 27245 19212 27292 19214
rect 27356 19212 27362 19276
rect 30281 19274 30347 19277
rect 31661 19274 31727 19277
rect 30281 19272 31727 19274
rect 30281 19216 30286 19272
rect 30342 19216 31666 19272
rect 31722 19216 31727 19272
rect 30281 19214 31727 19216
rect 27245 19211 27311 19212
rect 30281 19211 30347 19214
rect 31661 19211 31727 19214
rect 0 19138 800 19168
rect 1761 19138 1827 19141
rect 0 19136 1827 19138
rect 0 19080 1766 19136
rect 1822 19080 1827 19136
rect 0 19078 1827 19080
rect 0 19048 800 19078
rect 1761 19075 1827 19078
rect 11646 19076 11652 19140
rect 11716 19138 11722 19140
rect 14273 19138 14339 19141
rect 11716 19136 14339 19138
rect 11716 19080 14278 19136
rect 14334 19080 14339 19136
rect 11716 19078 14339 19080
rect 11716 19076 11722 19078
rect 14273 19075 14339 19078
rect 15653 19138 15719 19141
rect 19374 19138 19380 19140
rect 15653 19136 19380 19138
rect 15653 19080 15658 19136
rect 15714 19080 19380 19136
rect 15653 19078 19380 19080
rect 15653 19075 15719 19078
rect 19374 19076 19380 19078
rect 19444 19076 19450 19140
rect 19701 19138 19767 19141
rect 20713 19138 20779 19141
rect 19701 19136 20779 19138
rect 19701 19080 19706 19136
rect 19762 19080 20718 19136
rect 20774 19080 20779 19136
rect 19701 19078 20779 19080
rect 19701 19075 19767 19078
rect 20713 19075 20779 19078
rect 24761 19138 24827 19141
rect 28441 19138 28507 19141
rect 24761 19136 28507 19138
rect 24761 19080 24766 19136
rect 24822 19080 28446 19136
rect 28502 19080 28507 19136
rect 24761 19078 28507 19080
rect 24761 19075 24827 19078
rect 28441 19075 28507 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 12566 18940 12572 19004
rect 12636 19002 12642 19004
rect 19149 19002 19215 19005
rect 22502 19002 22508 19004
rect 12636 18942 19074 19002
rect 12636 18940 12642 18942
rect 2037 18866 2103 18869
rect 2814 18866 2820 18868
rect 2037 18864 2820 18866
rect 2037 18808 2042 18864
rect 2098 18808 2820 18864
rect 2037 18806 2820 18808
rect 2037 18803 2103 18806
rect 2814 18804 2820 18806
rect 2884 18804 2890 18868
rect 4521 18866 4587 18869
rect 5441 18866 5507 18869
rect 4521 18864 5507 18866
rect 4521 18808 4526 18864
rect 4582 18808 5446 18864
rect 5502 18808 5507 18864
rect 4521 18806 5507 18808
rect 4521 18803 4587 18806
rect 5441 18803 5507 18806
rect 11329 18866 11395 18869
rect 12157 18866 12223 18869
rect 14089 18866 14155 18869
rect 11329 18864 14155 18866
rect 11329 18808 11334 18864
rect 11390 18808 12162 18864
rect 12218 18808 14094 18864
rect 14150 18808 14155 18864
rect 11329 18806 14155 18808
rect 11329 18803 11395 18806
rect 12157 18803 12223 18806
rect 14089 18803 14155 18806
rect 15193 18866 15259 18869
rect 18873 18866 18939 18869
rect 15193 18864 18939 18866
rect 15193 18808 15198 18864
rect 15254 18808 18878 18864
rect 18934 18808 18939 18864
rect 15193 18806 18939 18808
rect 19014 18866 19074 18942
rect 19149 19000 22508 19002
rect 19149 18944 19154 19000
rect 19210 18944 22508 19000
rect 19149 18942 22508 18944
rect 19149 18939 19215 18942
rect 22502 18940 22508 18942
rect 22572 19002 22578 19004
rect 24945 19002 25011 19005
rect 22572 19000 25011 19002
rect 22572 18944 24950 19000
rect 25006 18944 25011 19000
rect 22572 18942 25011 18944
rect 22572 18940 22578 18942
rect 24945 18939 25011 18942
rect 20437 18866 20503 18869
rect 19014 18864 20503 18866
rect 19014 18808 20442 18864
rect 20498 18808 20503 18864
rect 19014 18806 20503 18808
rect 15193 18803 15259 18806
rect 18873 18803 18939 18806
rect 20437 18803 20503 18806
rect 20662 18804 20668 18868
rect 20732 18866 20738 18868
rect 24945 18866 25011 18869
rect 20732 18864 25011 18866
rect 20732 18808 24950 18864
rect 25006 18808 25011 18864
rect 20732 18806 25011 18808
rect 20732 18804 20738 18806
rect 24945 18803 25011 18806
rect 2998 18668 3004 18732
rect 3068 18730 3074 18732
rect 5942 18730 5948 18732
rect 3068 18670 5948 18730
rect 3068 18668 3074 18670
rect 5942 18668 5948 18670
rect 6012 18668 6018 18732
rect 7281 18730 7347 18733
rect 6088 18728 7347 18730
rect 6088 18672 7286 18728
rect 7342 18672 7347 18728
rect 6088 18670 7347 18672
rect 0 18594 800 18624
rect 3693 18594 3759 18597
rect 0 18592 3759 18594
rect 0 18536 3698 18592
rect 3754 18536 3759 18592
rect 0 18534 3759 18536
rect 0 18504 800 18534
rect 3693 18531 3759 18534
rect 4153 18594 4219 18597
rect 6088 18594 6148 18670
rect 7281 18667 7347 18670
rect 8661 18730 8727 18733
rect 19793 18730 19859 18733
rect 8661 18728 19859 18730
rect 8661 18672 8666 18728
rect 8722 18672 19798 18728
rect 19854 18672 19859 18728
rect 8661 18670 19859 18672
rect 8661 18667 8727 18670
rect 19793 18667 19859 18670
rect 20294 18668 20300 18732
rect 20364 18730 20370 18732
rect 21817 18730 21883 18733
rect 20364 18728 21883 18730
rect 20364 18672 21822 18728
rect 21878 18672 21883 18728
rect 20364 18670 21883 18672
rect 20364 18668 20370 18670
rect 21817 18667 21883 18670
rect 24853 18730 24919 18733
rect 28022 18730 28028 18732
rect 24853 18728 28028 18730
rect 24853 18672 24858 18728
rect 24914 18672 28028 18728
rect 24853 18670 28028 18672
rect 24853 18667 24919 18670
rect 28022 18668 28028 18670
rect 28092 18668 28098 18732
rect 4153 18592 6148 18594
rect 4153 18536 4158 18592
rect 4214 18536 6148 18592
rect 4153 18534 6148 18536
rect 6545 18594 6611 18597
rect 10961 18594 11027 18597
rect 6545 18592 11027 18594
rect 6545 18536 6550 18592
rect 6606 18536 10966 18592
rect 11022 18536 11027 18592
rect 6545 18534 11027 18536
rect 4153 18531 4219 18534
rect 6545 18531 6611 18534
rect 10961 18531 11027 18534
rect 11278 18532 11284 18596
rect 11348 18594 11354 18596
rect 11697 18594 11763 18597
rect 11348 18592 11763 18594
rect 11348 18536 11702 18592
rect 11758 18536 11763 18592
rect 11348 18534 11763 18536
rect 11348 18532 11354 18534
rect 11697 18531 11763 18534
rect 15510 18532 15516 18596
rect 15580 18594 15586 18596
rect 16665 18594 16731 18597
rect 15580 18592 16731 18594
rect 15580 18536 16670 18592
rect 16726 18536 16731 18592
rect 15580 18534 16731 18536
rect 15580 18532 15586 18534
rect 16665 18531 16731 18534
rect 16798 18532 16804 18596
rect 16868 18594 16874 18596
rect 18045 18594 18111 18597
rect 26601 18596 26667 18597
rect 16868 18592 18111 18594
rect 16868 18536 18050 18592
rect 18106 18536 18111 18592
rect 16868 18534 18111 18536
rect 16868 18532 16874 18534
rect 18045 18531 18111 18534
rect 26550 18532 26556 18596
rect 26620 18594 26667 18596
rect 26620 18592 26712 18594
rect 26662 18536 26712 18592
rect 26620 18534 26712 18536
rect 26620 18532 26667 18534
rect 26601 18531 26667 18532
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3141 18458 3207 18461
rect 5206 18458 5212 18460
rect 3141 18456 5212 18458
rect 3141 18400 3146 18456
rect 3202 18400 5212 18456
rect 3141 18398 5212 18400
rect 3141 18395 3207 18398
rect 5206 18396 5212 18398
rect 5276 18396 5282 18460
rect 8937 18458 9003 18461
rect 17125 18458 17191 18461
rect 8937 18456 17191 18458
rect 8937 18400 8942 18456
rect 8998 18400 17130 18456
rect 17186 18400 17191 18456
rect 8937 18398 17191 18400
rect 8937 18395 9003 18398
rect 17125 18395 17191 18398
rect 17769 18458 17835 18461
rect 18873 18458 18939 18461
rect 21449 18458 21515 18461
rect 17769 18456 18939 18458
rect 17769 18400 17774 18456
rect 17830 18400 18878 18456
rect 18934 18400 18939 18456
rect 17769 18398 18939 18400
rect 17769 18395 17835 18398
rect 18873 18395 18939 18398
rect 20118 18456 21515 18458
rect 20118 18400 21454 18456
rect 21510 18400 21515 18456
rect 20118 18398 21515 18400
rect 3969 18322 4035 18325
rect 16021 18322 16087 18325
rect 3969 18320 16087 18322
rect 3969 18264 3974 18320
rect 4030 18264 16026 18320
rect 16082 18264 16087 18320
rect 3969 18262 16087 18264
rect 3969 18259 4035 18262
rect 16021 18259 16087 18262
rect 17217 18322 17283 18325
rect 20118 18322 20178 18398
rect 21449 18395 21515 18398
rect 22921 18458 22987 18461
rect 24894 18458 24900 18460
rect 22921 18456 24900 18458
rect 22921 18400 22926 18456
rect 22982 18400 24900 18456
rect 22921 18398 24900 18400
rect 22921 18395 22987 18398
rect 24894 18396 24900 18398
rect 24964 18396 24970 18460
rect 17217 18320 20178 18322
rect 17217 18264 17222 18320
rect 17278 18264 20178 18320
rect 17217 18262 20178 18264
rect 20345 18322 20411 18325
rect 23197 18322 23263 18325
rect 20345 18320 23263 18322
rect 20345 18264 20350 18320
rect 20406 18264 23202 18320
rect 23258 18264 23263 18320
rect 20345 18262 23263 18264
rect 17217 18259 17283 18262
rect 20345 18259 20411 18262
rect 23197 18259 23263 18262
rect 23381 18322 23447 18325
rect 24894 18322 24900 18324
rect 23381 18320 24900 18322
rect 23381 18264 23386 18320
rect 23442 18264 24900 18320
rect 23381 18262 24900 18264
rect 23381 18259 23447 18262
rect 24894 18260 24900 18262
rect 24964 18260 24970 18324
rect 25497 18322 25563 18325
rect 26734 18322 26740 18324
rect 25497 18320 26740 18322
rect 25497 18264 25502 18320
rect 25558 18264 26740 18320
rect 25497 18262 26740 18264
rect 25497 18259 25563 18262
rect 26734 18260 26740 18262
rect 26804 18260 26810 18324
rect 31661 18322 31727 18325
rect 32254 18322 32260 18324
rect 31661 18320 32260 18322
rect 31661 18264 31666 18320
rect 31722 18264 32260 18320
rect 31661 18262 32260 18264
rect 31661 18259 31727 18262
rect 32254 18260 32260 18262
rect 32324 18260 32330 18324
rect 2681 18186 2747 18189
rect 7557 18186 7623 18189
rect 2681 18184 7623 18186
rect 2681 18128 2686 18184
rect 2742 18128 7562 18184
rect 7618 18128 7623 18184
rect 2681 18126 7623 18128
rect 2681 18123 2747 18126
rect 7557 18123 7623 18126
rect 8569 18186 8635 18189
rect 28165 18186 28231 18189
rect 32438 18186 32444 18188
rect 8569 18184 24042 18186
rect 8569 18128 8574 18184
rect 8630 18128 24042 18184
rect 8569 18126 24042 18128
rect 8569 18123 8635 18126
rect 3550 17988 3556 18052
rect 3620 18050 3626 18052
rect 3693 18050 3759 18053
rect 5349 18050 5415 18053
rect 5993 18050 6059 18053
rect 3620 18048 3986 18050
rect 3620 17992 3698 18048
rect 3754 17992 3986 18048
rect 3620 17990 3986 17992
rect 3620 17988 3626 17990
rect 3693 17987 3759 17990
rect 0 17914 800 17944
rect 2957 17914 3023 17917
rect 0 17912 3023 17914
rect 0 17856 2962 17912
rect 3018 17856 3023 17912
rect 0 17854 3023 17856
rect 0 17824 800 17854
rect 2957 17851 3023 17854
rect 3926 17778 3986 17990
rect 5349 18048 6059 18050
rect 5349 17992 5354 18048
rect 5410 17992 5998 18048
rect 6054 17992 6059 18048
rect 5349 17990 6059 17992
rect 5349 17987 5415 17990
rect 5993 17987 6059 17990
rect 12934 17988 12940 18052
rect 13004 18050 13010 18052
rect 13169 18050 13235 18053
rect 13004 18048 13235 18050
rect 13004 17992 13174 18048
rect 13230 17992 13235 18048
rect 13004 17990 13235 17992
rect 13004 17988 13010 17990
rect 13169 17987 13235 17990
rect 13353 18050 13419 18053
rect 16665 18050 16731 18053
rect 17493 18050 17559 18053
rect 18137 18052 18203 18053
rect 18086 18050 18092 18052
rect 13353 18048 17559 18050
rect 13353 17992 13358 18048
rect 13414 17992 16670 18048
rect 16726 17992 17498 18048
rect 17554 17992 17559 18048
rect 13353 17990 17559 17992
rect 18046 17990 18092 18050
rect 18156 18048 18203 18052
rect 18198 17992 18203 18048
rect 13353 17987 13419 17990
rect 16665 17987 16731 17990
rect 17493 17987 17559 17990
rect 18086 17988 18092 17990
rect 18156 17988 18203 17992
rect 18137 17987 18203 17988
rect 18321 18050 18387 18053
rect 20110 18050 20116 18052
rect 18321 18048 20116 18050
rect 18321 17992 18326 18048
rect 18382 17992 20116 18048
rect 18321 17990 20116 17992
rect 18321 17987 18387 17990
rect 20110 17988 20116 17990
rect 20180 17988 20186 18052
rect 20437 18050 20503 18053
rect 22686 18050 22692 18052
rect 20437 18048 22692 18050
rect 20437 17992 20442 18048
rect 20498 17992 22692 18048
rect 20437 17990 22692 17992
rect 20437 17987 20503 17990
rect 22686 17988 22692 17990
rect 22756 17988 22762 18052
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 7097 17914 7163 17917
rect 5398 17912 7163 17914
rect 5398 17856 7102 17912
rect 7158 17856 7163 17912
rect 5398 17854 7163 17856
rect 5398 17778 5458 17854
rect 7097 17851 7163 17854
rect 11329 17914 11395 17917
rect 17125 17916 17191 17917
rect 15510 17914 15516 17916
rect 11329 17912 15516 17914
rect 11329 17856 11334 17912
rect 11390 17856 15516 17912
rect 11329 17854 15516 17856
rect 11329 17851 11395 17854
rect 15510 17852 15516 17854
rect 15580 17852 15586 17916
rect 17125 17914 17172 17916
rect 17080 17912 17172 17914
rect 17080 17856 17130 17912
rect 17080 17854 17172 17856
rect 17125 17852 17172 17854
rect 17236 17852 17242 17916
rect 17902 17852 17908 17916
rect 17972 17914 17978 17916
rect 18137 17914 18203 17917
rect 20294 17914 20300 17916
rect 17972 17912 18203 17914
rect 17972 17856 18142 17912
rect 18198 17856 18203 17912
rect 17972 17854 18203 17856
rect 17972 17852 17978 17854
rect 17125 17851 17191 17852
rect 18137 17851 18203 17854
rect 18278 17854 20300 17914
rect 3926 17718 5458 17778
rect 5533 17778 5599 17781
rect 6729 17778 6795 17781
rect 5533 17776 6795 17778
rect 5533 17720 5538 17776
rect 5594 17720 6734 17776
rect 6790 17720 6795 17776
rect 5533 17718 6795 17720
rect 5533 17715 5599 17718
rect 6729 17715 6795 17718
rect 12433 17778 12499 17781
rect 18045 17778 18111 17781
rect 12433 17776 18111 17778
rect 12433 17720 12438 17776
rect 12494 17720 18050 17776
rect 18106 17720 18111 17776
rect 12433 17718 18111 17720
rect 12433 17715 12499 17718
rect 18045 17715 18111 17718
rect 8702 17580 8708 17644
rect 8772 17642 8778 17644
rect 10133 17642 10199 17645
rect 8772 17640 10199 17642
rect 8772 17584 10138 17640
rect 10194 17584 10199 17640
rect 8772 17582 10199 17584
rect 8772 17580 8778 17582
rect 10133 17579 10199 17582
rect 16021 17642 16087 17645
rect 17493 17642 17559 17645
rect 16021 17640 17559 17642
rect 16021 17584 16026 17640
rect 16082 17584 17498 17640
rect 17554 17584 17559 17640
rect 16021 17582 17559 17584
rect 16021 17579 16087 17582
rect 17493 17579 17559 17582
rect 17718 17580 17724 17644
rect 17788 17642 17794 17644
rect 18278 17642 18338 17854
rect 20294 17852 20300 17854
rect 20364 17852 20370 17916
rect 20437 17914 20503 17917
rect 20662 17914 20668 17916
rect 20437 17912 20668 17914
rect 20437 17856 20442 17912
rect 20498 17856 20668 17912
rect 20437 17854 20668 17856
rect 20437 17851 20503 17854
rect 20662 17852 20668 17854
rect 20732 17852 20738 17916
rect 20897 17914 20963 17917
rect 21030 17914 21036 17916
rect 20897 17912 21036 17914
rect 20897 17856 20902 17912
rect 20958 17856 21036 17912
rect 20897 17854 21036 17856
rect 20897 17851 20963 17854
rect 21030 17852 21036 17854
rect 21100 17852 21106 17916
rect 21725 17914 21791 17917
rect 22502 17914 22508 17916
rect 21725 17912 22508 17914
rect 21725 17856 21730 17912
rect 21786 17856 22508 17912
rect 21725 17854 22508 17856
rect 21725 17851 21791 17854
rect 22502 17852 22508 17854
rect 22572 17852 22578 17916
rect 23982 17914 24042 18126
rect 28165 18184 32444 18186
rect 28165 18128 28170 18184
rect 28226 18128 32444 18184
rect 28165 18126 32444 18128
rect 28165 18123 28231 18126
rect 32438 18124 32444 18126
rect 32508 18124 32514 18188
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 24301 17914 24367 17917
rect 23982 17912 24367 17914
rect 23982 17856 24306 17912
rect 24362 17856 24367 17912
rect 23982 17854 24367 17856
rect 24301 17851 24367 17854
rect 27654 17852 27660 17916
rect 27724 17914 27730 17916
rect 28257 17914 28323 17917
rect 27724 17912 28323 17914
rect 27724 17856 28262 17912
rect 28318 17856 28323 17912
rect 27724 17854 28323 17856
rect 27724 17852 27730 17854
rect 28257 17851 28323 17854
rect 18505 17778 18571 17781
rect 19701 17778 19767 17781
rect 18505 17776 19767 17778
rect 18505 17720 18510 17776
rect 18566 17720 19706 17776
rect 19762 17720 19767 17776
rect 18505 17718 19767 17720
rect 18505 17715 18571 17718
rect 19701 17715 19767 17718
rect 19977 17778 20043 17781
rect 23289 17778 23355 17781
rect 19977 17776 23355 17778
rect 19977 17720 19982 17776
rect 20038 17720 23294 17776
rect 23350 17720 23355 17776
rect 19977 17718 23355 17720
rect 19977 17715 20043 17718
rect 23289 17715 23355 17718
rect 18965 17644 19031 17645
rect 18965 17642 19012 17644
rect 17788 17582 18338 17642
rect 18920 17640 19012 17642
rect 18920 17584 18970 17640
rect 18920 17582 19012 17584
rect 17788 17580 17794 17582
rect 18965 17580 19012 17582
rect 19076 17580 19082 17644
rect 19609 17642 19675 17645
rect 19152 17640 19675 17642
rect 19152 17584 19614 17640
rect 19670 17584 19675 17640
rect 19152 17582 19675 17584
rect 18965 17579 19031 17580
rect 4981 17506 5047 17509
rect 14549 17506 14615 17509
rect 19152 17506 19212 17582
rect 19609 17579 19675 17582
rect 20662 17580 20668 17644
rect 20732 17642 20738 17644
rect 22461 17642 22527 17645
rect 20732 17640 22527 17642
rect 20732 17584 22466 17640
rect 22522 17584 22527 17640
rect 20732 17582 22527 17584
rect 20732 17580 20738 17582
rect 22461 17579 22527 17582
rect 4981 17504 12450 17506
rect 4981 17448 4986 17504
rect 5042 17448 12450 17504
rect 4981 17446 12450 17448
rect 4981 17443 5047 17446
rect 0 17370 800 17400
rect 4061 17370 4127 17373
rect 0 17368 4127 17370
rect 0 17312 4066 17368
rect 4122 17312 4127 17368
rect 0 17310 4127 17312
rect 0 17280 800 17310
rect 4061 17307 4127 17310
rect 7557 17370 7623 17373
rect 12390 17370 12450 17446
rect 14549 17504 19212 17506
rect 14549 17448 14554 17504
rect 14610 17448 19212 17504
rect 14549 17446 19212 17448
rect 19977 17506 20043 17509
rect 24761 17506 24827 17509
rect 19977 17504 24827 17506
rect 19977 17448 19982 17504
rect 20038 17448 24766 17504
rect 24822 17448 24827 17504
rect 19977 17446 24827 17448
rect 14549 17443 14615 17446
rect 19977 17443 20043 17446
rect 24761 17443 24827 17446
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 14273 17370 14339 17373
rect 7557 17368 11530 17370
rect 7557 17312 7562 17368
rect 7618 17312 11530 17368
rect 7557 17310 11530 17312
rect 12390 17368 14339 17370
rect 12390 17312 14278 17368
rect 14334 17312 14339 17368
rect 12390 17310 14339 17312
rect 7557 17307 7623 17310
rect 1669 17234 1735 17237
rect 3233 17234 3299 17237
rect 11470 17234 11530 17310
rect 14273 17307 14339 17310
rect 17401 17370 17467 17373
rect 18597 17370 18663 17373
rect 17401 17368 18663 17370
rect 17401 17312 17406 17368
rect 17462 17312 18602 17368
rect 18658 17312 18663 17368
rect 17401 17310 18663 17312
rect 17401 17307 17467 17310
rect 18597 17307 18663 17310
rect 18781 17370 18847 17373
rect 19190 17370 19196 17372
rect 18781 17368 19196 17370
rect 18781 17312 18786 17368
rect 18842 17312 19196 17368
rect 18781 17310 19196 17312
rect 18781 17307 18847 17310
rect 19190 17308 19196 17310
rect 19260 17308 19266 17372
rect 20805 17370 20871 17373
rect 27654 17370 27660 17372
rect 20805 17368 27660 17370
rect 20805 17312 20810 17368
rect 20866 17312 27660 17368
rect 20805 17310 27660 17312
rect 20805 17307 20871 17310
rect 27654 17308 27660 17310
rect 27724 17308 27730 17372
rect 16665 17234 16731 17237
rect 1669 17232 3299 17234
rect 1669 17176 1674 17232
rect 1730 17176 3238 17232
rect 3294 17176 3299 17232
rect 1669 17174 3299 17176
rect 1669 17171 1735 17174
rect 3233 17171 3299 17174
rect 3742 17174 11346 17234
rect 11470 17232 16731 17234
rect 11470 17176 16670 17232
rect 16726 17176 16731 17232
rect 11470 17174 16731 17176
rect 13 17098 79 17101
rect 1158 17098 1164 17100
rect 13 17096 1164 17098
rect 13 17040 18 17096
rect 74 17040 1164 17096
rect 13 17038 1164 17040
rect 13 17035 79 17038
rect 1158 17036 1164 17038
rect 1228 17036 1234 17100
rect 2129 17098 2195 17101
rect 3742 17098 3802 17174
rect 11145 17098 11211 17101
rect 2129 17096 3802 17098
rect 2129 17040 2134 17096
rect 2190 17040 3802 17096
rect 2129 17038 3802 17040
rect 3926 17096 11211 17098
rect 3926 17040 11150 17096
rect 11206 17040 11211 17096
rect 3926 17038 11211 17040
rect 11286 17098 11346 17174
rect 16665 17171 16731 17174
rect 16941 17234 17007 17237
rect 19701 17234 19767 17237
rect 16941 17232 19767 17234
rect 16941 17176 16946 17232
rect 17002 17176 19706 17232
rect 19762 17176 19767 17232
rect 16941 17174 19767 17176
rect 16941 17171 17007 17174
rect 19701 17171 19767 17174
rect 20253 17234 20319 17237
rect 23105 17234 23171 17237
rect 20253 17232 23171 17234
rect 20253 17176 20258 17232
rect 20314 17176 23110 17232
rect 23166 17176 23171 17232
rect 20253 17174 23171 17176
rect 20253 17171 20319 17174
rect 23105 17171 23171 17174
rect 27521 17234 27587 17237
rect 27981 17234 28047 17237
rect 27521 17232 28047 17234
rect 27521 17176 27526 17232
rect 27582 17176 27986 17232
rect 28042 17176 28047 17232
rect 27521 17174 28047 17176
rect 27521 17171 27587 17174
rect 27981 17171 28047 17174
rect 22461 17098 22527 17101
rect 11286 17096 22527 17098
rect 11286 17040 22466 17096
rect 22522 17040 22527 17096
rect 11286 17038 22527 17040
rect 1166 16962 1226 17036
rect 2129 17035 2195 17038
rect 3926 16962 3986 17038
rect 11145 17035 11211 17038
rect 22461 17035 22527 17038
rect 22921 17098 22987 17101
rect 28993 17098 29059 17101
rect 22921 17096 29059 17098
rect 22921 17040 22926 17096
rect 22982 17040 28998 17096
rect 29054 17040 29059 17096
rect 22921 17038 29059 17040
rect 22921 17035 22987 17038
rect 28993 17035 29059 17038
rect 1166 16902 3986 16962
rect 5533 16962 5599 16965
rect 8017 16962 8083 16965
rect 5533 16960 8083 16962
rect 5533 16904 5538 16960
rect 5594 16904 8022 16960
rect 8078 16904 8083 16960
rect 5533 16902 8083 16904
rect 5533 16899 5599 16902
rect 8017 16899 8083 16902
rect 12382 16900 12388 16964
rect 12452 16962 12458 16964
rect 18454 16962 18460 16964
rect 12452 16902 18460 16962
rect 12452 16900 12458 16902
rect 18454 16900 18460 16902
rect 18524 16900 18530 16964
rect 18597 16962 18663 16965
rect 24025 16962 24091 16965
rect 18597 16960 24091 16962
rect 18597 16904 18602 16960
rect 18658 16904 24030 16960
rect 24086 16904 24091 16960
rect 18597 16902 24091 16904
rect 18597 16899 18663 16902
rect 24025 16899 24091 16902
rect 4208 16896 4528 16897
rect 0 16826 800 16856
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 3509 16826 3575 16829
rect 0 16824 3575 16826
rect 0 16768 3514 16824
rect 3570 16768 3575 16824
rect 0 16766 3575 16768
rect 0 16736 800 16766
rect 3509 16763 3575 16766
rect 6269 16826 6335 16829
rect 10542 16826 10548 16828
rect 6269 16824 10548 16826
rect 6269 16768 6274 16824
rect 6330 16768 10548 16824
rect 6269 16766 10548 16768
rect 6269 16763 6335 16766
rect 10542 16764 10548 16766
rect 10612 16764 10618 16828
rect 10685 16826 10751 16829
rect 16389 16826 16455 16829
rect 10685 16824 16455 16826
rect 10685 16768 10690 16824
rect 10746 16768 16394 16824
rect 16450 16768 16455 16824
rect 10685 16766 16455 16768
rect 10685 16763 10751 16766
rect 16389 16763 16455 16766
rect 18413 16826 18479 16829
rect 19149 16826 19215 16829
rect 22093 16828 22159 16829
rect 18413 16824 19215 16826
rect 18413 16768 18418 16824
rect 18474 16768 19154 16824
rect 19210 16768 19215 16824
rect 18413 16766 19215 16768
rect 18413 16763 18479 16766
rect 19149 16763 19215 16766
rect 19374 16764 19380 16828
rect 19444 16826 19450 16828
rect 20294 16826 20300 16828
rect 19444 16766 20300 16826
rect 19444 16764 19450 16766
rect 20294 16764 20300 16766
rect 20364 16764 20370 16828
rect 22093 16824 22140 16828
rect 22204 16826 22210 16828
rect 22461 16826 22527 16829
rect 23289 16826 23355 16829
rect 27061 16826 27127 16829
rect 29453 16826 29519 16829
rect 22093 16768 22098 16824
rect 22093 16764 22140 16768
rect 22204 16766 22250 16826
rect 22461 16824 22754 16826
rect 22461 16768 22466 16824
rect 22522 16768 22754 16824
rect 22461 16766 22754 16768
rect 22204 16764 22210 16766
rect 22093 16763 22159 16764
rect 22461 16763 22527 16766
rect 3233 16690 3299 16693
rect 7373 16690 7439 16693
rect 7557 16692 7623 16693
rect 7557 16690 7604 16692
rect 3233 16688 7439 16690
rect 3233 16632 3238 16688
rect 3294 16632 7378 16688
rect 7434 16632 7439 16688
rect 3233 16630 7439 16632
rect 7512 16688 7604 16690
rect 7512 16632 7562 16688
rect 7512 16630 7604 16632
rect 3233 16627 3299 16630
rect 7373 16627 7439 16630
rect 7557 16628 7604 16630
rect 7668 16628 7674 16692
rect 10225 16690 10291 16693
rect 13169 16690 13235 16693
rect 10225 16688 13235 16690
rect 10225 16632 10230 16688
rect 10286 16632 13174 16688
rect 13230 16632 13235 16688
rect 10225 16630 13235 16632
rect 7557 16627 7623 16628
rect 10225 16627 10291 16630
rect 10872 16557 10932 16630
rect 13169 16627 13235 16630
rect 13670 16628 13676 16692
rect 13740 16690 13746 16692
rect 16021 16690 16087 16693
rect 13740 16688 16087 16690
rect 13740 16632 16026 16688
rect 16082 16632 16087 16688
rect 13740 16630 16087 16632
rect 13740 16628 13746 16630
rect 16021 16627 16087 16630
rect 16297 16690 16363 16693
rect 19057 16692 19123 16693
rect 19006 16690 19012 16692
rect 16297 16688 18752 16690
rect 16297 16632 16302 16688
rect 16358 16632 18752 16688
rect 16297 16630 18752 16632
rect 18966 16630 19012 16690
rect 19076 16688 19123 16692
rect 19118 16632 19123 16688
rect 16297 16627 16363 16630
rect 18692 16557 18752 16630
rect 19006 16628 19012 16630
rect 19076 16628 19123 16632
rect 19374 16628 19380 16692
rect 19444 16690 19450 16692
rect 19793 16690 19859 16693
rect 19444 16688 19859 16690
rect 19444 16632 19798 16688
rect 19854 16632 19859 16688
rect 19444 16630 19859 16632
rect 19444 16628 19450 16630
rect 19057 16627 19123 16628
rect 19793 16627 19859 16630
rect 20846 16628 20852 16692
rect 20916 16690 20922 16692
rect 21817 16690 21883 16693
rect 22001 16690 22067 16693
rect 22694 16690 22754 16766
rect 23289 16824 29519 16826
rect 23289 16768 23294 16824
rect 23350 16768 27066 16824
rect 27122 16768 29458 16824
rect 29514 16768 29519 16824
rect 23289 16766 29519 16768
rect 23289 16763 23355 16766
rect 27061 16763 27127 16766
rect 29453 16763 29519 16766
rect 29545 16690 29611 16693
rect 20916 16688 21883 16690
rect 20916 16632 21822 16688
rect 21878 16632 21883 16688
rect 20916 16630 21883 16632
rect 21966 16688 22570 16690
rect 21966 16632 22006 16688
rect 22062 16632 22570 16688
rect 21966 16630 22570 16632
rect 22694 16688 29611 16690
rect 22694 16632 29550 16688
rect 29606 16632 29611 16688
rect 22694 16630 29611 16632
rect 20916 16628 20922 16630
rect 21817 16627 21883 16630
rect 22001 16627 22067 16630
rect 22510 16557 22570 16630
rect 29545 16627 29611 16630
rect 2681 16554 2747 16557
rect 7189 16556 7255 16557
rect 5574 16554 5580 16556
rect 2681 16552 5580 16554
rect 2681 16496 2686 16552
rect 2742 16496 5580 16552
rect 2681 16494 5580 16496
rect 2681 16491 2747 16494
rect 5574 16492 5580 16494
rect 5644 16554 5650 16556
rect 6494 16554 6500 16556
rect 5644 16494 6500 16554
rect 5644 16492 5650 16494
rect 6494 16492 6500 16494
rect 6564 16492 6570 16556
rect 7189 16552 7236 16556
rect 7300 16554 7306 16556
rect 9029 16554 9095 16557
rect 9622 16554 9628 16556
rect 7189 16496 7194 16552
rect 7189 16492 7236 16496
rect 7300 16494 7346 16554
rect 9029 16552 9628 16554
rect 9029 16496 9034 16552
rect 9090 16496 9628 16552
rect 9029 16494 9628 16496
rect 7300 16492 7306 16494
rect 7189 16491 7255 16492
rect 9029 16491 9095 16494
rect 9622 16492 9628 16494
rect 9692 16492 9698 16556
rect 10869 16552 10935 16557
rect 10869 16496 10874 16552
rect 10930 16496 10935 16552
rect 10869 16491 10935 16496
rect 12801 16554 12867 16557
rect 16665 16554 16731 16557
rect 12801 16552 16731 16554
rect 12801 16496 12806 16552
rect 12862 16496 16670 16552
rect 16726 16496 16731 16552
rect 12801 16494 16731 16496
rect 12801 16491 12867 16494
rect 16665 16491 16731 16494
rect 18689 16552 18755 16557
rect 18689 16496 18694 16552
rect 18750 16496 18755 16552
rect 18689 16491 18755 16496
rect 18822 16492 18828 16556
rect 18892 16554 18898 16556
rect 21214 16554 21220 16556
rect 18892 16494 21220 16554
rect 18892 16492 18898 16494
rect 21214 16492 21220 16494
rect 21284 16492 21290 16556
rect 22461 16552 22570 16557
rect 22461 16496 22466 16552
rect 22522 16496 22570 16552
rect 22461 16494 22570 16496
rect 22461 16491 22527 16494
rect 2129 16418 2195 16421
rect 10910 16418 10916 16420
rect 2129 16416 10916 16418
rect 2129 16360 2134 16416
rect 2190 16360 10916 16416
rect 2129 16358 10916 16360
rect 2129 16355 2195 16358
rect 10910 16356 10916 16358
rect 10980 16356 10986 16420
rect 11329 16418 11395 16421
rect 13169 16418 13235 16421
rect 11329 16416 13235 16418
rect 11329 16360 11334 16416
rect 11390 16360 13174 16416
rect 13230 16360 13235 16416
rect 11329 16358 13235 16360
rect 11329 16355 11395 16358
rect 13169 16355 13235 16358
rect 14365 16418 14431 16421
rect 16389 16418 16455 16421
rect 14365 16416 16455 16418
rect 14365 16360 14370 16416
rect 14426 16360 16394 16416
rect 16450 16360 16455 16416
rect 14365 16358 16455 16360
rect 14365 16355 14431 16358
rect 16389 16355 16455 16358
rect 18229 16418 18295 16421
rect 19006 16418 19012 16420
rect 18229 16416 19012 16418
rect 18229 16360 18234 16416
rect 18290 16360 19012 16416
rect 18229 16358 19012 16360
rect 18229 16355 18295 16358
rect 19006 16356 19012 16358
rect 19076 16356 19082 16420
rect 20069 16418 20135 16421
rect 20529 16418 20595 16421
rect 20069 16416 20595 16418
rect 20069 16360 20074 16416
rect 20130 16360 20534 16416
rect 20590 16360 20595 16416
rect 20069 16358 20595 16360
rect 20069 16355 20135 16358
rect 20529 16355 20595 16358
rect 20846 16356 20852 16420
rect 20916 16418 20922 16420
rect 24577 16418 24643 16421
rect 20916 16416 24643 16418
rect 20916 16360 24582 16416
rect 24638 16360 24643 16416
rect 20916 16358 24643 16360
rect 20916 16356 20922 16358
rect 24577 16355 24643 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 1669 16284 1735 16285
rect 1669 16282 1716 16284
rect 1588 16280 1716 16282
rect 1780 16282 1786 16284
rect 11605 16282 11671 16285
rect 15469 16282 15535 16285
rect 16113 16282 16179 16285
rect 1780 16280 11671 16282
rect 1588 16224 1674 16280
rect 1780 16224 11610 16280
rect 11666 16224 11671 16280
rect 1588 16222 1716 16224
rect 1669 16220 1716 16222
rect 1780 16222 11671 16224
rect 1780 16220 1786 16222
rect 1669 16219 1735 16220
rect 11605 16219 11671 16222
rect 12390 16280 16179 16282
rect 12390 16224 15474 16280
rect 15530 16224 16118 16280
rect 16174 16224 16179 16280
rect 12390 16222 16179 16224
rect 0 16146 800 16176
rect 1301 16146 1367 16149
rect 12390 16146 12450 16222
rect 15469 16219 15535 16222
rect 16113 16219 16179 16222
rect 18086 16220 18092 16284
rect 18156 16282 18162 16284
rect 18229 16282 18295 16285
rect 18156 16280 18295 16282
rect 18156 16224 18234 16280
rect 18290 16224 18295 16280
rect 18156 16222 18295 16224
rect 18156 16220 18162 16222
rect 18229 16219 18295 16222
rect 18873 16280 18939 16285
rect 18873 16224 18878 16280
rect 18934 16224 18939 16280
rect 18873 16219 18939 16224
rect 19977 16282 20043 16285
rect 25313 16282 25379 16285
rect 19977 16280 25379 16282
rect 19977 16224 19982 16280
rect 20038 16224 25318 16280
rect 25374 16224 25379 16280
rect 19977 16222 25379 16224
rect 19977 16219 20043 16222
rect 25313 16219 25379 16222
rect 26325 16282 26391 16285
rect 31569 16282 31635 16285
rect 26325 16280 31635 16282
rect 26325 16224 26330 16280
rect 26386 16224 31574 16280
rect 31630 16224 31635 16280
rect 26325 16222 31635 16224
rect 26325 16219 26391 16222
rect 31569 16219 31635 16222
rect 0 16144 1367 16146
rect 0 16088 1306 16144
rect 1362 16088 1367 16144
rect 0 16086 1367 16088
rect 0 16056 800 16086
rect 1301 16083 1367 16086
rect 2730 16086 12450 16146
rect 15929 16146 15995 16149
rect 18876 16146 18936 16219
rect 24025 16146 24091 16149
rect 15929 16144 18936 16146
rect 15929 16088 15934 16144
rect 15990 16088 18936 16144
rect 15929 16086 18936 16088
rect 19014 16144 24091 16146
rect 19014 16088 24030 16144
rect 24086 16088 24091 16144
rect 19014 16086 24091 16088
rect 1577 16012 1643 16013
rect 1526 16010 1532 16012
rect 1450 15950 1532 16010
rect 1596 16010 1643 16012
rect 2730 16010 2790 16086
rect 15929 16083 15995 16086
rect 6729 16012 6795 16013
rect 1596 16008 2790 16010
rect 1638 15952 2790 16008
rect 1526 15948 1532 15950
rect 1596 15950 2790 15952
rect 1596 15948 1643 15950
rect 6678 15948 6684 16012
rect 6748 16010 6795 16012
rect 9121 16010 9187 16013
rect 18873 16010 18939 16013
rect 19014 16010 19074 16086
rect 24025 16083 24091 16086
rect 6748 16008 6840 16010
rect 6790 15952 6840 16008
rect 6748 15950 6840 15952
rect 9121 16008 19074 16010
rect 9121 15952 9126 16008
rect 9182 15952 18878 16008
rect 18934 15952 19074 16008
rect 9121 15950 19074 15952
rect 20529 16010 20595 16013
rect 23473 16010 23539 16013
rect 26325 16010 26391 16013
rect 20529 16008 26391 16010
rect 20529 15952 20534 16008
rect 20590 15952 23478 16008
rect 23534 15952 26330 16008
rect 26386 15952 26391 16008
rect 20529 15950 26391 15952
rect 6748 15948 6795 15950
rect 1577 15947 1643 15948
rect 6729 15947 6795 15948
rect 9121 15947 9187 15950
rect 18873 15947 18939 15950
rect 20529 15947 20595 15950
rect 23473 15947 23539 15950
rect 26325 15947 26391 15950
rect 15101 15874 15167 15877
rect 16062 15874 16068 15876
rect 15101 15872 16068 15874
rect 15101 15816 15106 15872
rect 15162 15816 16068 15872
rect 15101 15814 16068 15816
rect 15101 15811 15167 15814
rect 16062 15812 16068 15814
rect 16132 15812 16138 15876
rect 16481 15874 16547 15877
rect 19057 15874 19123 15877
rect 16481 15872 19123 15874
rect 16481 15816 16486 15872
rect 16542 15816 19062 15872
rect 19118 15816 19123 15872
rect 16481 15814 19123 15816
rect 16481 15811 16547 15814
rect 19057 15811 19123 15814
rect 19609 15874 19675 15877
rect 19977 15874 20043 15877
rect 26141 15874 26207 15877
rect 19609 15872 26207 15874
rect 19609 15816 19614 15872
rect 19670 15816 19982 15872
rect 20038 15816 26146 15872
rect 26202 15816 26207 15872
rect 19609 15814 26207 15816
rect 19609 15811 19675 15814
rect 19977 15811 20043 15814
rect 26141 15811 26207 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 8150 15676 8156 15740
rect 8220 15738 8226 15740
rect 9213 15738 9279 15741
rect 8220 15736 9279 15738
rect 8220 15680 9218 15736
rect 9274 15680 9279 15736
rect 8220 15678 9279 15680
rect 8220 15676 8226 15678
rect 9213 15675 9279 15678
rect 10869 15738 10935 15741
rect 14181 15738 14247 15741
rect 10869 15736 14247 15738
rect 10869 15680 10874 15736
rect 10930 15680 14186 15736
rect 14242 15680 14247 15736
rect 10869 15678 14247 15680
rect 10869 15675 10935 15678
rect 14181 15675 14247 15678
rect 14457 15738 14523 15741
rect 16205 15738 16271 15741
rect 17677 15738 17743 15741
rect 14457 15736 17743 15738
rect 14457 15680 14462 15736
rect 14518 15680 16210 15736
rect 16266 15680 17682 15736
rect 17738 15680 17743 15736
rect 14457 15678 17743 15680
rect 14457 15675 14523 15678
rect 16205 15675 16271 15678
rect 17677 15675 17743 15678
rect 18086 15676 18092 15740
rect 18156 15738 18162 15740
rect 20805 15738 20871 15741
rect 18156 15736 20871 15738
rect 18156 15680 20810 15736
rect 20866 15680 20871 15736
rect 18156 15678 20871 15680
rect 18156 15676 18162 15678
rect 20805 15675 20871 15678
rect 21633 15738 21699 15741
rect 24393 15738 24459 15741
rect 21633 15736 24459 15738
rect 21633 15680 21638 15736
rect 21694 15680 24398 15736
rect 24454 15680 24459 15736
rect 21633 15678 24459 15680
rect 21633 15675 21699 15678
rect 24393 15675 24459 15678
rect 26325 15738 26391 15741
rect 30414 15738 30420 15740
rect 26325 15736 30420 15738
rect 26325 15680 26330 15736
rect 26386 15680 30420 15736
rect 26325 15678 30420 15680
rect 26325 15675 26391 15678
rect 30414 15676 30420 15678
rect 30484 15676 30490 15740
rect 0 15602 800 15632
rect 3601 15602 3667 15605
rect 0 15600 3667 15602
rect 0 15544 3606 15600
rect 3662 15544 3667 15600
rect 0 15542 3667 15544
rect 0 15512 800 15542
rect 3601 15539 3667 15542
rect 4613 15602 4679 15605
rect 19241 15602 19307 15605
rect 4613 15600 19307 15602
rect 4613 15544 4618 15600
rect 4674 15544 19246 15600
rect 19302 15544 19307 15600
rect 4613 15542 19307 15544
rect 4613 15539 4679 15542
rect 19241 15539 19307 15542
rect 20069 15602 20135 15605
rect 20529 15602 20595 15605
rect 20069 15600 20595 15602
rect 20069 15544 20074 15600
rect 20130 15544 20534 15600
rect 20590 15544 20595 15600
rect 20069 15542 20595 15544
rect 20069 15539 20135 15542
rect 20529 15539 20595 15542
rect 20713 15602 20779 15605
rect 21541 15602 21607 15605
rect 24485 15602 24551 15605
rect 20713 15600 24551 15602
rect 20713 15544 20718 15600
rect 20774 15544 21546 15600
rect 21602 15544 24490 15600
rect 24546 15544 24551 15600
rect 20713 15542 24551 15544
rect 20713 15539 20779 15542
rect 21541 15539 21607 15542
rect 24485 15539 24551 15542
rect 2129 15466 2195 15469
rect 2262 15466 2268 15468
rect 2129 15464 2268 15466
rect 2129 15408 2134 15464
rect 2190 15408 2268 15464
rect 2129 15406 2268 15408
rect 2129 15403 2195 15406
rect 2262 15404 2268 15406
rect 2332 15404 2338 15468
rect 4705 15466 4771 15469
rect 20253 15466 20319 15469
rect 4705 15464 20319 15466
rect 4705 15408 4710 15464
rect 4766 15408 20258 15464
rect 20314 15408 20319 15464
rect 4705 15406 20319 15408
rect 4705 15403 4771 15406
rect 20253 15403 20319 15406
rect 21265 15466 21331 15469
rect 25313 15466 25379 15469
rect 21265 15464 25379 15466
rect 21265 15408 21270 15464
rect 21326 15408 25318 15464
rect 25374 15408 25379 15464
rect 21265 15406 25379 15408
rect 21265 15403 21331 15406
rect 25313 15403 25379 15406
rect 6453 15330 6519 15333
rect 8385 15330 8451 15333
rect 6453 15328 8451 15330
rect 6453 15272 6458 15328
rect 6514 15272 8390 15328
rect 8446 15272 8451 15328
rect 6453 15270 8451 15272
rect 6453 15267 6519 15270
rect 8385 15267 8451 15270
rect 13445 15330 13511 15333
rect 16798 15330 16804 15332
rect 13445 15328 16804 15330
rect 13445 15272 13450 15328
rect 13506 15272 16804 15328
rect 13445 15270 16804 15272
rect 13445 15267 13511 15270
rect 16798 15268 16804 15270
rect 16868 15268 16874 15332
rect 17401 15330 17467 15333
rect 19425 15330 19491 15333
rect 17401 15328 19491 15330
rect 17401 15272 17406 15328
rect 17462 15272 19430 15328
rect 19486 15272 19491 15328
rect 17401 15270 19491 15272
rect 17401 15267 17467 15270
rect 19425 15267 19491 15270
rect 20161 15330 20227 15333
rect 20294 15330 20300 15332
rect 20161 15328 20300 15330
rect 20161 15272 20166 15328
rect 20222 15272 20300 15328
rect 20161 15270 20300 15272
rect 20161 15267 20227 15270
rect 20294 15268 20300 15270
rect 20364 15268 20370 15332
rect 20989 15330 21055 15333
rect 22829 15330 22895 15333
rect 26049 15330 26115 15333
rect 20989 15328 22895 15330
rect 20989 15272 20994 15328
rect 21050 15272 22834 15328
rect 22890 15272 22895 15328
rect 20989 15270 22895 15272
rect 20989 15267 21055 15270
rect 22829 15267 22895 15270
rect 23062 15328 26115 15330
rect 23062 15272 26054 15328
rect 26110 15272 26115 15328
rect 23062 15270 26115 15272
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 5022 15132 5028 15196
rect 5092 15194 5098 15196
rect 9397 15194 9463 15197
rect 5092 15192 9463 15194
rect 5092 15136 9402 15192
rect 9458 15136 9463 15192
rect 5092 15134 9463 15136
rect 5092 15132 5098 15134
rect 9397 15131 9463 15134
rect 11697 15194 11763 15197
rect 17902 15194 17908 15196
rect 11697 15192 17908 15194
rect 11697 15136 11702 15192
rect 11758 15136 17908 15192
rect 11697 15134 17908 15136
rect 11697 15131 11763 15134
rect 17902 15132 17908 15134
rect 17972 15132 17978 15196
rect 18597 15194 18663 15197
rect 19190 15194 19196 15196
rect 18597 15192 19196 15194
rect 18597 15136 18602 15192
rect 18658 15136 19196 15192
rect 18597 15134 19196 15136
rect 18597 15131 18663 15134
rect 19190 15132 19196 15134
rect 19260 15132 19266 15196
rect 19977 15194 20043 15197
rect 20805 15196 20871 15197
rect 20805 15194 20852 15196
rect 19977 15192 20546 15194
rect 19977 15136 19982 15192
rect 20038 15136 20546 15192
rect 19977 15134 20546 15136
rect 20760 15192 20852 15194
rect 20760 15136 20810 15192
rect 20760 15134 20852 15136
rect 19977 15131 20043 15134
rect 0 15058 800 15088
rect 4061 15058 4127 15061
rect 0 15056 4127 15058
rect 0 15000 4066 15056
rect 4122 15000 4127 15056
rect 0 14998 4127 15000
rect 0 14968 800 14998
rect 4061 14995 4127 14998
rect 8201 15058 8267 15061
rect 20345 15058 20411 15061
rect 8201 15056 20411 15058
rect 8201 15000 8206 15056
rect 8262 15000 20350 15056
rect 20406 15000 20411 15056
rect 8201 14998 20411 15000
rect 20486 15058 20546 15134
rect 20805 15132 20852 15134
rect 20916 15132 20922 15196
rect 21582 15132 21588 15196
rect 21652 15194 21658 15196
rect 22001 15194 22067 15197
rect 21652 15192 22067 15194
rect 21652 15136 22006 15192
rect 22062 15136 22067 15192
rect 21652 15134 22067 15136
rect 21652 15132 21658 15134
rect 20805 15131 20871 15132
rect 22001 15131 22067 15134
rect 23062 15058 23122 15270
rect 26049 15267 26115 15270
rect 24209 15194 24275 15197
rect 24894 15194 24900 15196
rect 24209 15192 24900 15194
rect 24209 15136 24214 15192
rect 24270 15136 24900 15192
rect 24209 15134 24900 15136
rect 24209 15131 24275 15134
rect 24894 15132 24900 15134
rect 24964 15132 24970 15196
rect 25078 15132 25084 15196
rect 25148 15194 25154 15196
rect 25221 15194 25287 15197
rect 25148 15192 25287 15194
rect 25148 15136 25226 15192
rect 25282 15136 25287 15192
rect 25148 15134 25287 15136
rect 25148 15132 25154 15134
rect 25221 15131 25287 15134
rect 25497 15194 25563 15197
rect 27838 15194 27844 15196
rect 25497 15192 27844 15194
rect 25497 15136 25502 15192
rect 25558 15136 27844 15192
rect 25497 15134 27844 15136
rect 25497 15131 25563 15134
rect 27838 15132 27844 15134
rect 27908 15132 27914 15196
rect 20486 14998 23122 15058
rect 23289 15058 23355 15061
rect 27705 15058 27771 15061
rect 23289 15056 27771 15058
rect 23289 15000 23294 15056
rect 23350 15000 27710 15056
rect 27766 15000 27771 15056
rect 23289 14998 27771 15000
rect 8201 14995 8267 14998
rect 20345 14995 20411 14998
rect 23289 14995 23355 14998
rect 27705 14995 27771 14998
rect 1301 14922 1367 14925
rect 8109 14922 8175 14925
rect 1301 14920 8175 14922
rect 1301 14864 1306 14920
rect 1362 14864 8114 14920
rect 8170 14864 8175 14920
rect 1301 14862 8175 14864
rect 1301 14859 1367 14862
rect 8109 14859 8175 14862
rect 11605 14922 11671 14925
rect 16205 14922 16271 14925
rect 11605 14920 16271 14922
rect 11605 14864 11610 14920
rect 11666 14864 16210 14920
rect 16266 14864 16271 14920
rect 11605 14862 16271 14864
rect 11605 14859 11671 14862
rect 16205 14859 16271 14862
rect 18597 14922 18663 14925
rect 20989 14922 21055 14925
rect 24025 14924 24091 14925
rect 18597 14920 21055 14922
rect 18597 14864 18602 14920
rect 18658 14864 20994 14920
rect 21050 14864 21055 14920
rect 18597 14862 21055 14864
rect 18597 14859 18663 14862
rect 20989 14859 21055 14862
rect 23974 14860 23980 14924
rect 24044 14922 24091 14924
rect 24044 14920 24136 14922
rect 24086 14864 24136 14920
rect 24044 14862 24136 14864
rect 24044 14860 24091 14862
rect 30230 14860 30236 14924
rect 30300 14922 30306 14924
rect 42057 14922 42123 14925
rect 30300 14920 42123 14922
rect 30300 14864 42062 14920
rect 42118 14864 42123 14920
rect 30300 14862 42123 14864
rect 30300 14860 30306 14862
rect 24025 14859 24091 14860
rect 42057 14859 42123 14862
rect 16113 14786 16179 14789
rect 9630 14784 16179 14786
rect 9630 14728 16118 14784
rect 16174 14728 16179 14784
rect 9630 14726 16179 14728
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 9213 14650 9279 14653
rect 9630 14650 9690 14726
rect 16113 14723 16179 14726
rect 17166 14724 17172 14788
rect 17236 14786 17242 14788
rect 19374 14786 19380 14788
rect 17236 14726 19380 14786
rect 17236 14724 17242 14726
rect 19374 14724 19380 14726
rect 19444 14724 19450 14788
rect 19517 14786 19583 14789
rect 20294 14786 20300 14788
rect 19517 14784 20300 14786
rect 19517 14728 19522 14784
rect 19578 14728 20300 14784
rect 19517 14726 20300 14728
rect 19517 14723 19583 14726
rect 20294 14724 20300 14726
rect 20364 14786 20370 14788
rect 20529 14786 20595 14789
rect 21817 14786 21883 14789
rect 20364 14784 20595 14786
rect 20364 14728 20534 14784
rect 20590 14728 20595 14784
rect 20364 14726 20595 14728
rect 20364 14724 20370 14726
rect 20529 14723 20595 14726
rect 20670 14784 21883 14786
rect 20670 14728 21822 14784
rect 21878 14728 21883 14784
rect 20670 14726 21883 14728
rect 9213 14648 9690 14650
rect 9213 14592 9218 14648
rect 9274 14592 9690 14648
rect 9213 14590 9690 14592
rect 13169 14650 13235 14653
rect 13486 14650 13492 14652
rect 13169 14648 13492 14650
rect 13169 14592 13174 14648
rect 13230 14592 13492 14648
rect 13169 14590 13492 14592
rect 9213 14587 9279 14590
rect 13169 14587 13235 14590
rect 13486 14588 13492 14590
rect 13556 14588 13562 14652
rect 18454 14588 18460 14652
rect 18524 14650 18530 14652
rect 18689 14650 18755 14653
rect 18524 14648 18755 14650
rect 18524 14592 18694 14648
rect 18750 14592 18755 14648
rect 18524 14590 18755 14592
rect 18524 14588 18530 14590
rect 18689 14587 18755 14590
rect 19149 14650 19215 14653
rect 20670 14650 20730 14726
rect 21817 14723 21883 14726
rect 22737 14786 22803 14789
rect 26969 14786 27035 14789
rect 31109 14786 31175 14789
rect 22737 14784 31175 14786
rect 22737 14728 22742 14784
rect 22798 14728 26974 14784
rect 27030 14728 31114 14784
rect 31170 14728 31175 14784
rect 22737 14726 31175 14728
rect 22737 14723 22803 14726
rect 26969 14723 27035 14726
rect 31109 14723 31175 14726
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 19149 14648 20730 14650
rect 19149 14592 19154 14648
rect 19210 14592 20730 14648
rect 19149 14590 20730 14592
rect 20805 14650 20871 14653
rect 27429 14652 27495 14653
rect 27429 14650 27476 14652
rect 20805 14648 24916 14650
rect 20805 14592 20810 14648
rect 20866 14592 24916 14648
rect 20805 14590 24916 14592
rect 27384 14648 27476 14650
rect 27384 14592 27434 14648
rect 27384 14590 27476 14592
rect 19149 14587 19215 14590
rect 20805 14587 20871 14590
rect 1669 14514 1735 14517
rect 4337 14514 4403 14517
rect 5533 14514 5599 14517
rect 1669 14512 4124 14514
rect 1669 14456 1674 14512
rect 1730 14456 4124 14512
rect 1669 14454 4124 14456
rect 1669 14451 1735 14454
rect 0 14378 800 14408
rect 4064 14381 4124 14454
rect 4337 14512 5599 14514
rect 4337 14456 4342 14512
rect 4398 14456 5538 14512
rect 5594 14456 5599 14512
rect 4337 14454 5599 14456
rect 4337 14451 4403 14454
rect 5533 14451 5599 14454
rect 6453 14514 6519 14517
rect 7741 14514 7807 14517
rect 6453 14512 7807 14514
rect 6453 14456 6458 14512
rect 6514 14456 7746 14512
rect 7802 14456 7807 14512
rect 6453 14454 7807 14456
rect 6453 14451 6519 14454
rect 7741 14451 7807 14454
rect 10777 14514 10843 14517
rect 12617 14514 12683 14517
rect 13077 14516 13143 14517
rect 13077 14514 13124 14516
rect 10777 14512 12683 14514
rect 10777 14456 10782 14512
rect 10838 14456 12622 14512
rect 12678 14456 12683 14512
rect 10777 14454 12683 14456
rect 13032 14512 13124 14514
rect 13032 14456 13082 14512
rect 13032 14454 13124 14456
rect 10777 14451 10843 14454
rect 12617 14451 12683 14454
rect 13077 14452 13124 14454
rect 13188 14452 13194 14516
rect 13905 14514 13971 14517
rect 24669 14514 24735 14517
rect 13905 14512 24735 14514
rect 13905 14456 13910 14512
rect 13966 14456 24674 14512
rect 24730 14456 24735 14512
rect 13905 14454 24735 14456
rect 24856 14514 24916 14590
rect 27429 14588 27476 14590
rect 27540 14588 27546 14652
rect 27429 14587 27495 14588
rect 28625 14514 28691 14517
rect 24856 14512 28691 14514
rect 24856 14456 28630 14512
rect 28686 14456 28691 14512
rect 24856 14454 28691 14456
rect 13077 14451 13143 14452
rect 13905 14451 13971 14454
rect 24669 14451 24735 14454
rect 28625 14451 28691 14454
rect 1158 14378 1164 14380
rect 0 14318 1164 14378
rect 0 14288 800 14318
rect 1158 14316 1164 14318
rect 1228 14378 1234 14380
rect 3417 14378 3483 14381
rect 1228 14376 3483 14378
rect 1228 14320 3422 14376
rect 3478 14320 3483 14376
rect 1228 14318 3483 14320
rect 1228 14316 1234 14318
rect 3417 14315 3483 14318
rect 4061 14378 4127 14381
rect 5390 14378 5396 14380
rect 4061 14376 5396 14378
rect 4061 14320 4066 14376
rect 4122 14320 5396 14376
rect 4061 14318 5396 14320
rect 4061 14315 4127 14318
rect 5390 14316 5396 14318
rect 5460 14316 5466 14380
rect 6729 14378 6795 14381
rect 21265 14378 21331 14381
rect 6729 14376 21331 14378
rect 6729 14320 6734 14376
rect 6790 14320 21270 14376
rect 21326 14320 21331 14376
rect 6729 14318 21331 14320
rect 6729 14315 6795 14318
rect 21265 14315 21331 14318
rect 23197 14378 23263 14381
rect 27521 14378 27587 14381
rect 23197 14376 27587 14378
rect 23197 14320 23202 14376
rect 23258 14320 27526 14376
rect 27582 14320 27587 14376
rect 23197 14318 27587 14320
rect 23197 14315 23263 14318
rect 27521 14315 27587 14318
rect 28942 14316 28948 14380
rect 29012 14378 29018 14380
rect 35893 14378 35959 14381
rect 29012 14376 35959 14378
rect 29012 14320 35898 14376
rect 35954 14320 35959 14376
rect 29012 14318 35959 14320
rect 29012 14316 29018 14318
rect 35893 14315 35959 14318
rect 3877 14244 3943 14245
rect 3877 14240 3924 14244
rect 3988 14242 3994 14244
rect 5809 14242 5875 14245
rect 11513 14242 11579 14245
rect 3877 14184 3882 14240
rect 3877 14180 3924 14184
rect 3988 14182 4034 14242
rect 5809 14240 11579 14242
rect 5809 14184 5814 14240
rect 5870 14184 11518 14240
rect 11574 14184 11579 14240
rect 5809 14182 11579 14184
rect 3988 14180 3994 14182
rect 3877 14179 3943 14180
rect 5809 14179 5875 14182
rect 11513 14179 11579 14182
rect 13169 14242 13235 14245
rect 17861 14242 17927 14245
rect 13169 14240 17927 14242
rect 13169 14184 13174 14240
rect 13230 14184 17866 14240
rect 17922 14184 17927 14240
rect 13169 14182 17927 14184
rect 13169 14179 13235 14182
rect 17861 14179 17927 14182
rect 18045 14242 18111 14245
rect 19425 14242 19491 14245
rect 18045 14240 19491 14242
rect 18045 14184 18050 14240
rect 18106 14184 19430 14240
rect 19486 14184 19491 14240
rect 18045 14182 19491 14184
rect 18045 14179 18111 14182
rect 19425 14179 19491 14182
rect 20069 14242 20135 14245
rect 23565 14242 23631 14245
rect 20069 14240 23631 14242
rect 20069 14184 20074 14240
rect 20130 14184 23570 14240
rect 23626 14184 23631 14240
rect 20069 14182 23631 14184
rect 20069 14179 20135 14182
rect 23565 14179 23631 14182
rect 27429 14242 27495 14245
rect 28942 14242 28948 14244
rect 27429 14240 28948 14242
rect 27429 14184 27434 14240
rect 27490 14184 28948 14240
rect 27429 14182 28948 14184
rect 27429 14179 27495 14182
rect 28942 14180 28948 14182
rect 29012 14180 29018 14244
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 1025 14106 1091 14109
rect 11053 14106 11119 14109
rect 1025 14104 11119 14106
rect 1025 14048 1030 14104
rect 1086 14048 11058 14104
rect 11114 14048 11119 14104
rect 1025 14046 11119 14048
rect 1025 14043 1091 14046
rect 11053 14043 11119 14046
rect 12198 14044 12204 14108
rect 12268 14106 12274 14108
rect 14365 14106 14431 14109
rect 15745 14108 15811 14109
rect 12268 14104 14431 14106
rect 12268 14048 14370 14104
rect 14426 14048 14431 14104
rect 12268 14046 14431 14048
rect 12268 14044 12274 14046
rect 14365 14043 14431 14046
rect 15694 14044 15700 14108
rect 15764 14106 15811 14108
rect 15764 14104 15856 14106
rect 15806 14048 15856 14104
rect 15764 14046 15856 14048
rect 15764 14044 15811 14046
rect 16982 14044 16988 14108
rect 17052 14106 17058 14108
rect 18638 14106 18644 14108
rect 17052 14046 18644 14106
rect 17052 14044 17058 14046
rect 18638 14044 18644 14046
rect 18708 14106 18714 14108
rect 19149 14106 19215 14109
rect 20805 14106 20871 14109
rect 18708 14104 19215 14106
rect 18708 14048 19154 14104
rect 19210 14048 19215 14104
rect 18708 14046 19215 14048
rect 18708 14044 18714 14046
rect 15745 14043 15811 14044
rect 19149 14043 19215 14046
rect 19980 14104 20871 14106
rect 19980 14048 20810 14104
rect 20866 14048 20871 14104
rect 19980 14046 20871 14048
rect 19980 14004 20040 14046
rect 20805 14043 20871 14046
rect 21081 14106 21147 14109
rect 22737 14106 22803 14109
rect 23381 14108 23447 14109
rect 29269 14108 29335 14109
rect 23381 14106 23428 14108
rect 21081 14104 22803 14106
rect 21081 14048 21086 14104
rect 21142 14048 22742 14104
rect 22798 14048 22803 14104
rect 21081 14046 22803 14048
rect 23336 14104 23428 14106
rect 23336 14048 23386 14104
rect 23336 14046 23428 14048
rect 21081 14043 21147 14046
rect 22737 14043 22803 14046
rect 23381 14044 23428 14046
rect 23492 14044 23498 14108
rect 29269 14106 29316 14108
rect 29224 14104 29316 14106
rect 29224 14048 29274 14104
rect 29224 14046 29316 14048
rect 29269 14044 29316 14046
rect 29380 14044 29386 14108
rect 23381 14043 23447 14044
rect 29269 14043 29335 14044
rect 2313 13970 2379 13973
rect 2630 13970 2636 13972
rect 2313 13968 2636 13970
rect 2313 13912 2318 13968
rect 2374 13912 2636 13968
rect 2313 13910 2636 13912
rect 2313 13907 2379 13910
rect 2630 13908 2636 13910
rect 2700 13908 2706 13972
rect 2773 13970 2839 13973
rect 7230 13970 7236 13972
rect 2773 13968 7236 13970
rect 2773 13912 2778 13968
rect 2834 13912 7236 13968
rect 2773 13910 7236 13912
rect 2773 13907 2839 13910
rect 7230 13908 7236 13910
rect 7300 13970 7306 13972
rect 10777 13970 10843 13973
rect 7300 13968 10843 13970
rect 7300 13912 10782 13968
rect 10838 13912 10843 13968
rect 7300 13910 10843 13912
rect 7300 13908 7306 13910
rect 10777 13907 10843 13910
rect 10918 13910 13876 13970
rect 0 13834 800 13864
rect 2865 13834 2931 13837
rect 5257 13834 5323 13837
rect 0 13832 5323 13834
rect 0 13776 2870 13832
rect 2926 13776 5262 13832
rect 5318 13776 5323 13832
rect 0 13774 5323 13776
rect 0 13744 800 13774
rect 2865 13771 2931 13774
rect 5257 13771 5323 13774
rect 9857 13834 9923 13837
rect 10918 13834 10978 13910
rect 9857 13832 10978 13834
rect 9857 13776 9862 13832
rect 9918 13776 10978 13832
rect 9857 13774 10978 13776
rect 9857 13771 9923 13774
rect 12750 13772 12756 13836
rect 12820 13834 12826 13836
rect 13353 13834 13419 13837
rect 12820 13832 13419 13834
rect 12820 13776 13358 13832
rect 13414 13776 13419 13832
rect 12820 13774 13419 13776
rect 12820 13772 12826 13774
rect 13353 13771 13419 13774
rect 13537 13834 13603 13837
rect 13670 13834 13676 13836
rect 13537 13832 13676 13834
rect 13537 13776 13542 13832
rect 13598 13776 13676 13832
rect 13537 13774 13676 13776
rect 13537 13771 13603 13774
rect 13670 13772 13676 13774
rect 13740 13772 13746 13836
rect 13816 13834 13876 13910
rect 14222 13908 14228 13972
rect 14292 13970 14298 13972
rect 19704 13970 20040 14004
rect 14292 13944 20040 13970
rect 14292 13910 19764 13944
rect 14292 13908 14298 13910
rect 20846 13908 20852 13972
rect 20916 13970 20922 13972
rect 21449 13970 21515 13973
rect 20916 13968 21515 13970
rect 20916 13912 21454 13968
rect 21510 13912 21515 13968
rect 20916 13910 21515 13912
rect 20916 13908 20922 13910
rect 21449 13907 21515 13910
rect 23422 13908 23428 13972
rect 23492 13970 23498 13972
rect 23657 13970 23723 13973
rect 23492 13968 23723 13970
rect 23492 13912 23662 13968
rect 23718 13912 23723 13968
rect 23492 13910 23723 13912
rect 23492 13908 23498 13910
rect 23657 13907 23723 13910
rect 15285 13834 15351 13837
rect 13816 13832 15351 13834
rect 13816 13776 15290 13832
rect 15346 13776 15351 13832
rect 13816 13774 15351 13776
rect 15285 13771 15351 13774
rect 16389 13834 16455 13837
rect 19701 13834 19767 13837
rect 19977 13834 20043 13837
rect 16389 13832 20043 13834
rect 16389 13776 16394 13832
rect 16450 13776 19706 13832
rect 19762 13776 19982 13832
rect 20038 13776 20043 13832
rect 16389 13774 20043 13776
rect 16389 13771 16455 13774
rect 19701 13771 19767 13774
rect 19977 13771 20043 13774
rect 20161 13834 20227 13837
rect 29269 13834 29335 13837
rect 20161 13832 29335 13834
rect 20161 13776 20166 13832
rect 20222 13776 29274 13832
rect 29330 13776 29335 13832
rect 20161 13774 29335 13776
rect 20161 13771 20227 13774
rect 29269 13771 29335 13774
rect 1761 13698 1827 13701
rect 1894 13698 1900 13700
rect 1761 13696 1900 13698
rect 1761 13640 1766 13696
rect 1822 13640 1900 13696
rect 1761 13638 1900 13640
rect 1761 13635 1827 13638
rect 1894 13636 1900 13638
rect 1964 13636 1970 13700
rect 5533 13698 5599 13701
rect 5942 13698 5948 13700
rect 5533 13696 5948 13698
rect 5533 13640 5538 13696
rect 5594 13640 5948 13696
rect 5533 13638 5948 13640
rect 5533 13635 5599 13638
rect 5942 13636 5948 13638
rect 6012 13636 6018 13700
rect 6545 13698 6611 13701
rect 8334 13698 8340 13700
rect 6545 13696 8340 13698
rect 6545 13640 6550 13696
rect 6606 13640 8340 13696
rect 6545 13638 8340 13640
rect 6545 13635 6611 13638
rect 8334 13636 8340 13638
rect 8404 13636 8410 13700
rect 10317 13698 10383 13701
rect 12801 13698 12867 13701
rect 10317 13696 12867 13698
rect 10317 13640 10322 13696
rect 10378 13640 12806 13696
rect 12862 13640 12867 13696
rect 10317 13638 12867 13640
rect 10317 13635 10383 13638
rect 12801 13635 12867 13638
rect 12985 13698 13051 13701
rect 19517 13698 19583 13701
rect 12985 13696 19583 13698
rect 12985 13640 12990 13696
rect 13046 13640 19522 13696
rect 19578 13640 19583 13696
rect 12985 13638 19583 13640
rect 12985 13635 13051 13638
rect 19517 13635 19583 13638
rect 20805 13698 20871 13701
rect 28257 13698 28323 13701
rect 20805 13696 28323 13698
rect 20805 13640 20810 13696
rect 20866 13640 28262 13696
rect 28318 13640 28323 13696
rect 20805 13638 28323 13640
rect 20805 13635 20871 13638
rect 28257 13635 28323 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 5390 13500 5396 13564
rect 5460 13562 5466 13564
rect 8150 13562 8156 13564
rect 5460 13502 8156 13562
rect 5460 13500 5466 13502
rect 8150 13500 8156 13502
rect 8220 13500 8226 13564
rect 9438 13500 9444 13564
rect 9508 13562 9514 13564
rect 12249 13562 12315 13565
rect 9508 13560 12315 13562
rect 9508 13504 12254 13560
rect 12310 13504 12315 13560
rect 9508 13502 12315 13504
rect 9508 13500 9514 13502
rect 12249 13499 12315 13502
rect 14641 13562 14707 13565
rect 15837 13562 15903 13565
rect 19241 13562 19307 13565
rect 21817 13562 21883 13565
rect 14641 13560 21883 13562
rect 14641 13504 14646 13560
rect 14702 13504 15842 13560
rect 15898 13504 19246 13560
rect 19302 13504 21822 13560
rect 21878 13504 21883 13560
rect 14641 13502 21883 13504
rect 14641 13499 14707 13502
rect 15837 13499 15903 13502
rect 19241 13499 19307 13502
rect 21817 13499 21883 13502
rect 22093 13564 22159 13565
rect 22093 13560 22140 13564
rect 22204 13562 22210 13564
rect 22645 13562 22711 13565
rect 30373 13562 30439 13565
rect 22093 13504 22098 13560
rect 22093 13500 22140 13504
rect 22204 13502 22250 13562
rect 22645 13560 30439 13562
rect 22645 13504 22650 13560
rect 22706 13504 30378 13560
rect 30434 13504 30439 13560
rect 22645 13502 30439 13504
rect 22204 13500 22210 13502
rect 22093 13499 22159 13500
rect 22645 13499 22711 13502
rect 30373 13499 30439 13502
rect 3877 13426 3943 13429
rect 7414 13426 7420 13428
rect 3877 13424 7420 13426
rect 3877 13368 3882 13424
rect 3938 13368 7420 13424
rect 3877 13366 7420 13368
rect 3877 13363 3943 13366
rect 7414 13364 7420 13366
rect 7484 13364 7490 13428
rect 9673 13426 9739 13429
rect 18137 13426 18203 13429
rect 21725 13426 21791 13429
rect 22553 13428 22619 13429
rect 9673 13424 21791 13426
rect 9673 13368 9678 13424
rect 9734 13368 18142 13424
rect 18198 13368 21730 13424
rect 21786 13368 21791 13424
rect 9673 13366 21791 13368
rect 9673 13363 9739 13366
rect 18137 13363 18203 13366
rect 21725 13363 21791 13366
rect 22502 13364 22508 13428
rect 22572 13426 22619 13428
rect 22737 13426 22803 13429
rect 23657 13426 23723 13429
rect 22572 13424 22664 13426
rect 22614 13368 22664 13424
rect 22572 13366 22664 13368
rect 22737 13424 23723 13426
rect 22737 13368 22742 13424
rect 22798 13368 23662 13424
rect 23718 13368 23723 13424
rect 22737 13366 23723 13368
rect 22572 13364 22619 13366
rect 22553 13363 22619 13364
rect 22737 13363 22803 13366
rect 23657 13363 23723 13366
rect 23841 13426 23907 13429
rect 30465 13426 30531 13429
rect 23841 13424 30531 13426
rect 23841 13368 23846 13424
rect 23902 13368 30470 13424
rect 30526 13368 30531 13424
rect 23841 13366 30531 13368
rect 23841 13363 23907 13366
rect 30465 13363 30531 13366
rect 0 13290 800 13320
rect 2998 13290 3004 13292
rect 0 13230 3004 13290
rect 0 13200 800 13230
rect 2998 13228 3004 13230
rect 3068 13228 3074 13292
rect 3877 13290 3943 13293
rect 5206 13290 5212 13292
rect 3877 13288 5212 13290
rect 3877 13232 3882 13288
rect 3938 13232 5212 13288
rect 3877 13230 5212 13232
rect 3877 13227 3943 13230
rect 5206 13228 5212 13230
rect 5276 13228 5282 13292
rect 7598 13228 7604 13292
rect 7668 13290 7674 13292
rect 15193 13290 15259 13293
rect 7668 13288 15259 13290
rect 7668 13232 15198 13288
rect 15254 13232 15259 13288
rect 7668 13230 15259 13232
rect 7668 13228 7674 13230
rect 15193 13227 15259 13230
rect 15745 13290 15811 13293
rect 18454 13290 18460 13292
rect 15745 13288 18460 13290
rect 15745 13232 15750 13288
rect 15806 13232 18460 13288
rect 15745 13230 18460 13232
rect 15745 13227 15811 13230
rect 18454 13228 18460 13230
rect 18524 13228 18530 13292
rect 18597 13290 18663 13293
rect 21449 13290 21515 13293
rect 23565 13290 23631 13293
rect 25313 13290 25379 13293
rect 18597 13288 25379 13290
rect 18597 13232 18602 13288
rect 18658 13232 21454 13288
rect 21510 13232 23570 13288
rect 23626 13232 25318 13288
rect 25374 13232 25379 13288
rect 18597 13230 25379 13232
rect 18597 13227 18663 13230
rect 21449 13227 21515 13230
rect 23565 13227 23631 13230
rect 25313 13227 25379 13230
rect 26049 13290 26115 13293
rect 27889 13290 27955 13293
rect 26049 13288 27955 13290
rect 26049 13232 26054 13288
rect 26110 13232 27894 13288
rect 27950 13232 27955 13288
rect 26049 13230 27955 13232
rect 26049 13227 26115 13230
rect 27889 13227 27955 13230
rect 3509 13156 3575 13157
rect 3509 13152 3556 13156
rect 3620 13154 3626 13156
rect 4153 13154 4219 13157
rect 9254 13154 9260 13156
rect 3509 13096 3514 13152
rect 3509 13092 3556 13096
rect 3620 13094 3666 13154
rect 4153 13152 9260 13154
rect 4153 13096 4158 13152
rect 4214 13096 9260 13152
rect 4153 13094 9260 13096
rect 3620 13092 3626 13094
rect 3509 13091 3575 13092
rect 4153 13091 4219 13094
rect 9254 13092 9260 13094
rect 9324 13092 9330 13156
rect 10358 13092 10364 13156
rect 10428 13154 10434 13156
rect 12341 13154 12407 13157
rect 10428 13152 12407 13154
rect 10428 13096 12346 13152
rect 12402 13096 12407 13152
rect 10428 13094 12407 13096
rect 10428 13092 10434 13094
rect 12341 13091 12407 13094
rect 12801 13154 12867 13157
rect 18454 13154 18460 13156
rect 12801 13152 18460 13154
rect 12801 13096 12806 13152
rect 12862 13096 18460 13152
rect 12801 13094 18460 13096
rect 12801 13091 12867 13094
rect 18454 13092 18460 13094
rect 18524 13092 18530 13156
rect 18873 13154 18939 13157
rect 19374 13154 19380 13156
rect 18873 13152 19380 13154
rect 18873 13096 18878 13152
rect 18934 13096 19380 13152
rect 18873 13094 19380 13096
rect 18873 13091 18939 13094
rect 19374 13092 19380 13094
rect 19444 13092 19450 13156
rect 21909 13154 21975 13157
rect 25957 13154 26023 13157
rect 21909 13152 26023 13154
rect 21909 13096 21914 13152
rect 21970 13096 25962 13152
rect 26018 13096 26023 13152
rect 21909 13094 26023 13096
rect 21909 13091 21975 13094
rect 25957 13091 26023 13094
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 3509 13018 3575 13021
rect 7925 13018 7991 13021
rect 10593 13020 10659 13021
rect 3509 13016 7991 13018
rect 3509 12960 3514 13016
rect 3570 12960 7930 13016
rect 7986 12960 7991 13016
rect 3509 12958 7991 12960
rect 3509 12955 3575 12958
rect 7925 12955 7991 12958
rect 10542 12956 10548 13020
rect 10612 13018 10659 13020
rect 12893 13018 12959 13021
rect 21817 13018 21883 13021
rect 23565 13018 23631 13021
rect 10612 13016 10704 13018
rect 10654 12960 10704 13016
rect 10612 12958 10704 12960
rect 12893 13016 19488 13018
rect 12893 12960 12898 13016
rect 12954 12960 19488 13016
rect 12893 12958 19488 12960
rect 10612 12956 10659 12958
rect 10593 12955 10659 12956
rect 12893 12955 12959 12958
rect 5901 12882 5967 12885
rect 4846 12880 5967 12882
rect 4846 12824 5906 12880
rect 5962 12824 5967 12880
rect 4846 12822 5967 12824
rect 1669 12746 1735 12749
rect 3509 12746 3575 12749
rect 4846 12746 4906 12822
rect 5901 12819 5967 12822
rect 7373 12882 7439 12885
rect 10869 12882 10935 12885
rect 15285 12882 15351 12885
rect 7373 12880 10935 12882
rect 7373 12824 7378 12880
rect 7434 12824 10874 12880
rect 10930 12824 10935 12880
rect 7373 12822 10935 12824
rect 7373 12819 7439 12822
rect 10869 12819 10935 12822
rect 11102 12880 15351 12882
rect 11102 12824 15290 12880
rect 15346 12824 15351 12880
rect 11102 12822 15351 12824
rect 11102 12746 11162 12822
rect 15285 12819 15351 12822
rect 16798 12820 16804 12884
rect 16868 12882 16874 12884
rect 17493 12882 17559 12885
rect 18086 12882 18092 12884
rect 16868 12880 18092 12882
rect 16868 12824 17498 12880
rect 17554 12824 18092 12880
rect 16868 12822 18092 12824
rect 16868 12820 16874 12822
rect 17493 12819 17559 12822
rect 18086 12820 18092 12822
rect 18156 12820 18162 12884
rect 19428 12882 19488 12958
rect 21817 13016 23631 13018
rect 21817 12960 21822 13016
rect 21878 12960 23570 13016
rect 23626 12960 23631 13016
rect 21817 12958 23631 12960
rect 21817 12955 21883 12958
rect 23565 12955 23631 12958
rect 23749 13018 23815 13021
rect 29729 13018 29795 13021
rect 23749 13016 29795 13018
rect 23749 12960 23754 13016
rect 23810 12960 29734 13016
rect 29790 12960 29795 13016
rect 23749 12958 29795 12960
rect 23749 12955 23815 12958
rect 29729 12955 29795 12958
rect 19701 12882 19767 12885
rect 19428 12880 19767 12882
rect 19428 12824 19706 12880
rect 19762 12824 19767 12880
rect 19428 12822 19767 12824
rect 19701 12819 19767 12822
rect 25865 12882 25931 12885
rect 28257 12882 28323 12885
rect 25865 12880 28323 12882
rect 25865 12824 25870 12880
rect 25926 12824 28262 12880
rect 28318 12824 28323 12880
rect 25865 12822 28323 12824
rect 25865 12819 25931 12822
rect 28257 12819 28323 12822
rect 17217 12746 17283 12749
rect 21725 12746 21791 12749
rect 1669 12744 4906 12746
rect 1669 12688 1674 12744
rect 1730 12688 3514 12744
rect 3570 12688 4906 12744
rect 1669 12686 4906 12688
rect 4984 12686 11162 12746
rect 12390 12744 21791 12746
rect 12390 12688 17222 12744
rect 17278 12688 21730 12744
rect 21786 12688 21791 12744
rect 12390 12686 21791 12688
rect 1669 12683 1735 12686
rect 3509 12683 3575 12686
rect 0 12610 800 12640
rect 3785 12610 3851 12613
rect 0 12608 3851 12610
rect 0 12552 3790 12608
rect 3846 12552 3851 12608
rect 0 12550 3851 12552
rect 0 12520 800 12550
rect 3785 12547 3851 12550
rect 4654 12548 4660 12612
rect 4724 12610 4730 12612
rect 4984 12610 5044 12686
rect 4724 12550 5044 12610
rect 4724 12548 4730 12550
rect 5574 12548 5580 12612
rect 5644 12610 5650 12612
rect 8937 12610 9003 12613
rect 12390 12610 12450 12686
rect 17217 12683 17283 12686
rect 21725 12683 21791 12686
rect 23473 12746 23539 12749
rect 32305 12746 32371 12749
rect 23473 12744 32371 12746
rect 23473 12688 23478 12744
rect 23534 12688 32310 12744
rect 32366 12688 32371 12744
rect 23473 12686 32371 12688
rect 23473 12683 23539 12686
rect 32305 12683 32371 12686
rect 5644 12608 12450 12610
rect 5644 12552 8942 12608
rect 8998 12552 12450 12608
rect 5644 12550 12450 12552
rect 5644 12548 5650 12550
rect 8937 12547 9003 12550
rect 13854 12548 13860 12612
rect 13924 12610 13930 12612
rect 14089 12610 14155 12613
rect 13924 12608 14155 12610
rect 13924 12552 14094 12608
rect 14150 12552 14155 12608
rect 13924 12550 14155 12552
rect 13924 12548 13930 12550
rect 14089 12547 14155 12550
rect 16205 12610 16271 12613
rect 17861 12610 17927 12613
rect 16205 12608 17927 12610
rect 16205 12552 16210 12608
rect 16266 12552 17866 12608
rect 17922 12552 17927 12608
rect 16205 12550 17927 12552
rect 16205 12547 16271 12550
rect 17861 12547 17927 12550
rect 18413 12610 18479 12613
rect 19609 12610 19675 12613
rect 18413 12608 19675 12610
rect 18413 12552 18418 12608
rect 18474 12552 19614 12608
rect 19670 12552 19675 12608
rect 18413 12550 19675 12552
rect 18413 12547 18479 12550
rect 19609 12547 19675 12550
rect 21173 12610 21239 12613
rect 22318 12610 22324 12612
rect 21173 12608 22324 12610
rect 21173 12552 21178 12608
rect 21234 12552 22324 12608
rect 21173 12550 22324 12552
rect 21173 12547 21239 12550
rect 22318 12548 22324 12550
rect 22388 12548 22394 12612
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 4981 12474 5047 12477
rect 5390 12474 5396 12476
rect 4981 12472 5396 12474
rect 4981 12416 4986 12472
rect 5042 12416 5396 12472
rect 4981 12414 5396 12416
rect 4981 12411 5047 12414
rect 5390 12412 5396 12414
rect 5460 12412 5466 12476
rect 6678 12412 6684 12476
rect 6748 12474 6754 12476
rect 8569 12474 8635 12477
rect 6748 12472 8635 12474
rect 6748 12416 8574 12472
rect 8630 12416 8635 12472
rect 6748 12414 8635 12416
rect 6748 12412 6754 12414
rect 8569 12411 8635 12414
rect 9857 12474 9923 12477
rect 11421 12474 11487 12477
rect 9857 12472 11487 12474
rect 9857 12416 9862 12472
rect 9918 12416 11426 12472
rect 11482 12416 11487 12472
rect 9857 12414 11487 12416
rect 9857 12411 9923 12414
rect 11421 12411 11487 12414
rect 12985 12474 13051 12477
rect 15009 12474 15075 12477
rect 18045 12474 18111 12477
rect 12985 12472 15075 12474
rect 12985 12416 12990 12472
rect 13046 12416 15014 12472
rect 15070 12416 15075 12472
rect 12985 12414 15075 12416
rect 12985 12411 13051 12414
rect 15009 12411 15075 12414
rect 16530 12472 18111 12474
rect 16530 12416 18050 12472
rect 18106 12416 18111 12472
rect 16530 12414 18111 12416
rect 1853 12338 1919 12341
rect 8753 12338 8819 12341
rect 1853 12336 8819 12338
rect 1853 12280 1858 12336
rect 1914 12280 8758 12336
rect 8814 12280 8819 12336
rect 1853 12278 8819 12280
rect 1853 12275 1919 12278
rect 8753 12275 8819 12278
rect 10501 12338 10567 12341
rect 16530 12338 16590 12414
rect 18045 12411 18111 12414
rect 18321 12474 18387 12477
rect 18638 12474 18644 12476
rect 18321 12472 18644 12474
rect 18321 12416 18326 12472
rect 18382 12416 18644 12472
rect 18321 12414 18644 12416
rect 18321 12411 18387 12414
rect 18638 12412 18644 12414
rect 18708 12412 18714 12476
rect 20621 12474 20687 12477
rect 25681 12474 25747 12477
rect 28165 12474 28231 12477
rect 31661 12476 31727 12477
rect 31661 12474 31708 12476
rect 20621 12472 28231 12474
rect 20621 12416 20626 12472
rect 20682 12416 25686 12472
rect 25742 12416 28170 12472
rect 28226 12416 28231 12472
rect 20621 12414 28231 12416
rect 31616 12472 31708 12474
rect 31616 12416 31666 12472
rect 31616 12414 31708 12416
rect 20621 12411 20687 12414
rect 25681 12411 25747 12414
rect 28165 12411 28231 12414
rect 31661 12412 31708 12414
rect 31772 12412 31778 12476
rect 31661 12411 31727 12412
rect 10501 12336 16590 12338
rect 10501 12280 10506 12336
rect 10562 12280 16590 12336
rect 10501 12278 16590 12280
rect 10501 12275 10567 12278
rect 16982 12276 16988 12340
rect 17052 12338 17058 12340
rect 17309 12338 17375 12341
rect 17052 12336 17375 12338
rect 17052 12280 17314 12336
rect 17370 12280 17375 12336
rect 17052 12278 17375 12280
rect 17052 12276 17058 12278
rect 17309 12275 17375 12278
rect 17585 12338 17651 12341
rect 17902 12338 17908 12340
rect 17585 12336 17908 12338
rect 17585 12280 17590 12336
rect 17646 12280 17908 12336
rect 17585 12278 17908 12280
rect 17585 12275 17651 12278
rect 17902 12276 17908 12278
rect 17972 12276 17978 12340
rect 19701 12338 19767 12341
rect 20662 12338 20668 12340
rect 19701 12336 20668 12338
rect 19701 12280 19706 12336
rect 19762 12280 20668 12336
rect 19701 12278 20668 12280
rect 19701 12275 19767 12278
rect 20662 12276 20668 12278
rect 20732 12276 20738 12340
rect 26233 12338 26299 12341
rect 22050 12336 26299 12338
rect 22050 12280 26238 12336
rect 26294 12280 26299 12336
rect 22050 12278 26299 12280
rect 4521 12202 4587 12205
rect 6269 12202 6335 12205
rect 4521 12200 6335 12202
rect 4521 12144 4526 12200
rect 4582 12144 6274 12200
rect 6330 12144 6335 12200
rect 4521 12142 6335 12144
rect 4521 12139 4587 12142
rect 6269 12139 6335 12142
rect 7189 12202 7255 12205
rect 16941 12202 17007 12205
rect 7189 12200 17007 12202
rect 7189 12144 7194 12200
rect 7250 12144 16946 12200
rect 17002 12144 17007 12200
rect 7189 12142 17007 12144
rect 7189 12139 7255 12142
rect 16941 12139 17007 12142
rect 17534 12140 17540 12204
rect 17604 12202 17610 12204
rect 20478 12202 20484 12204
rect 17604 12142 20484 12202
rect 17604 12140 17610 12142
rect 20478 12140 20484 12142
rect 20548 12140 20554 12204
rect 20621 12202 20687 12205
rect 20989 12202 21055 12205
rect 20621 12200 21055 12202
rect 20621 12144 20626 12200
rect 20682 12144 20994 12200
rect 21050 12144 21055 12200
rect 20621 12142 21055 12144
rect 20621 12139 20687 12142
rect 20989 12139 21055 12142
rect 21817 12202 21883 12205
rect 22050 12202 22110 12278
rect 26233 12275 26299 12278
rect 27654 12276 27660 12340
rect 27724 12338 27730 12340
rect 29545 12338 29611 12341
rect 31661 12340 31727 12341
rect 31661 12338 31708 12340
rect 27724 12336 29611 12338
rect 27724 12280 29550 12336
rect 29606 12280 29611 12336
rect 27724 12278 29611 12280
rect 31616 12336 31708 12338
rect 31616 12280 31666 12336
rect 31616 12278 31708 12280
rect 27724 12276 27730 12278
rect 29545 12275 29611 12278
rect 31661 12276 31708 12278
rect 31772 12276 31778 12340
rect 31661 12275 31727 12276
rect 21817 12200 22110 12202
rect 21817 12144 21822 12200
rect 21878 12144 22110 12200
rect 21817 12142 22110 12144
rect 21817 12139 21883 12142
rect 0 12066 800 12096
rect 1342 12066 1348 12068
rect 0 12006 1348 12066
rect 0 11976 800 12006
rect 1342 12004 1348 12006
rect 1412 12066 1418 12068
rect 3141 12066 3207 12069
rect 6545 12066 6611 12069
rect 1412 12064 3207 12066
rect 1412 12008 3146 12064
rect 3202 12008 3207 12064
rect 1412 12006 3207 12008
rect 1412 12004 1418 12006
rect 3141 12003 3207 12006
rect 3328 12064 6611 12066
rect 3328 12008 6550 12064
rect 6606 12008 6611 12064
rect 3328 12006 6611 12008
rect 2405 11930 2471 11933
rect 3328 11930 3388 12006
rect 6545 12003 6611 12006
rect 10542 12004 10548 12068
rect 10612 12066 10618 12068
rect 17493 12066 17559 12069
rect 18597 12068 18663 12069
rect 18597 12066 18644 12068
rect 10612 12064 17559 12066
rect 10612 12008 17498 12064
rect 17554 12008 17559 12064
rect 10612 12006 17559 12008
rect 18552 12064 18644 12066
rect 18552 12008 18602 12064
rect 18552 12006 18644 12008
rect 10612 12004 10618 12006
rect 17493 12003 17559 12006
rect 18597 12004 18644 12006
rect 18708 12004 18714 12068
rect 19425 12064 19491 12069
rect 19425 12008 19430 12064
rect 19486 12008 19491 12064
rect 18597 12003 18663 12004
rect 19425 12003 19491 12008
rect 20662 12004 20668 12068
rect 20732 12066 20738 12068
rect 20805 12066 20871 12069
rect 20732 12064 20871 12066
rect 20732 12008 20810 12064
rect 20866 12008 20871 12064
rect 20732 12006 20871 12008
rect 20732 12004 20738 12006
rect 20805 12003 20871 12006
rect 21030 12004 21036 12068
rect 21100 12066 21106 12068
rect 21173 12066 21239 12069
rect 21100 12064 21239 12066
rect 21100 12008 21178 12064
rect 21234 12008 21239 12064
rect 21100 12006 21239 12008
rect 21100 12004 21106 12006
rect 21173 12003 21239 12006
rect 21449 12066 21515 12069
rect 27429 12066 27495 12069
rect 34789 12066 34855 12069
rect 21449 12064 26986 12066
rect 21449 12008 21454 12064
rect 21510 12008 26986 12064
rect 21449 12006 26986 12008
rect 21449 12003 21515 12006
rect 2405 11928 3388 11930
rect 2405 11872 2410 11928
rect 2466 11872 3388 11928
rect 2405 11870 3388 11872
rect 2405 11867 2471 11870
rect 5574 11868 5580 11932
rect 5644 11930 5650 11932
rect 5717 11930 5783 11933
rect 5644 11928 5783 11930
rect 5644 11872 5722 11928
rect 5778 11872 5783 11928
rect 5644 11870 5783 11872
rect 5644 11868 5650 11870
rect 5717 11867 5783 11870
rect 7782 11868 7788 11932
rect 7852 11930 7858 11932
rect 11329 11930 11395 11933
rect 7852 11928 11395 11930
rect 7852 11872 11334 11928
rect 11390 11872 11395 11928
rect 7852 11870 11395 11872
rect 7852 11868 7858 11870
rect 11329 11867 11395 11870
rect 13353 11930 13419 11933
rect 18321 11930 18387 11933
rect 13353 11928 18387 11930
rect 13353 11872 13358 11928
rect 13414 11872 18326 11928
rect 18382 11872 18387 11928
rect 13353 11870 18387 11872
rect 13353 11867 13419 11870
rect 18321 11867 18387 11870
rect 18597 11930 18663 11933
rect 19006 11930 19012 11932
rect 18597 11928 19012 11930
rect 18597 11872 18602 11928
rect 18658 11872 19012 11928
rect 18597 11870 19012 11872
rect 18597 11867 18663 11870
rect 19006 11868 19012 11870
rect 19076 11868 19082 11932
rect 19428 11797 19488 12003
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 20478 11868 20484 11932
rect 20548 11930 20554 11932
rect 25221 11930 25287 11933
rect 20548 11928 25287 11930
rect 20548 11872 25226 11928
rect 25282 11872 25287 11928
rect 20548 11870 25287 11872
rect 26926 11930 26986 12006
rect 27429 12064 34855 12066
rect 27429 12008 27434 12064
rect 27490 12008 34794 12064
rect 34850 12008 34855 12064
rect 27429 12006 34855 12008
rect 27429 12003 27495 12006
rect 34789 12003 34855 12006
rect 33225 11930 33291 11933
rect 26926 11928 33291 11930
rect 26926 11872 33230 11928
rect 33286 11872 33291 11928
rect 26926 11870 33291 11872
rect 20548 11868 20554 11870
rect 25221 11867 25287 11870
rect 33225 11867 33291 11870
rect 841 11794 907 11797
rect 6545 11794 6611 11797
rect 841 11792 6611 11794
rect 841 11736 846 11792
rect 902 11736 6550 11792
rect 6606 11736 6611 11792
rect 841 11734 6611 11736
rect 841 11731 907 11734
rect 6545 11731 6611 11734
rect 9489 11794 9555 11797
rect 13854 11794 13860 11796
rect 9489 11792 13860 11794
rect 9489 11736 9494 11792
rect 9550 11736 13860 11792
rect 9489 11734 13860 11736
rect 9489 11731 9555 11734
rect 13854 11732 13860 11734
rect 13924 11794 13930 11796
rect 15561 11794 15627 11797
rect 13924 11792 15627 11794
rect 13924 11736 15566 11792
rect 15622 11736 15627 11792
rect 13924 11734 15627 11736
rect 13924 11732 13930 11734
rect 15561 11731 15627 11734
rect 16021 11794 16087 11797
rect 17401 11794 17467 11797
rect 16021 11792 17467 11794
rect 16021 11736 16026 11792
rect 16082 11736 17406 11792
rect 17462 11736 17467 11792
rect 16021 11734 17467 11736
rect 16021 11731 16087 11734
rect 17401 11731 17467 11734
rect 19425 11792 19491 11797
rect 19425 11736 19430 11792
rect 19486 11736 19491 11792
rect 19425 11731 19491 11736
rect 19609 11794 19675 11797
rect 20294 11794 20300 11796
rect 19609 11792 20300 11794
rect 19609 11736 19614 11792
rect 19670 11736 20300 11792
rect 19609 11734 20300 11736
rect 19609 11731 19675 11734
rect 20294 11732 20300 11734
rect 20364 11732 20370 11796
rect 27981 11794 28047 11797
rect 20486 11792 28047 11794
rect 20486 11736 27986 11792
rect 28042 11736 28047 11792
rect 20486 11734 28047 11736
rect 3969 11658 4035 11661
rect 4981 11658 5047 11661
rect 3969 11656 5047 11658
rect 3969 11600 3974 11656
rect 4030 11600 4986 11656
rect 5042 11600 5047 11656
rect 3969 11598 5047 11600
rect 3969 11595 4035 11598
rect 4981 11595 5047 11598
rect 7833 11658 7899 11661
rect 20253 11658 20319 11661
rect 7833 11656 20319 11658
rect 7833 11600 7838 11656
rect 7894 11600 20258 11656
rect 20314 11600 20319 11656
rect 7833 11598 20319 11600
rect 7833 11595 7899 11598
rect 20253 11595 20319 11598
rect 0 11522 800 11552
rect 3785 11522 3851 11525
rect 0 11520 3851 11522
rect 0 11464 3790 11520
rect 3846 11464 3851 11520
rect 0 11462 3851 11464
rect 0 11432 800 11462
rect 3785 11459 3851 11462
rect 4838 11460 4844 11524
rect 4908 11522 4914 11524
rect 11881 11522 11947 11525
rect 4908 11520 11947 11522
rect 4908 11464 11886 11520
rect 11942 11464 11947 11520
rect 4908 11462 11947 11464
rect 4908 11460 4914 11462
rect 11881 11459 11947 11462
rect 14273 11522 14339 11525
rect 15745 11522 15811 11525
rect 20486 11522 20546 11734
rect 27981 11731 28047 11734
rect 29126 11732 29132 11796
rect 29196 11794 29202 11796
rect 42517 11794 42583 11797
rect 29196 11792 42583 11794
rect 29196 11736 42522 11792
rect 42578 11736 42583 11792
rect 29196 11734 42583 11736
rect 29196 11732 29202 11734
rect 42517 11731 42583 11734
rect 20805 11658 20871 11661
rect 30925 11658 30991 11661
rect 20805 11656 30991 11658
rect 20805 11600 20810 11656
rect 20866 11600 30930 11656
rect 30986 11600 30991 11656
rect 20805 11598 30991 11600
rect 20805 11595 20871 11598
rect 30925 11595 30991 11598
rect 31334 11596 31340 11660
rect 31404 11658 31410 11660
rect 42241 11658 42307 11661
rect 31404 11656 42307 11658
rect 31404 11600 42246 11656
rect 42302 11600 42307 11656
rect 31404 11598 42307 11600
rect 31404 11596 31410 11598
rect 42241 11595 42307 11598
rect 23565 11524 23631 11525
rect 23565 11522 23612 11524
rect 14273 11520 15811 11522
rect 14273 11464 14278 11520
rect 14334 11464 15750 11520
rect 15806 11464 15811 11520
rect 14273 11462 15811 11464
rect 14273 11459 14339 11462
rect 15745 11459 15811 11462
rect 16990 11462 20546 11522
rect 23520 11520 23612 11522
rect 23520 11464 23570 11520
rect 23520 11462 23612 11464
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 16990 11389 17050 11462
rect 23565 11460 23612 11462
rect 23676 11460 23682 11524
rect 23790 11460 23796 11524
rect 23860 11522 23866 11524
rect 24393 11522 24459 11525
rect 23860 11520 24459 11522
rect 23860 11464 24398 11520
rect 24454 11464 24459 11520
rect 23860 11462 24459 11464
rect 23860 11460 23866 11462
rect 23565 11459 23631 11460
rect 24393 11459 24459 11462
rect 29913 11522 29979 11525
rect 33910 11522 33916 11524
rect 29913 11520 33916 11522
rect 29913 11464 29918 11520
rect 29974 11464 33916 11520
rect 29913 11462 33916 11464
rect 29913 11459 29979 11462
rect 33910 11460 33916 11462
rect 33980 11460 33986 11524
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 2865 11384 2931 11389
rect 4889 11388 4955 11389
rect 2865 11328 2870 11384
rect 2926 11328 2931 11384
rect 2865 11323 2931 11328
rect 4838 11324 4844 11388
rect 4908 11386 4955 11388
rect 6269 11386 6335 11389
rect 4908 11384 5000 11386
rect 4950 11328 5000 11384
rect 4908 11326 5000 11328
rect 5766 11384 6335 11386
rect 5766 11328 6274 11384
rect 6330 11328 6335 11384
rect 5766 11326 6335 11328
rect 4908 11324 4955 11326
rect 4889 11323 4955 11324
rect 2868 11114 2928 11323
rect 4705 11114 4771 11117
rect 2868 11112 4771 11114
rect 2868 11056 4710 11112
rect 4766 11056 4771 11112
rect 2868 11054 4771 11056
rect 4705 11051 4771 11054
rect 5022 11052 5028 11116
rect 5092 11114 5098 11116
rect 5766 11114 5826 11326
rect 6269 11323 6335 11326
rect 7649 11386 7715 11389
rect 11278 11386 11284 11388
rect 7649 11384 11284 11386
rect 7649 11328 7654 11384
rect 7710 11328 11284 11384
rect 7649 11326 11284 11328
rect 7649 11323 7715 11326
rect 11278 11324 11284 11326
rect 11348 11324 11354 11388
rect 16990 11386 17099 11389
rect 12390 11384 17099 11386
rect 12390 11328 17038 11384
rect 17094 11328 17099 11384
rect 12390 11326 17099 11328
rect 5993 11250 6059 11253
rect 9949 11250 10015 11253
rect 5993 11248 10015 11250
rect 5993 11192 5998 11248
rect 6054 11192 9954 11248
rect 10010 11192 10015 11248
rect 5993 11190 10015 11192
rect 5993 11187 6059 11190
rect 9949 11187 10015 11190
rect 10174 11188 10180 11252
rect 10244 11250 10250 11252
rect 11421 11250 11487 11253
rect 10244 11248 11487 11250
rect 10244 11192 11426 11248
rect 11482 11192 11487 11248
rect 10244 11190 11487 11192
rect 10244 11188 10250 11190
rect 11421 11187 11487 11190
rect 6637 11114 6703 11117
rect 5092 11112 6703 11114
rect 5092 11056 6642 11112
rect 6698 11056 6703 11112
rect 5092 11054 6703 11056
rect 5092 11052 5098 11054
rect 6637 11051 6703 11054
rect 9765 11112 9831 11117
rect 9765 11056 9770 11112
rect 9826 11056 9831 11112
rect 9765 11051 9831 11056
rect 11329 11114 11395 11117
rect 12390 11114 12450 11326
rect 17033 11323 17099 11326
rect 17350 11324 17356 11388
rect 17420 11386 17426 11388
rect 17861 11386 17927 11389
rect 19885 11386 19951 11389
rect 17420 11384 17927 11386
rect 17420 11328 17866 11384
rect 17922 11328 17927 11384
rect 17420 11326 17927 11328
rect 17420 11324 17426 11326
rect 17861 11323 17927 11326
rect 18278 11384 19951 11386
rect 18278 11328 19890 11384
rect 19946 11328 19951 11384
rect 18278 11326 19951 11328
rect 12893 11252 12959 11253
rect 12893 11250 12940 11252
rect 12848 11248 12940 11250
rect 12848 11192 12898 11248
rect 12848 11190 12940 11192
rect 12893 11188 12940 11190
rect 13004 11188 13010 11252
rect 13997 11250 14063 11253
rect 14222 11250 14228 11252
rect 13997 11248 14228 11250
rect 13997 11192 14002 11248
rect 14058 11192 14228 11248
rect 13997 11190 14228 11192
rect 12893 11187 12959 11188
rect 13997 11187 14063 11190
rect 14222 11188 14228 11190
rect 14292 11188 14298 11252
rect 14406 11188 14412 11252
rect 14476 11250 14482 11252
rect 14825 11250 14891 11253
rect 16757 11250 16823 11253
rect 18278 11250 18338 11326
rect 19885 11323 19951 11326
rect 20069 11386 20135 11389
rect 21398 11386 21404 11388
rect 20069 11384 21404 11386
rect 20069 11328 20074 11384
rect 20130 11328 21404 11384
rect 20069 11326 21404 11328
rect 20069 11323 20135 11326
rect 21398 11324 21404 11326
rect 21468 11324 21474 11388
rect 24393 11386 24459 11389
rect 24526 11386 24532 11388
rect 24393 11384 24532 11386
rect 24393 11328 24398 11384
rect 24454 11328 24532 11384
rect 24393 11326 24532 11328
rect 24393 11323 24459 11326
rect 24526 11324 24532 11326
rect 24596 11324 24602 11388
rect 14476 11248 18338 11250
rect 14476 11192 14830 11248
rect 14886 11192 16762 11248
rect 16818 11192 18338 11248
rect 14476 11190 18338 11192
rect 18413 11250 18479 11253
rect 26233 11250 26299 11253
rect 18413 11248 26299 11250
rect 18413 11192 18418 11248
rect 18474 11192 26238 11248
rect 26294 11192 26299 11248
rect 18413 11190 26299 11192
rect 14476 11188 14482 11190
rect 14825 11187 14891 11190
rect 16757 11187 16823 11190
rect 18413 11187 18479 11190
rect 26233 11187 26299 11190
rect 16665 11114 16731 11117
rect 20253 11114 20319 11117
rect 20989 11114 21055 11117
rect 21449 11114 21515 11117
rect 11329 11112 12450 11114
rect 11329 11056 11334 11112
rect 11390 11056 12450 11112
rect 11329 11054 12450 11056
rect 14782 11112 16731 11114
rect 14782 11056 16670 11112
rect 16726 11056 16731 11112
rect 14782 11054 16731 11056
rect 11329 11051 11395 11054
rect 2630 10916 2636 10980
rect 2700 10978 2706 10980
rect 6361 10978 6427 10981
rect 2700 10976 6427 10978
rect 2700 10920 6366 10976
rect 6422 10920 6427 10976
rect 2700 10918 6427 10920
rect 9768 10978 9828 11051
rect 13169 10978 13235 10981
rect 14782 10978 14842 11054
rect 16665 11051 16731 11054
rect 19382 11054 20040 11114
rect 9768 10918 12450 10978
rect 2700 10916 2706 10918
rect 6361 10915 6427 10918
rect 0 10842 800 10872
rect 3141 10842 3207 10845
rect 0 10840 3207 10842
rect 0 10784 3146 10840
rect 3202 10784 3207 10840
rect 0 10782 3207 10784
rect 0 10752 800 10782
rect 3141 10779 3207 10782
rect 4153 10842 4219 10845
rect 4654 10842 4660 10844
rect 4153 10840 4660 10842
rect 4153 10784 4158 10840
rect 4214 10784 4660 10840
rect 4153 10782 4660 10784
rect 4153 10779 4219 10782
rect 4654 10780 4660 10782
rect 4724 10780 4730 10844
rect 6126 10780 6132 10844
rect 6196 10842 6202 10844
rect 6269 10842 6335 10845
rect 6196 10840 6335 10842
rect 6196 10784 6274 10840
rect 6330 10784 6335 10840
rect 6196 10782 6335 10784
rect 6196 10780 6202 10782
rect 6269 10779 6335 10782
rect 6453 10844 6519 10845
rect 6453 10840 6500 10844
rect 6564 10842 6570 10844
rect 7046 10842 7052 10844
rect 6453 10784 6458 10840
rect 6453 10780 6500 10784
rect 6564 10782 7052 10842
rect 6564 10780 6570 10782
rect 7046 10780 7052 10782
rect 7116 10780 7122 10844
rect 8201 10842 8267 10845
rect 9305 10842 9371 10845
rect 8201 10840 9371 10842
rect 8201 10784 8206 10840
rect 8262 10784 9310 10840
rect 9366 10784 9371 10840
rect 8201 10782 9371 10784
rect 12390 10842 12450 10918
rect 13169 10976 14842 10978
rect 13169 10920 13174 10976
rect 13230 10920 14842 10976
rect 13169 10918 14842 10920
rect 15009 10978 15075 10981
rect 16389 10978 16455 10981
rect 19057 10978 19123 10981
rect 15009 10976 19123 10978
rect 15009 10920 15014 10976
rect 15070 10920 16394 10976
rect 16450 10920 19062 10976
rect 19118 10920 19123 10976
rect 15009 10918 19123 10920
rect 13169 10915 13235 10918
rect 15009 10915 15075 10918
rect 16389 10915 16455 10918
rect 19057 10915 19123 10918
rect 15101 10842 15167 10845
rect 12390 10840 15167 10842
rect 12390 10784 15106 10840
rect 15162 10784 15167 10840
rect 12390 10782 15167 10784
rect 6453 10779 6519 10780
rect 8201 10779 8267 10782
rect 9305 10779 9371 10782
rect 15101 10779 15167 10782
rect 17217 10842 17283 10845
rect 19241 10844 19307 10845
rect 17534 10842 17540 10844
rect 17217 10840 17540 10842
rect 17217 10784 17222 10840
rect 17278 10784 17540 10840
rect 17217 10782 17540 10784
rect 17217 10779 17283 10782
rect 17534 10780 17540 10782
rect 17604 10780 17610 10844
rect 19190 10842 19196 10844
rect 19150 10782 19196 10842
rect 19260 10840 19307 10844
rect 19302 10784 19307 10840
rect 19190 10780 19196 10782
rect 19260 10780 19307 10784
rect 19241 10779 19307 10780
rect 1577 10706 1643 10709
rect 10777 10706 10843 10709
rect 1577 10704 10843 10706
rect 1577 10648 1582 10704
rect 1638 10648 10782 10704
rect 10838 10648 10843 10704
rect 1577 10646 10843 10648
rect 1577 10643 1643 10646
rect 10777 10643 10843 10646
rect 11094 10644 11100 10708
rect 11164 10706 11170 10708
rect 15285 10706 15351 10709
rect 19382 10706 19442 11054
rect 19980 10978 20040 11054
rect 20253 11112 21515 11114
rect 20253 11056 20258 11112
rect 20314 11056 20994 11112
rect 21050 11056 21454 11112
rect 21510 11056 21515 11112
rect 20253 11054 21515 11056
rect 20253 11051 20319 11054
rect 20989 11051 21055 11054
rect 21449 11051 21515 11054
rect 22553 11114 22619 11117
rect 30782 11114 30788 11116
rect 22553 11112 30788 11114
rect 22553 11056 22558 11112
rect 22614 11056 30788 11112
rect 22553 11054 30788 11056
rect 22553 11051 22619 11054
rect 30782 11052 30788 11054
rect 30852 11052 30858 11116
rect 20529 10978 20595 10981
rect 19980 10976 20595 10978
rect 19980 10920 20534 10976
rect 20590 10920 20595 10976
rect 19980 10918 20595 10920
rect 20529 10915 20595 10918
rect 20805 10978 20871 10981
rect 23422 10978 23428 10980
rect 20805 10976 23428 10978
rect 20805 10920 20810 10976
rect 20866 10920 23428 10976
rect 20805 10918 23428 10920
rect 20805 10915 20871 10918
rect 23422 10916 23428 10918
rect 23492 10916 23498 10980
rect 25681 10978 25747 10981
rect 43253 10978 43319 10981
rect 25681 10976 43319 10978
rect 25681 10920 25686 10976
rect 25742 10920 43258 10976
rect 43314 10920 43319 10976
rect 25681 10918 43319 10920
rect 25681 10915 25747 10918
rect 43253 10915 43319 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 19977 10842 20043 10845
rect 27705 10842 27771 10845
rect 19977 10840 27771 10842
rect 19977 10784 19982 10840
rect 20038 10784 27710 10840
rect 27766 10784 27771 10840
rect 19977 10782 27771 10784
rect 19977 10779 20043 10782
rect 27705 10779 27771 10782
rect 11164 10704 15351 10706
rect 11164 10648 15290 10704
rect 15346 10648 15351 10704
rect 11164 10646 15351 10648
rect 11164 10644 11170 10646
rect 15285 10643 15351 10646
rect 15518 10646 19442 10706
rect 19885 10706 19951 10709
rect 25221 10706 25287 10709
rect 19885 10704 25287 10706
rect 19885 10648 19890 10704
rect 19946 10648 25226 10704
rect 25282 10648 25287 10704
rect 19885 10646 25287 10648
rect 1577 10570 1643 10573
rect 1577 10568 7666 10570
rect 1577 10512 1582 10568
rect 1638 10512 7666 10568
rect 1577 10510 7666 10512
rect 1577 10507 1643 10510
rect 7606 10434 7666 10510
rect 7966 10508 7972 10572
rect 8036 10570 8042 10572
rect 9121 10570 9187 10573
rect 8036 10568 9187 10570
rect 8036 10512 9126 10568
rect 9182 10512 9187 10568
rect 8036 10510 9187 10512
rect 8036 10508 8042 10510
rect 9121 10507 9187 10510
rect 10225 10570 10291 10573
rect 12433 10570 12499 10573
rect 10225 10568 12499 10570
rect 10225 10512 10230 10568
rect 10286 10512 12438 10568
rect 12494 10512 12499 10568
rect 10225 10510 12499 10512
rect 10225 10507 10291 10510
rect 12433 10507 12499 10510
rect 12934 10508 12940 10572
rect 13004 10570 13010 10572
rect 13537 10570 13603 10573
rect 13997 10572 14063 10573
rect 13997 10570 14044 10572
rect 13004 10568 13603 10570
rect 13004 10512 13542 10568
rect 13598 10512 13603 10568
rect 13004 10510 13603 10512
rect 13952 10568 14044 10570
rect 13952 10512 14002 10568
rect 13952 10510 14044 10512
rect 13004 10508 13010 10510
rect 13537 10507 13603 10510
rect 13997 10508 14044 10510
rect 14108 10508 14114 10572
rect 14549 10570 14615 10573
rect 14774 10570 14780 10572
rect 14549 10568 14780 10570
rect 14549 10512 14554 10568
rect 14610 10512 14780 10568
rect 14549 10510 14780 10512
rect 13997 10507 14063 10508
rect 14549 10507 14615 10510
rect 14774 10508 14780 10510
rect 14844 10570 14850 10572
rect 15518 10570 15578 10646
rect 19885 10643 19951 10646
rect 25221 10643 25287 10646
rect 14844 10510 15578 10570
rect 16757 10570 16823 10573
rect 24669 10570 24735 10573
rect 35433 10570 35499 10573
rect 43345 10570 43411 10573
rect 16757 10568 22110 10570
rect 16757 10512 16762 10568
rect 16818 10512 22110 10568
rect 16757 10510 22110 10512
rect 14844 10508 14850 10510
rect 16757 10507 16823 10510
rect 14273 10434 14339 10437
rect 7606 10432 14339 10434
rect 7606 10376 14278 10432
rect 14334 10376 14339 10432
rect 7606 10374 14339 10376
rect 14273 10371 14339 10374
rect 15009 10434 15075 10437
rect 20897 10434 20963 10437
rect 21582 10434 21588 10436
rect 15009 10432 21588 10434
rect 15009 10376 15014 10432
rect 15070 10376 20902 10432
rect 20958 10376 21588 10432
rect 15009 10374 21588 10376
rect 15009 10371 15075 10374
rect 20897 10371 20963 10374
rect 21582 10372 21588 10374
rect 21652 10372 21658 10436
rect 21766 10372 21772 10436
rect 21836 10434 21842 10436
rect 21909 10434 21975 10437
rect 21836 10432 21975 10434
rect 21836 10376 21914 10432
rect 21970 10376 21975 10432
rect 21836 10374 21975 10376
rect 22050 10434 22110 10510
rect 24669 10568 43411 10570
rect 24669 10512 24674 10568
rect 24730 10512 35438 10568
rect 35494 10512 43350 10568
rect 43406 10512 43411 10568
rect 24669 10510 43411 10512
rect 24669 10507 24735 10510
rect 35433 10507 35499 10510
rect 43345 10507 43411 10510
rect 24945 10434 25011 10437
rect 22050 10432 25011 10434
rect 22050 10376 24950 10432
rect 25006 10376 25011 10432
rect 22050 10374 25011 10376
rect 21836 10372 21842 10374
rect 21909 10371 21975 10374
rect 24945 10371 25011 10374
rect 25221 10434 25287 10437
rect 33685 10434 33751 10437
rect 25221 10432 33751 10434
rect 25221 10376 25226 10432
rect 25282 10376 33690 10432
rect 33746 10376 33751 10432
rect 25221 10374 33751 10376
rect 25221 10371 25287 10374
rect 33685 10371 33751 10374
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 1853 10298 1919 10301
rect 0 10296 1919 10298
rect 0 10240 1858 10296
rect 1914 10240 1919 10296
rect 0 10238 1919 10240
rect 0 10208 800 10238
rect 1853 10235 1919 10238
rect 7414 10236 7420 10300
rect 7484 10298 7490 10300
rect 8017 10298 8083 10301
rect 7484 10296 8083 10298
rect 7484 10240 8022 10296
rect 8078 10240 8083 10296
rect 7484 10238 8083 10240
rect 7484 10236 7490 10238
rect 8017 10235 8083 10238
rect 8937 10298 9003 10301
rect 9254 10298 9260 10300
rect 8937 10296 9260 10298
rect 8937 10240 8942 10296
rect 8998 10240 9260 10296
rect 8937 10238 9260 10240
rect 8937 10235 9003 10238
rect 9254 10236 9260 10238
rect 9324 10236 9330 10300
rect 9806 10236 9812 10300
rect 9876 10298 9882 10300
rect 11053 10298 11119 10301
rect 16665 10298 16731 10301
rect 9876 10296 11119 10298
rect 9876 10240 11058 10296
rect 11114 10240 11119 10296
rect 9876 10238 11119 10240
rect 9876 10236 9882 10238
rect 11053 10235 11119 10238
rect 11286 10296 16731 10298
rect 11286 10240 16670 10296
rect 16726 10240 16731 10296
rect 11286 10238 16731 10240
rect 2129 10162 2195 10165
rect 2446 10162 2452 10164
rect 2129 10160 2452 10162
rect 2129 10104 2134 10160
rect 2190 10104 2452 10160
rect 2129 10102 2452 10104
rect 2129 10099 2195 10102
rect 2446 10100 2452 10102
rect 2516 10100 2522 10164
rect 2589 10162 2655 10165
rect 11145 10162 11211 10165
rect 2589 10160 11211 10162
rect 2589 10104 2594 10160
rect 2650 10104 11150 10160
rect 11206 10104 11211 10160
rect 2589 10102 11211 10104
rect 2589 10099 2655 10102
rect 11145 10099 11211 10102
rect 3601 10026 3667 10029
rect 4654 10026 4660 10028
rect 3601 10024 4660 10026
rect 3601 9968 3606 10024
rect 3662 9968 4660 10024
rect 3601 9966 4660 9968
rect 3601 9963 3667 9966
rect 4654 9964 4660 9966
rect 4724 10026 4730 10028
rect 6913 10026 6979 10029
rect 8017 10026 8083 10029
rect 4724 10024 8083 10026
rect 4724 9968 6918 10024
rect 6974 9968 8022 10024
rect 8078 9968 8083 10024
rect 4724 9966 8083 9968
rect 4724 9964 4730 9966
rect 6913 9963 6979 9966
rect 8017 9963 8083 9966
rect 8150 9964 8156 10028
rect 8220 10026 8226 10028
rect 9029 10026 9095 10029
rect 11286 10026 11346 10238
rect 16665 10235 16731 10238
rect 16849 10298 16915 10301
rect 17350 10298 17356 10300
rect 16849 10296 17356 10298
rect 16849 10240 16854 10296
rect 16910 10240 17356 10296
rect 16849 10238 17356 10240
rect 16849 10235 16915 10238
rect 17350 10236 17356 10238
rect 17420 10236 17426 10300
rect 18137 10298 18203 10301
rect 20478 10298 20484 10300
rect 18137 10296 20484 10298
rect 18137 10240 18142 10296
rect 18198 10240 20484 10296
rect 18137 10238 20484 10240
rect 18137 10235 18203 10238
rect 20478 10236 20484 10238
rect 20548 10236 20554 10300
rect 21173 10298 21239 10301
rect 31518 10298 31524 10300
rect 21173 10296 31524 10298
rect 21173 10240 21178 10296
rect 21234 10240 31524 10296
rect 21173 10238 31524 10240
rect 21173 10235 21239 10238
rect 31518 10236 31524 10238
rect 31588 10236 31594 10300
rect 12433 10162 12499 10165
rect 13169 10162 13235 10165
rect 12433 10160 13235 10162
rect 12433 10104 12438 10160
rect 12494 10104 13174 10160
rect 13230 10104 13235 10160
rect 12433 10102 13235 10104
rect 12433 10099 12499 10102
rect 13169 10099 13235 10102
rect 14457 10162 14523 10165
rect 20069 10162 20135 10165
rect 14457 10160 20135 10162
rect 14457 10104 14462 10160
rect 14518 10104 20074 10160
rect 20130 10104 20135 10160
rect 14457 10102 20135 10104
rect 14457 10099 14523 10102
rect 20069 10099 20135 10102
rect 20529 10162 20595 10165
rect 25681 10162 25747 10165
rect 27153 10162 27219 10165
rect 28993 10164 29059 10165
rect 20529 10160 25747 10162
rect 20529 10104 20534 10160
rect 20590 10104 25686 10160
rect 25742 10104 25747 10160
rect 20529 10102 25747 10104
rect 20529 10099 20595 10102
rect 25681 10099 25747 10102
rect 25822 10160 27219 10162
rect 25822 10104 27158 10160
rect 27214 10104 27219 10160
rect 25822 10102 27219 10104
rect 8220 10024 11346 10026
rect 8220 9968 9034 10024
rect 9090 9968 11346 10024
rect 8220 9966 11346 9968
rect 11881 10026 11947 10029
rect 12382 10026 12388 10028
rect 11881 10024 12388 10026
rect 11881 9968 11886 10024
rect 11942 9968 12388 10024
rect 11881 9966 12388 9968
rect 8220 9964 8226 9966
rect 9029 9963 9095 9966
rect 11881 9963 11947 9966
rect 12382 9964 12388 9966
rect 12452 9964 12458 10028
rect 12985 10026 13051 10029
rect 15929 10026 15995 10029
rect 12985 10024 15995 10026
rect 12985 9968 12990 10024
rect 13046 9968 15934 10024
rect 15990 9968 15995 10024
rect 12985 9966 15995 9968
rect 12985 9963 13051 9966
rect 15929 9963 15995 9966
rect 16113 10026 16179 10029
rect 17217 10026 17283 10029
rect 16113 10024 17283 10026
rect 16113 9968 16118 10024
rect 16174 9968 17222 10024
rect 17278 9968 17283 10024
rect 16113 9966 17283 9968
rect 16113 9963 16179 9966
rect 17217 9963 17283 9966
rect 18781 10026 18847 10029
rect 25822 10026 25882 10102
rect 27153 10099 27219 10102
rect 28942 10100 28948 10164
rect 29012 10162 29059 10164
rect 29012 10160 29104 10162
rect 29054 10104 29104 10160
rect 29012 10102 29104 10104
rect 29012 10100 29059 10102
rect 28993 10099 29059 10100
rect 18781 10024 25882 10026
rect 18781 9968 18786 10024
rect 18842 9968 25882 10024
rect 18781 9966 25882 9968
rect 26233 10026 26299 10029
rect 38009 10026 38075 10029
rect 26233 10024 38075 10026
rect 26233 9968 26238 10024
rect 26294 9968 38014 10024
rect 38070 9968 38075 10024
rect 26233 9966 38075 9968
rect 18781 9963 18847 9966
rect 26233 9963 26299 9966
rect 38009 9963 38075 9966
rect 44081 10026 44147 10029
rect 45200 10026 46000 10056
rect 44081 10024 46000 10026
rect 44081 9968 44086 10024
rect 44142 9968 46000 10024
rect 44081 9966 46000 9968
rect 44081 9963 44147 9966
rect 45200 9936 46000 9966
rect 5206 9828 5212 9892
rect 5276 9890 5282 9892
rect 8702 9890 8708 9892
rect 5276 9830 8708 9890
rect 5276 9828 5282 9830
rect 8702 9828 8708 9830
rect 8772 9890 8778 9892
rect 8937 9890 9003 9893
rect 8772 9888 9003 9890
rect 8772 9832 8942 9888
rect 8998 9832 9003 9888
rect 8772 9830 9003 9832
rect 8772 9828 8778 9830
rect 8937 9827 9003 9830
rect 9213 9890 9279 9893
rect 9438 9890 9444 9892
rect 9213 9888 9444 9890
rect 9213 9832 9218 9888
rect 9274 9832 9444 9888
rect 9213 9830 9444 9832
rect 9213 9827 9279 9830
rect 9438 9828 9444 9830
rect 9508 9828 9514 9892
rect 9949 9890 10015 9893
rect 11513 9890 11579 9893
rect 9949 9888 12450 9890
rect 9949 9832 9954 9888
rect 10010 9832 11518 9888
rect 11574 9832 12450 9888
rect 9949 9830 12450 9832
rect 9949 9827 10015 9830
rect 11513 9827 11579 9830
rect 0 9754 800 9784
rect 2865 9754 2931 9757
rect 3601 9756 3667 9757
rect 3182 9754 3188 9756
rect 0 9752 3188 9754
rect 0 9696 2870 9752
rect 2926 9696 3188 9752
rect 0 9694 3188 9696
rect 0 9664 800 9694
rect 2865 9691 2931 9694
rect 3182 9692 3188 9694
rect 3252 9692 3258 9756
rect 3550 9692 3556 9756
rect 3620 9754 3667 9756
rect 3877 9754 3943 9757
rect 10317 9754 10383 9757
rect 3620 9752 3712 9754
rect 3662 9696 3712 9752
rect 3620 9694 3712 9696
rect 3877 9752 10383 9754
rect 3877 9696 3882 9752
rect 3938 9696 10322 9752
rect 10378 9696 10383 9752
rect 3877 9694 10383 9696
rect 3620 9692 3667 9694
rect 3601 9691 3667 9692
rect 3877 9691 3943 9694
rect 10317 9691 10383 9694
rect 11973 9754 12039 9757
rect 12390 9754 12450 9830
rect 13302 9828 13308 9892
rect 13372 9890 13378 9892
rect 13629 9890 13695 9893
rect 14457 9892 14523 9893
rect 13372 9888 13695 9890
rect 13372 9832 13634 9888
rect 13690 9832 13695 9888
rect 13372 9830 13695 9832
rect 13372 9828 13378 9830
rect 13629 9827 13695 9830
rect 14406 9828 14412 9892
rect 14476 9890 14523 9892
rect 16757 9890 16823 9893
rect 19006 9890 19012 9892
rect 14476 9888 14568 9890
rect 14518 9832 14568 9888
rect 14476 9830 14568 9832
rect 16757 9888 19012 9890
rect 16757 9832 16762 9888
rect 16818 9832 19012 9888
rect 16757 9830 19012 9832
rect 14476 9828 14523 9830
rect 14457 9827 14523 9828
rect 16757 9827 16823 9830
rect 19006 9828 19012 9830
rect 19076 9828 19082 9892
rect 20294 9828 20300 9892
rect 20364 9890 20370 9892
rect 20529 9890 20595 9893
rect 20364 9888 20595 9890
rect 20364 9832 20534 9888
rect 20590 9832 20595 9888
rect 20364 9830 20595 9832
rect 20364 9828 20370 9830
rect 20529 9827 20595 9830
rect 20897 9890 20963 9893
rect 21173 9890 21239 9893
rect 20897 9888 21239 9890
rect 20897 9832 20902 9888
rect 20958 9832 21178 9888
rect 21234 9832 21239 9888
rect 20897 9830 21239 9832
rect 20897 9827 20963 9830
rect 21173 9827 21239 9830
rect 25497 9890 25563 9893
rect 31845 9890 31911 9893
rect 25497 9888 31911 9890
rect 25497 9832 25502 9888
rect 25558 9832 31850 9888
rect 31906 9832 31911 9888
rect 25497 9830 31911 9832
rect 25497 9827 25563 9830
rect 31845 9827 31911 9830
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 16665 9754 16731 9757
rect 11973 9752 12266 9754
rect 11973 9696 11978 9752
rect 12034 9696 12266 9752
rect 11973 9694 12266 9696
rect 12390 9752 16731 9754
rect 12390 9696 16670 9752
rect 16726 9696 16731 9752
rect 12390 9694 16731 9696
rect 11973 9691 12039 9694
rect 1158 9556 1164 9620
rect 1228 9618 1234 9620
rect 1485 9618 1551 9621
rect 1228 9616 1551 9618
rect 1228 9560 1490 9616
rect 1546 9560 1551 9616
rect 1228 9558 1551 9560
rect 1228 9556 1234 9558
rect 1485 9555 1551 9558
rect 3877 9618 3943 9621
rect 4521 9618 4587 9621
rect 3877 9616 4587 9618
rect 3877 9560 3882 9616
rect 3938 9560 4526 9616
rect 4582 9560 4587 9616
rect 3877 9558 4587 9560
rect 3877 9555 3943 9558
rect 4521 9555 4587 9558
rect 5533 9618 5599 9621
rect 6085 9618 6151 9621
rect 5533 9616 6151 9618
rect 5533 9560 5538 9616
rect 5594 9560 6090 9616
rect 6146 9560 6151 9616
rect 5533 9558 6151 9560
rect 5533 9555 5599 9558
rect 6085 9555 6151 9558
rect 6913 9618 6979 9621
rect 7782 9618 7788 9620
rect 6913 9616 7788 9618
rect 6913 9560 6918 9616
rect 6974 9560 7788 9616
rect 6913 9558 7788 9560
rect 6913 9555 6979 9558
rect 7782 9556 7788 9558
rect 7852 9556 7858 9620
rect 8017 9618 8083 9621
rect 11605 9618 11671 9621
rect 8017 9616 11671 9618
rect 8017 9560 8022 9616
rect 8078 9560 11610 9616
rect 11666 9560 11671 9616
rect 8017 9558 11671 9560
rect 8017 9555 8083 9558
rect 11605 9555 11671 9558
rect 11973 9620 12039 9621
rect 11973 9616 12020 9620
rect 12084 9618 12090 9620
rect 12206 9618 12266 9694
rect 16665 9691 16731 9694
rect 18505 9754 18571 9757
rect 19425 9754 19491 9757
rect 18505 9752 19491 9754
rect 18505 9696 18510 9752
rect 18566 9696 19430 9752
rect 19486 9696 19491 9752
rect 18505 9694 19491 9696
rect 18505 9691 18571 9694
rect 19425 9691 19491 9694
rect 20478 9692 20484 9756
rect 20548 9754 20554 9756
rect 21030 9754 21036 9756
rect 20548 9694 21036 9754
rect 20548 9692 20554 9694
rect 21030 9692 21036 9694
rect 21100 9692 21106 9756
rect 15745 9618 15811 9621
rect 11973 9560 11978 9616
rect 11973 9556 12020 9560
rect 12084 9558 12130 9618
rect 12206 9616 15811 9618
rect 12206 9560 15750 9616
rect 15806 9560 15811 9616
rect 12206 9558 15811 9560
rect 12084 9556 12090 9558
rect 11973 9555 12039 9556
rect 15745 9555 15811 9558
rect 16941 9618 17007 9621
rect 24209 9620 24275 9621
rect 17166 9618 17172 9620
rect 16941 9616 17172 9618
rect 16941 9560 16946 9616
rect 17002 9560 17172 9616
rect 16941 9558 17172 9560
rect 16941 9555 17007 9558
rect 17166 9556 17172 9558
rect 17236 9556 17242 9620
rect 18822 9618 18828 9620
rect 17358 9558 18828 9618
rect 3509 9482 3575 9485
rect 11789 9482 11855 9485
rect 14917 9482 14983 9485
rect 3509 9480 11855 9482
rect 3509 9424 3514 9480
rect 3570 9424 11794 9480
rect 11850 9424 11855 9480
rect 3509 9422 11855 9424
rect 3509 9419 3575 9422
rect 11789 9419 11855 9422
rect 11976 9480 14983 9482
rect 11976 9424 14922 9480
rect 14978 9424 14983 9480
rect 11976 9422 14983 9424
rect 5349 9346 5415 9349
rect 8845 9346 8911 9349
rect 9121 9346 9187 9349
rect 5349 9344 8402 9346
rect 5349 9288 5354 9344
rect 5410 9288 8402 9344
rect 5349 9286 8402 9288
rect 5349 9283 5415 9286
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 5942 9148 5948 9212
rect 6012 9210 6018 9212
rect 6085 9210 6151 9213
rect 6637 9210 6703 9213
rect 7741 9210 7807 9213
rect 6012 9208 6151 9210
rect 6012 9152 6090 9208
rect 6146 9152 6151 9208
rect 6012 9150 6151 9152
rect 6012 9148 6018 9150
rect 6085 9147 6151 9150
rect 6502 9208 6703 9210
rect 6502 9152 6642 9208
rect 6698 9152 6703 9208
rect 6502 9150 6703 9152
rect 0 9074 800 9104
rect 6502 9074 6562 9150
rect 6637 9147 6703 9150
rect 6870 9208 7807 9210
rect 6870 9152 7746 9208
rect 7802 9152 7807 9208
rect 6870 9150 7807 9152
rect 0 9014 6562 9074
rect 0 8984 800 9014
rect 1393 8940 1459 8941
rect 1342 8938 1348 8940
rect 1302 8878 1348 8938
rect 1412 8936 1459 8940
rect 5574 8938 5580 8940
rect 1454 8880 1459 8936
rect 1342 8876 1348 8878
rect 1412 8876 1459 8880
rect 1393 8875 1459 8876
rect 1534 8878 5580 8938
rect 974 8740 980 8804
rect 1044 8802 1050 8804
rect 1534 8802 1594 8878
rect 5574 8876 5580 8878
rect 5644 8938 5650 8940
rect 6177 8938 6243 8941
rect 5644 8936 6243 8938
rect 5644 8880 6182 8936
rect 6238 8880 6243 8936
rect 5644 8878 6243 8880
rect 6870 8938 6930 9150
rect 7741 9147 7807 9150
rect 7966 9148 7972 9212
rect 8036 9210 8042 9212
rect 8109 9210 8175 9213
rect 8036 9208 8175 9210
rect 8036 9152 8114 9208
rect 8170 9152 8175 9208
rect 8036 9150 8175 9152
rect 8342 9210 8402 9286
rect 8845 9344 9187 9346
rect 8845 9288 8850 9344
rect 8906 9288 9126 9344
rect 9182 9288 9187 9344
rect 8845 9286 9187 9288
rect 8845 9283 8911 9286
rect 9121 9283 9187 9286
rect 9397 9346 9463 9349
rect 11976 9346 12036 9422
rect 14917 9419 14983 9422
rect 15653 9482 15719 9485
rect 16614 9482 16620 9484
rect 15653 9480 16620 9482
rect 15653 9424 15658 9480
rect 15714 9424 16620 9480
rect 15653 9422 16620 9424
rect 15653 9419 15719 9422
rect 16614 9420 16620 9422
rect 16684 9420 16690 9484
rect 17033 9482 17099 9485
rect 17358 9482 17418 9558
rect 18822 9556 18828 9558
rect 18892 9556 18898 9620
rect 19006 9556 19012 9620
rect 19076 9618 19082 9620
rect 23422 9618 23428 9620
rect 19076 9558 23428 9618
rect 19076 9556 19082 9558
rect 23422 9556 23428 9558
rect 23492 9556 23498 9620
rect 24158 9556 24164 9620
rect 24228 9618 24275 9620
rect 24228 9616 24320 9618
rect 24270 9560 24320 9616
rect 24228 9558 24320 9560
rect 24228 9556 24275 9558
rect 25814 9556 25820 9620
rect 25884 9618 25890 9620
rect 25957 9618 26023 9621
rect 25884 9616 26023 9618
rect 25884 9560 25962 9616
rect 26018 9560 26023 9616
rect 25884 9558 26023 9560
rect 25884 9556 25890 9558
rect 24209 9555 24275 9556
rect 25957 9555 26023 9558
rect 17033 9480 17418 9482
rect 17033 9424 17038 9480
rect 17094 9424 17418 9480
rect 17033 9422 17418 9424
rect 17585 9482 17651 9485
rect 18597 9484 18663 9485
rect 18270 9482 18276 9484
rect 17585 9480 18276 9482
rect 17585 9424 17590 9480
rect 17646 9424 18276 9480
rect 17585 9422 18276 9424
rect 17033 9419 17099 9422
rect 17585 9419 17651 9422
rect 18270 9420 18276 9422
rect 18340 9420 18346 9484
rect 18597 9480 18644 9484
rect 18708 9482 18714 9484
rect 19517 9482 19583 9485
rect 24853 9482 24919 9485
rect 32070 9482 32076 9484
rect 18597 9424 18602 9480
rect 18597 9420 18644 9424
rect 18708 9422 18754 9482
rect 19517 9480 23306 9482
rect 19517 9424 19522 9480
rect 19578 9424 23306 9480
rect 19517 9422 23306 9424
rect 18708 9420 18714 9422
rect 18597 9419 18663 9420
rect 19517 9419 19583 9422
rect 12893 9346 12959 9349
rect 17718 9346 17724 9348
rect 9397 9344 12036 9346
rect 9397 9288 9402 9344
rect 9458 9288 12036 9344
rect 9397 9286 12036 9288
rect 12436 9344 12959 9346
rect 12436 9288 12898 9344
rect 12954 9288 12959 9344
rect 12436 9286 12959 9288
rect 9397 9283 9463 9286
rect 8477 9210 8543 9213
rect 8342 9208 8543 9210
rect 8342 9152 8482 9208
rect 8538 9152 8543 9208
rect 8342 9150 8543 9152
rect 8036 9148 8042 9150
rect 8109 9147 8175 9150
rect 8477 9147 8543 9150
rect 8661 9212 8727 9213
rect 8661 9208 8708 9212
rect 8772 9210 8778 9212
rect 12436 9210 12496 9286
rect 12893 9283 12959 9286
rect 16760 9286 17724 9346
rect 16760 9213 16820 9286
rect 17718 9284 17724 9286
rect 17788 9284 17794 9348
rect 17861 9346 17927 9349
rect 23054 9346 23060 9348
rect 17861 9344 23060 9346
rect 17861 9288 17866 9344
rect 17922 9288 23060 9344
rect 17861 9286 23060 9288
rect 17861 9283 17927 9286
rect 23054 9284 23060 9286
rect 23124 9284 23130 9348
rect 23246 9346 23306 9422
rect 24853 9480 32076 9482
rect 24853 9424 24858 9480
rect 24914 9424 32076 9480
rect 24853 9422 32076 9424
rect 24853 9419 24919 9422
rect 32070 9420 32076 9422
rect 32140 9420 32146 9484
rect 25037 9346 25103 9349
rect 23246 9344 25103 9346
rect 23246 9288 25042 9344
rect 25098 9288 25103 9344
rect 23246 9286 25103 9288
rect 25037 9283 25103 9286
rect 25221 9346 25287 9349
rect 31661 9346 31727 9349
rect 25221 9344 31727 9346
rect 25221 9288 25226 9344
rect 25282 9288 31666 9344
rect 31722 9288 31727 9344
rect 25221 9286 31727 9288
rect 25221 9283 25287 9286
rect 31661 9283 31727 9286
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 8661 9152 8666 9208
rect 8661 9148 8708 9152
rect 8772 9150 12496 9210
rect 12617 9210 12683 9213
rect 12750 9210 12756 9212
rect 12617 9208 12756 9210
rect 12617 9152 12622 9208
rect 12678 9152 12756 9208
rect 12617 9150 12756 9152
rect 8772 9148 8778 9150
rect 8661 9147 8727 9148
rect 12617 9147 12683 9150
rect 12750 9148 12756 9150
rect 12820 9148 12826 9212
rect 16246 9148 16252 9212
rect 16316 9210 16322 9212
rect 16481 9210 16547 9213
rect 16316 9208 16547 9210
rect 16316 9152 16486 9208
rect 16542 9152 16547 9208
rect 16316 9150 16547 9152
rect 16316 9148 16322 9150
rect 16481 9147 16547 9150
rect 16757 9208 16823 9213
rect 16757 9152 16762 9208
rect 16818 9152 16823 9208
rect 16757 9147 16823 9152
rect 17033 9210 17099 9213
rect 18045 9212 18111 9213
rect 17534 9210 17540 9212
rect 17033 9208 17540 9210
rect 17033 9152 17038 9208
rect 17094 9152 17540 9208
rect 17033 9150 17540 9152
rect 17033 9147 17099 9150
rect 17534 9148 17540 9150
rect 17604 9148 17610 9212
rect 18045 9208 18092 9212
rect 18156 9210 18162 9212
rect 19149 9210 19215 9213
rect 22093 9210 22159 9213
rect 18045 9152 18050 9208
rect 18045 9148 18092 9152
rect 18156 9150 18202 9210
rect 19149 9208 22159 9210
rect 19149 9152 19154 9208
rect 19210 9152 22098 9208
rect 22154 9152 22159 9208
rect 19149 9150 22159 9152
rect 18156 9148 18162 9150
rect 18045 9147 18111 9148
rect 19149 9147 19215 9150
rect 22093 9147 22159 9150
rect 22553 9210 22619 9213
rect 25262 9210 25268 9212
rect 22553 9208 25268 9210
rect 22553 9152 22558 9208
rect 22614 9152 25268 9208
rect 22553 9150 25268 9152
rect 22553 9147 22619 9150
rect 25262 9148 25268 9150
rect 25332 9148 25338 9212
rect 26182 9148 26188 9212
rect 26252 9210 26258 9212
rect 33593 9210 33659 9213
rect 26252 9208 33659 9210
rect 26252 9152 33598 9208
rect 33654 9152 33659 9208
rect 26252 9150 33659 9152
rect 26252 9148 26258 9150
rect 33593 9147 33659 9150
rect 7005 9074 7071 9077
rect 10133 9074 10199 9077
rect 7005 9072 10199 9074
rect 7005 9016 7010 9072
rect 7066 9016 10138 9072
rect 10194 9016 10199 9072
rect 7005 9014 10199 9016
rect 7005 9011 7071 9014
rect 10133 9011 10199 9014
rect 10542 9012 10548 9076
rect 10612 9074 10618 9076
rect 19057 9074 19123 9077
rect 10612 9072 19123 9074
rect 10612 9016 19062 9072
rect 19118 9016 19123 9072
rect 10612 9014 19123 9016
rect 10612 9012 10618 9014
rect 19057 9011 19123 9014
rect 19885 9074 19951 9077
rect 22185 9074 22251 9077
rect 19885 9072 22251 9074
rect 19885 9016 19890 9072
rect 19946 9016 22190 9072
rect 22246 9016 22251 9072
rect 19885 9014 22251 9016
rect 19885 9011 19951 9014
rect 22185 9011 22251 9014
rect 22553 9074 22619 9077
rect 34697 9074 34763 9077
rect 22553 9072 34763 9074
rect 22553 9016 22558 9072
rect 22614 9016 34702 9072
rect 34758 9016 34763 9072
rect 22553 9014 34763 9016
rect 22553 9011 22619 9014
rect 34697 9011 34763 9014
rect 7097 8938 7163 8941
rect 7373 8940 7439 8941
rect 7373 8938 7420 8940
rect 6870 8936 7163 8938
rect 6870 8880 7102 8936
rect 7158 8880 7163 8936
rect 6870 8878 7163 8880
rect 7328 8936 7420 8938
rect 7328 8880 7378 8936
rect 7328 8878 7420 8880
rect 5644 8876 5650 8878
rect 6177 8875 6243 8878
rect 7097 8875 7163 8878
rect 7373 8876 7420 8878
rect 7484 8876 7490 8940
rect 16798 8938 16804 8940
rect 7606 8878 16804 8938
rect 7373 8875 7439 8876
rect 1044 8742 1594 8802
rect 1945 8802 2011 8805
rect 7606 8802 7666 8878
rect 16798 8876 16804 8878
rect 16868 8876 16874 8940
rect 18321 8938 18387 8941
rect 21357 8938 21423 8941
rect 16990 8878 17786 8938
rect 1945 8800 7666 8802
rect 1945 8744 1950 8800
rect 2006 8744 7666 8800
rect 1945 8742 7666 8744
rect 7741 8802 7807 8805
rect 16990 8802 17050 8878
rect 7741 8800 17050 8802
rect 7741 8744 7746 8800
rect 7802 8744 17050 8800
rect 7741 8742 17050 8744
rect 17726 8802 17786 8878
rect 18321 8936 21423 8938
rect 18321 8880 18326 8936
rect 18382 8880 21362 8936
rect 21418 8880 21423 8936
rect 18321 8878 21423 8880
rect 18321 8875 18387 8878
rect 21357 8875 21423 8878
rect 24485 8938 24551 8941
rect 43069 8938 43135 8941
rect 24485 8936 43135 8938
rect 24485 8880 24490 8936
rect 24546 8880 43074 8936
rect 43130 8880 43135 8936
rect 24485 8878 43135 8880
rect 24485 8875 24551 8878
rect 43069 8875 43135 8878
rect 18965 8802 19031 8805
rect 17726 8800 19031 8802
rect 17726 8744 18970 8800
rect 19026 8744 19031 8800
rect 17726 8742 19031 8744
rect 1044 8740 1050 8742
rect 1945 8739 2011 8742
rect 7741 8739 7807 8742
rect 18965 8739 19031 8742
rect 21449 8802 21515 8805
rect 24853 8802 24919 8805
rect 21449 8800 24919 8802
rect 21449 8744 21454 8800
rect 21510 8744 24858 8800
rect 24914 8744 24919 8800
rect 21449 8742 24919 8744
rect 21449 8739 21515 8742
rect 24853 8739 24919 8742
rect 25037 8802 25103 8805
rect 32673 8802 32739 8805
rect 25037 8800 32739 8802
rect 25037 8744 25042 8800
rect 25098 8744 32678 8800
rect 32734 8744 32739 8800
rect 25037 8742 32739 8744
rect 25037 8739 25103 8742
rect 32673 8739 32739 8742
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 2221 8666 2287 8669
rect 2998 8666 3004 8668
rect 2221 8664 3004 8666
rect 2221 8608 2226 8664
rect 2282 8608 3004 8664
rect 2221 8606 3004 8608
rect 2221 8603 2287 8606
rect 2998 8604 3004 8606
rect 3068 8604 3074 8668
rect 3417 8666 3483 8669
rect 10869 8666 10935 8669
rect 3417 8664 10935 8666
rect 3417 8608 3422 8664
rect 3478 8608 10874 8664
rect 10930 8608 10935 8664
rect 3417 8606 10935 8608
rect 3417 8603 3483 8606
rect 10869 8603 10935 8606
rect 11053 8666 11119 8669
rect 13721 8666 13787 8669
rect 11053 8664 13787 8666
rect 11053 8608 11058 8664
rect 11114 8608 13726 8664
rect 13782 8608 13787 8664
rect 11053 8606 13787 8608
rect 11053 8603 11119 8606
rect 13721 8603 13787 8606
rect 14089 8666 14155 8669
rect 17401 8666 17467 8669
rect 19149 8666 19215 8669
rect 14089 8664 17280 8666
rect 14089 8608 14094 8664
rect 14150 8608 17280 8664
rect 14089 8606 17280 8608
rect 14089 8603 14155 8606
rect 0 8530 800 8560
rect 1761 8530 1827 8533
rect 6678 8530 6684 8532
rect 0 8528 1827 8530
rect 0 8472 1766 8528
rect 1822 8472 1827 8528
rect 0 8470 1827 8472
rect 0 8440 800 8470
rect 1761 8467 1827 8470
rect 3926 8470 6684 8530
rect 1894 8332 1900 8396
rect 1964 8394 1970 8396
rect 2037 8394 2103 8397
rect 1964 8392 2103 8394
rect 1964 8336 2042 8392
rect 2098 8336 2103 8392
rect 1964 8334 2103 8336
rect 1964 8332 1970 8334
rect 2037 8331 2103 8334
rect 2262 8196 2268 8260
rect 2332 8258 2338 8260
rect 2589 8258 2655 8261
rect 2332 8256 2655 8258
rect 2332 8200 2594 8256
rect 2650 8200 2655 8256
rect 2332 8198 2655 8200
rect 2332 8196 2338 8198
rect 2589 8195 2655 8198
rect 2681 8124 2747 8125
rect 2630 8122 2636 8124
rect 2590 8062 2636 8122
rect 2700 8120 2747 8124
rect 2742 8064 2747 8120
rect 2630 8060 2636 8062
rect 2700 8060 2747 8064
rect 2681 8059 2747 8060
rect 0 7986 800 8016
rect 3926 7986 3986 8470
rect 6678 8468 6684 8470
rect 6748 8530 6754 8532
rect 9949 8530 10015 8533
rect 6748 8528 10015 8530
rect 6748 8472 9954 8528
rect 10010 8472 10015 8528
rect 6748 8470 10015 8472
rect 6748 8468 6754 8470
rect 9949 8467 10015 8470
rect 10869 8530 10935 8533
rect 16941 8530 17007 8533
rect 10869 8528 17007 8530
rect 10869 8472 10874 8528
rect 10930 8472 16946 8528
rect 17002 8472 17007 8528
rect 10869 8470 17007 8472
rect 10869 8467 10935 8470
rect 16941 8467 17007 8470
rect 6177 8394 6243 8397
rect 9806 8394 9812 8396
rect 6177 8392 9812 8394
rect 6177 8336 6182 8392
rect 6238 8336 9812 8392
rect 6177 8334 9812 8336
rect 6177 8331 6243 8334
rect 9806 8332 9812 8334
rect 9876 8332 9882 8396
rect 12341 8394 12407 8397
rect 13997 8394 14063 8397
rect 14365 8394 14431 8397
rect 12341 8392 14431 8394
rect 12341 8336 12346 8392
rect 12402 8336 14002 8392
rect 14058 8336 14370 8392
rect 14426 8336 14431 8392
rect 12341 8334 14431 8336
rect 12341 8331 12407 8334
rect 13997 8331 14063 8334
rect 14365 8331 14431 8334
rect 15285 8396 15351 8397
rect 15285 8392 15332 8396
rect 15396 8394 15402 8396
rect 17220 8394 17280 8606
rect 17401 8664 19215 8666
rect 17401 8608 17406 8664
rect 17462 8608 19154 8664
rect 19210 8608 19215 8664
rect 17401 8606 19215 8608
rect 17401 8603 17467 8606
rect 19149 8603 19215 8606
rect 19977 8666 20043 8669
rect 23841 8666 23907 8669
rect 19977 8664 23907 8666
rect 19977 8608 19982 8664
rect 20038 8608 23846 8664
rect 23902 8608 23907 8664
rect 19977 8606 23907 8608
rect 19977 8603 20043 8606
rect 23841 8603 23907 8606
rect 18689 8530 18755 8533
rect 33409 8530 33475 8533
rect 18689 8528 33475 8530
rect 18689 8472 18694 8528
rect 18750 8472 33414 8528
rect 33470 8472 33475 8528
rect 18689 8470 33475 8472
rect 18689 8467 18755 8470
rect 33409 8467 33475 8470
rect 20621 8394 20687 8397
rect 15285 8336 15290 8392
rect 15285 8332 15332 8336
rect 15396 8334 15442 8394
rect 16070 8334 16682 8394
rect 17220 8392 20687 8394
rect 17220 8336 20626 8392
rect 20682 8336 20687 8392
rect 17220 8334 20687 8336
rect 15396 8332 15402 8334
rect 15285 8331 15351 8332
rect 7414 8196 7420 8260
rect 7484 8258 7490 8260
rect 9949 8258 10015 8261
rect 7484 8256 10015 8258
rect 7484 8200 9954 8256
rect 10010 8200 10015 8256
rect 7484 8198 10015 8200
rect 7484 8196 7490 8198
rect 9949 8195 10015 8198
rect 13854 8196 13860 8260
rect 13924 8258 13930 8260
rect 14089 8258 14155 8261
rect 15009 8260 15075 8261
rect 15561 8260 15627 8261
rect 14958 8258 14964 8260
rect 13924 8256 14155 8258
rect 13924 8200 14094 8256
rect 14150 8200 14155 8256
rect 13924 8198 14155 8200
rect 14918 8198 14964 8258
rect 15028 8256 15075 8260
rect 15510 8258 15516 8260
rect 15070 8200 15075 8256
rect 13924 8196 13930 8198
rect 14089 8195 14155 8198
rect 14958 8196 14964 8198
rect 15028 8196 15075 8200
rect 15470 8198 15516 8258
rect 15580 8256 15627 8260
rect 16070 8258 16130 8334
rect 15622 8200 15627 8256
rect 15510 8196 15516 8198
rect 15580 8196 15627 8200
rect 15009 8195 15075 8196
rect 15561 8195 15627 8196
rect 15886 8198 16130 8258
rect 16622 8258 16682 8334
rect 20621 8331 20687 8334
rect 25262 8332 25268 8396
rect 25332 8394 25338 8396
rect 25957 8394 26023 8397
rect 25332 8392 26023 8394
rect 25332 8336 25962 8392
rect 26018 8336 26023 8392
rect 25332 8334 26023 8336
rect 25332 8332 25338 8334
rect 25957 8331 26023 8334
rect 19374 8258 19380 8260
rect 16622 8198 19380 8258
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 5390 8060 5396 8124
rect 5460 8122 5466 8124
rect 9949 8122 10015 8125
rect 5460 8120 10015 8122
rect 5460 8064 9954 8120
rect 10010 8064 10015 8120
rect 5460 8062 10015 8064
rect 5460 8060 5466 8062
rect 9949 8059 10015 8062
rect 11462 8060 11468 8124
rect 11532 8122 11538 8124
rect 15886 8122 15946 8198
rect 19374 8196 19380 8198
rect 19444 8196 19450 8260
rect 19517 8258 19583 8261
rect 21449 8258 21515 8261
rect 19517 8256 21515 8258
rect 19517 8200 19522 8256
rect 19578 8200 21454 8256
rect 21510 8200 21515 8256
rect 19517 8198 21515 8200
rect 19517 8195 19583 8198
rect 21449 8195 21515 8198
rect 25037 8258 25103 8261
rect 31886 8258 31892 8260
rect 25037 8256 31892 8258
rect 25037 8200 25042 8256
rect 25098 8200 31892 8256
rect 25037 8198 31892 8200
rect 25037 8195 25103 8198
rect 31886 8196 31892 8198
rect 31956 8196 31962 8260
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 11532 8062 15946 8122
rect 11532 8060 11538 8062
rect 16062 8060 16068 8124
rect 16132 8122 16138 8124
rect 17401 8122 17467 8125
rect 16132 8120 17467 8122
rect 16132 8064 17406 8120
rect 17462 8064 17467 8120
rect 16132 8062 17467 8064
rect 16132 8060 16138 8062
rect 17401 8059 17467 8062
rect 18454 8060 18460 8124
rect 18524 8122 18530 8124
rect 18597 8122 18663 8125
rect 18524 8120 18663 8122
rect 18524 8064 18602 8120
rect 18658 8064 18663 8120
rect 18524 8062 18663 8064
rect 18524 8060 18530 8062
rect 18597 8059 18663 8062
rect 18965 8122 19031 8125
rect 20846 8122 20852 8124
rect 18965 8120 20852 8122
rect 18965 8064 18970 8120
rect 19026 8064 20852 8120
rect 18965 8062 20852 8064
rect 18965 8059 19031 8062
rect 20846 8060 20852 8062
rect 20916 8060 20922 8124
rect 22369 8122 22435 8125
rect 22686 8122 22692 8124
rect 22369 8120 22692 8122
rect 22369 8064 22374 8120
rect 22430 8064 22692 8120
rect 22369 8062 22692 8064
rect 22369 8059 22435 8062
rect 22686 8060 22692 8062
rect 22756 8060 22762 8124
rect 25589 8122 25655 8125
rect 34513 8122 34579 8125
rect 25589 8120 34579 8122
rect 25589 8064 25594 8120
rect 25650 8064 34518 8120
rect 34574 8064 34579 8120
rect 25589 8062 34579 8064
rect 25589 8059 25655 8062
rect 34513 8059 34579 8062
rect 0 7926 3986 7986
rect 0 7896 800 7926
rect 7046 7924 7052 7988
rect 7116 7986 7122 7988
rect 7189 7986 7255 7989
rect 9489 7988 9555 7989
rect 7116 7984 7255 7986
rect 7116 7928 7194 7984
rect 7250 7928 7255 7984
rect 7116 7926 7255 7928
rect 7116 7924 7122 7926
rect 7189 7923 7255 7926
rect 8342 7926 9322 7986
rect 4337 7850 4403 7853
rect 8150 7850 8156 7852
rect 4337 7848 8156 7850
rect 4337 7792 4342 7848
rect 4398 7792 8156 7848
rect 4337 7790 8156 7792
rect 4337 7787 4403 7790
rect 8150 7788 8156 7790
rect 8220 7788 8226 7852
rect 6545 7714 6611 7717
rect 7230 7714 7236 7716
rect 6545 7712 7236 7714
rect 6545 7656 6550 7712
rect 6606 7656 7236 7712
rect 6545 7654 7236 7656
rect 6545 7651 6611 7654
rect 7230 7652 7236 7654
rect 7300 7714 7306 7716
rect 8342 7714 8402 7926
rect 8937 7852 9003 7853
rect 8886 7788 8892 7852
rect 8956 7850 9003 7852
rect 9262 7850 9322 7926
rect 9438 7924 9444 7988
rect 9508 7986 9555 7988
rect 12341 7986 12407 7989
rect 21081 7986 21147 7989
rect 9508 7984 9600 7986
rect 9550 7928 9600 7984
rect 9508 7926 9600 7928
rect 12341 7984 21147 7986
rect 12341 7928 12346 7984
rect 12402 7928 21086 7984
rect 21142 7928 21147 7984
rect 12341 7926 21147 7928
rect 9508 7924 9555 7926
rect 9489 7923 9555 7924
rect 12341 7923 12407 7926
rect 21081 7923 21147 7926
rect 21909 7986 21975 7989
rect 31937 7986 32003 7989
rect 21909 7984 32003 7986
rect 21909 7928 21914 7984
rect 21970 7928 31942 7984
rect 31998 7928 32003 7984
rect 21909 7926 32003 7928
rect 21909 7923 21975 7926
rect 31937 7923 32003 7926
rect 13169 7850 13235 7853
rect 16113 7850 16179 7853
rect 8956 7848 9048 7850
rect 8998 7792 9048 7848
rect 8956 7790 9048 7792
rect 9262 7848 16179 7850
rect 9262 7792 13174 7848
rect 13230 7792 16118 7848
rect 16174 7792 16179 7848
rect 9262 7790 16179 7792
rect 8956 7788 9003 7790
rect 8937 7787 9003 7788
rect 13169 7787 13235 7790
rect 16113 7787 16179 7790
rect 16297 7850 16363 7853
rect 16430 7850 16436 7852
rect 16297 7848 16436 7850
rect 16297 7792 16302 7848
rect 16358 7792 16436 7848
rect 16297 7790 16436 7792
rect 16297 7787 16363 7790
rect 16430 7788 16436 7790
rect 16500 7788 16506 7852
rect 16941 7850 17007 7853
rect 17350 7850 17356 7852
rect 16941 7848 17356 7850
rect 16941 7792 16946 7848
rect 17002 7792 17356 7848
rect 16941 7790 17356 7792
rect 16941 7787 17007 7790
rect 17350 7788 17356 7790
rect 17420 7788 17426 7852
rect 19793 7850 19859 7853
rect 32949 7850 33015 7853
rect 19793 7848 33015 7850
rect 19793 7792 19798 7848
rect 19854 7792 32954 7848
rect 33010 7792 33015 7848
rect 19793 7790 33015 7792
rect 19793 7787 19859 7790
rect 32949 7787 33015 7790
rect 7300 7654 8402 7714
rect 7300 7652 7306 7654
rect 8518 7652 8524 7716
rect 8588 7714 8594 7716
rect 8845 7714 8911 7717
rect 8588 7712 8911 7714
rect 8588 7656 8850 7712
rect 8906 7656 8911 7712
rect 8588 7654 8911 7656
rect 8588 7652 8594 7654
rect 8845 7651 8911 7654
rect 9029 7714 9095 7717
rect 9489 7714 9555 7717
rect 11421 7714 11487 7717
rect 9029 7712 9555 7714
rect 9029 7656 9034 7712
rect 9090 7656 9494 7712
rect 9550 7656 9555 7712
rect 9029 7654 9555 7656
rect 9029 7651 9095 7654
rect 9489 7651 9555 7654
rect 9768 7712 11487 7714
rect 9768 7656 11426 7712
rect 11482 7656 11487 7712
rect 9768 7654 11487 7656
rect 790 7516 796 7580
rect 860 7578 866 7580
rect 860 7518 1042 7578
rect 860 7516 866 7518
rect 982 7442 1042 7518
rect 2446 7516 2452 7580
rect 2516 7578 2522 7580
rect 9581 7578 9647 7581
rect 2516 7576 9647 7578
rect 2516 7520 9586 7576
rect 9642 7520 9647 7576
rect 2516 7518 9647 7520
rect 2516 7516 2522 7518
rect 9581 7515 9647 7518
rect 9768 7442 9828 7654
rect 11421 7651 11487 7654
rect 15285 7714 15351 7717
rect 18965 7714 19031 7717
rect 15285 7712 19031 7714
rect 15285 7656 15290 7712
rect 15346 7656 18970 7712
rect 19026 7656 19031 7712
rect 15285 7654 19031 7656
rect 15285 7651 15351 7654
rect 18965 7651 19031 7654
rect 19977 7714 20043 7717
rect 26550 7714 26556 7716
rect 19977 7712 26556 7714
rect 19977 7656 19982 7712
rect 20038 7656 26556 7712
rect 19977 7654 26556 7656
rect 19977 7651 20043 7654
rect 26550 7652 26556 7654
rect 26620 7652 26626 7716
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 11513 7578 11579 7581
rect 11830 7578 11836 7580
rect 11513 7576 11836 7578
rect 11513 7520 11518 7576
rect 11574 7520 11836 7576
rect 11513 7518 11836 7520
rect 11513 7515 11579 7518
rect 11830 7516 11836 7518
rect 11900 7516 11906 7580
rect 14457 7578 14523 7581
rect 14590 7578 14596 7580
rect 14457 7576 14596 7578
rect 14457 7520 14462 7576
rect 14518 7520 14596 7576
rect 14457 7518 14596 7520
rect 14457 7515 14523 7518
rect 14590 7516 14596 7518
rect 14660 7516 14666 7580
rect 15142 7516 15148 7580
rect 15212 7578 15218 7580
rect 23841 7578 23907 7581
rect 34145 7578 34211 7581
rect 15212 7518 18154 7578
rect 15212 7516 15218 7518
rect 982 7382 9828 7442
rect 9990 7380 9996 7444
rect 10060 7442 10066 7444
rect 10777 7442 10843 7445
rect 17902 7442 17908 7444
rect 10060 7440 10843 7442
rect 10060 7384 10782 7440
rect 10838 7384 10843 7440
rect 10060 7382 10843 7384
rect 10060 7380 10066 7382
rect 10777 7379 10843 7382
rect 11470 7382 17908 7442
rect 0 7306 800 7336
rect 1393 7306 1459 7309
rect 0 7304 1459 7306
rect 0 7248 1398 7304
rect 1454 7248 1459 7304
rect 0 7246 1459 7248
rect 0 7216 800 7246
rect 1393 7243 1459 7246
rect 5073 7306 5139 7309
rect 5206 7306 5212 7308
rect 5073 7304 5212 7306
rect 5073 7248 5078 7304
rect 5134 7248 5212 7304
rect 5073 7246 5212 7248
rect 5073 7243 5139 7246
rect 5206 7244 5212 7246
rect 5276 7244 5282 7308
rect 7649 7306 7715 7309
rect 11470 7306 11530 7382
rect 17902 7380 17908 7382
rect 17972 7380 17978 7444
rect 7649 7304 11530 7306
rect 7649 7248 7654 7304
rect 7710 7248 11530 7304
rect 7649 7246 11530 7248
rect 11605 7306 11671 7309
rect 12566 7306 12572 7308
rect 11605 7304 12572 7306
rect 11605 7248 11610 7304
rect 11666 7248 12572 7304
rect 11605 7246 12572 7248
rect 7649 7243 7715 7246
rect 11605 7243 11671 7246
rect 12566 7244 12572 7246
rect 12636 7244 12642 7308
rect 15009 7306 15075 7309
rect 17309 7306 17375 7309
rect 15009 7304 17375 7306
rect 15009 7248 15014 7304
rect 15070 7248 17314 7304
rect 17370 7248 17375 7304
rect 15009 7246 17375 7248
rect 18094 7306 18154 7518
rect 23841 7576 34211 7578
rect 23841 7520 23846 7576
rect 23902 7520 34150 7576
rect 34206 7520 34211 7576
rect 23841 7518 34211 7520
rect 23841 7515 23907 7518
rect 34145 7515 34211 7518
rect 19425 7442 19491 7445
rect 20110 7442 20116 7444
rect 19425 7440 20116 7442
rect 19425 7384 19430 7440
rect 19486 7384 20116 7440
rect 19425 7382 20116 7384
rect 19425 7379 19491 7382
rect 20110 7380 20116 7382
rect 20180 7380 20186 7444
rect 21265 7442 21331 7445
rect 32857 7442 32923 7445
rect 21265 7440 32923 7442
rect 21265 7384 21270 7440
rect 21326 7384 32862 7440
rect 32918 7384 32923 7440
rect 21265 7382 32923 7384
rect 21265 7379 21331 7382
rect 32857 7379 32923 7382
rect 23105 7306 23171 7309
rect 18094 7304 23171 7306
rect 18094 7248 23110 7304
rect 23166 7248 23171 7304
rect 18094 7246 23171 7248
rect 15009 7243 15075 7246
rect 17309 7243 17375 7246
rect 23105 7243 23171 7246
rect 6637 7170 6703 7173
rect 11145 7170 11211 7173
rect 6637 7168 11211 7170
rect 6637 7112 6642 7168
rect 6698 7112 11150 7168
rect 11206 7112 11211 7168
rect 6637 7110 11211 7112
rect 6637 7107 6703 7110
rect 11145 7107 11211 7110
rect 11278 7108 11284 7172
rect 11348 7170 11354 7172
rect 11421 7170 11487 7173
rect 11348 7168 11487 7170
rect 11348 7112 11426 7168
rect 11482 7112 11487 7168
rect 11348 7110 11487 7112
rect 11348 7108 11354 7110
rect 11421 7107 11487 7110
rect 11605 7170 11671 7173
rect 14089 7170 14155 7173
rect 16297 7170 16363 7173
rect 26141 7170 26207 7173
rect 11605 7168 14155 7170
rect 11605 7112 11610 7168
rect 11666 7112 14094 7168
rect 14150 7112 14155 7168
rect 11605 7110 14155 7112
rect 11605 7107 11671 7110
rect 14089 7107 14155 7110
rect 16254 7168 26207 7170
rect 16254 7112 16302 7168
rect 16358 7112 26146 7168
rect 26202 7112 26207 7168
rect 16254 7110 26207 7112
rect 16254 7107 16363 7110
rect 26141 7107 26207 7110
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 4613 7034 4679 7037
rect 4838 7034 4844 7036
rect 4613 7032 4844 7034
rect 4613 6976 4618 7032
rect 4674 6976 4844 7032
rect 4613 6974 4844 6976
rect 4613 6971 4679 6974
rect 4838 6972 4844 6974
rect 4908 6972 4914 7036
rect 5758 6972 5764 7036
rect 5828 7034 5834 7036
rect 6361 7034 6427 7037
rect 5828 7032 6427 7034
rect 5828 6976 6366 7032
rect 6422 6976 6427 7032
rect 5828 6974 6427 6976
rect 5828 6972 5834 6974
rect 6361 6971 6427 6974
rect 8201 7034 8267 7037
rect 9070 7034 9076 7036
rect 8201 7032 9076 7034
rect 8201 6976 8206 7032
rect 8262 6976 9076 7032
rect 8201 6974 9076 6976
rect 8201 6971 8267 6974
rect 9070 6972 9076 6974
rect 9140 6972 9146 7036
rect 9489 7034 9555 7037
rect 10501 7034 10567 7037
rect 9489 7032 10567 7034
rect 9489 6976 9494 7032
rect 9550 6976 10506 7032
rect 10562 6976 10567 7032
rect 9489 6974 10567 6976
rect 9489 6971 9555 6974
rect 10501 6971 10567 6974
rect 11881 7034 11947 7037
rect 16254 7034 16314 7107
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 16982 7034 16988 7036
rect 11881 7032 16314 7034
rect 11881 6976 11886 7032
rect 11942 6976 16314 7032
rect 11881 6974 16314 6976
rect 16392 6974 16988 7034
rect 11881 6971 11947 6974
rect 4429 6898 4495 6901
rect 4654 6898 4660 6900
rect 4429 6896 4660 6898
rect 4429 6840 4434 6896
rect 4490 6840 4660 6896
rect 4429 6838 4660 6840
rect 4429 6835 4495 6838
rect 4654 6836 4660 6838
rect 4724 6836 4730 6900
rect 5165 6898 5231 6901
rect 5574 6898 5580 6900
rect 5165 6896 5580 6898
rect 5165 6840 5170 6896
rect 5226 6840 5580 6896
rect 5165 6838 5580 6840
rect 5165 6835 5231 6838
rect 5574 6836 5580 6838
rect 5644 6836 5650 6900
rect 9397 6898 9463 6901
rect 10358 6898 10364 6900
rect 9397 6896 10364 6898
rect 9397 6840 9402 6896
rect 9458 6840 10364 6896
rect 9397 6838 10364 6840
rect 9397 6835 9463 6838
rect 10358 6836 10364 6838
rect 10428 6836 10434 6900
rect 13077 6898 13143 6901
rect 15377 6898 15443 6901
rect 13077 6896 15443 6898
rect 13077 6840 13082 6896
rect 13138 6840 15382 6896
rect 15438 6840 15443 6896
rect 13077 6838 15443 6840
rect 13077 6835 13143 6838
rect 15377 6835 15443 6838
rect 0 6762 800 6792
rect 4613 6762 4679 6765
rect 5073 6764 5139 6765
rect 5022 6762 5028 6764
rect 0 6760 4679 6762
rect 0 6704 4618 6760
rect 4674 6704 4679 6760
rect 0 6702 4679 6704
rect 4982 6702 5028 6762
rect 5092 6760 5139 6764
rect 5134 6704 5139 6760
rect 0 6672 800 6702
rect 4613 6699 4679 6702
rect 5022 6700 5028 6702
rect 5092 6700 5139 6704
rect 5073 6699 5139 6700
rect 5349 6762 5415 6765
rect 6126 6762 6132 6764
rect 5349 6760 6132 6762
rect 5349 6704 5354 6760
rect 5410 6704 6132 6760
rect 5349 6702 6132 6704
rect 5349 6699 5415 6702
rect 6126 6700 6132 6702
rect 6196 6700 6202 6764
rect 7465 6762 7531 6765
rect 7598 6762 7604 6764
rect 7465 6760 7604 6762
rect 7465 6704 7470 6760
rect 7526 6704 7604 6760
rect 7465 6702 7604 6704
rect 7465 6699 7531 6702
rect 7598 6700 7604 6702
rect 7668 6700 7674 6764
rect 8293 6762 8359 6765
rect 9581 6762 9647 6765
rect 8293 6760 9647 6762
rect 8293 6704 8298 6760
rect 8354 6704 9586 6760
rect 9642 6704 9647 6760
rect 8293 6702 9647 6704
rect 8293 6699 8359 6702
rect 9581 6699 9647 6702
rect 10501 6762 10567 6765
rect 10726 6762 10732 6764
rect 10501 6760 10732 6762
rect 10501 6704 10506 6760
rect 10562 6704 10732 6760
rect 10501 6702 10732 6704
rect 10501 6699 10567 6702
rect 10726 6700 10732 6702
rect 10796 6700 10802 6764
rect 11881 6762 11947 6765
rect 16392 6762 16452 6974
rect 16982 6972 16988 6974
rect 17052 6972 17058 7036
rect 17902 6972 17908 7036
rect 17972 7034 17978 7036
rect 26182 7034 26188 7036
rect 17972 6974 26188 7034
rect 17972 6972 17978 6974
rect 26182 6972 26188 6974
rect 26252 6972 26258 7036
rect 17125 6898 17191 6901
rect 20621 6898 20687 6901
rect 17125 6896 20687 6898
rect 17125 6840 17130 6896
rect 17186 6840 20626 6896
rect 20682 6840 20687 6896
rect 17125 6838 20687 6840
rect 17125 6835 17191 6838
rect 20621 6835 20687 6838
rect 21909 6898 21975 6901
rect 22277 6898 22343 6901
rect 26877 6898 26943 6901
rect 32438 6898 32444 6900
rect 21909 6896 22343 6898
rect 21909 6840 21914 6896
rect 21970 6840 22282 6896
rect 22338 6840 22343 6896
rect 21909 6838 22343 6840
rect 21909 6835 21975 6838
rect 22277 6835 22343 6838
rect 22694 6838 24042 6898
rect 11881 6760 16452 6762
rect 11881 6704 11886 6760
rect 11942 6704 16452 6760
rect 11881 6702 16452 6704
rect 17217 6760 17283 6765
rect 17217 6704 17222 6760
rect 17278 6704 17283 6760
rect 11881 6699 11947 6702
rect 17217 6699 17283 6704
rect 19701 6762 19767 6765
rect 22694 6762 22754 6838
rect 19701 6760 22754 6762
rect 19701 6704 19706 6760
rect 19762 6704 22754 6760
rect 19701 6702 22754 6704
rect 22921 6762 22987 6765
rect 23841 6762 23907 6765
rect 22921 6760 23907 6762
rect 22921 6704 22926 6760
rect 22982 6704 23846 6760
rect 23902 6704 23907 6760
rect 22921 6702 23907 6704
rect 23982 6762 24042 6838
rect 26877 6896 32444 6898
rect 26877 6840 26882 6896
rect 26938 6840 32444 6896
rect 26877 6838 32444 6840
rect 26877 6835 26943 6838
rect 32438 6836 32444 6838
rect 32508 6836 32514 6900
rect 29085 6762 29151 6765
rect 23982 6760 29151 6762
rect 23982 6704 29090 6760
rect 29146 6704 29151 6760
rect 23982 6702 29151 6704
rect 19701 6699 19767 6702
rect 22921 6699 22987 6702
rect 23841 6699 23907 6702
rect 29085 6699 29151 6702
rect 5809 6626 5875 6629
rect 9949 6626 10015 6629
rect 5809 6624 10015 6626
rect 5809 6568 5814 6624
rect 5870 6568 9954 6624
rect 10010 6568 10015 6624
rect 5809 6566 10015 6568
rect 5809 6563 5875 6566
rect 9949 6563 10015 6566
rect 10593 6626 10659 6629
rect 17220 6626 17280 6699
rect 10593 6624 17280 6626
rect 10593 6568 10598 6624
rect 10654 6568 17280 6624
rect 10593 6566 17280 6568
rect 20069 6626 20135 6629
rect 37457 6626 37523 6629
rect 20069 6624 37523 6626
rect 20069 6568 20074 6624
rect 20130 6568 37462 6624
rect 37518 6568 37523 6624
rect 20069 6566 37523 6568
rect 10593 6563 10659 6566
rect 20069 6563 20135 6566
rect 37457 6563 37523 6566
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 3877 6492 3943 6493
rect 3877 6490 3924 6492
rect 3832 6488 3924 6490
rect 3832 6432 3882 6488
rect 3832 6430 3924 6432
rect 3877 6428 3924 6430
rect 3988 6428 3994 6492
rect 7465 6490 7531 6493
rect 13721 6490 13787 6493
rect 7465 6488 13787 6490
rect 7465 6432 7470 6488
rect 7526 6432 13726 6488
rect 13782 6432 13787 6488
rect 7465 6430 13787 6432
rect 3877 6427 3943 6428
rect 7465 6427 7531 6430
rect 13721 6427 13787 6430
rect 19977 6490 20043 6493
rect 26877 6490 26943 6493
rect 19977 6488 26943 6490
rect 19977 6432 19982 6488
rect 20038 6432 26882 6488
rect 26938 6432 26943 6488
rect 19977 6430 26943 6432
rect 19977 6427 20043 6430
rect 26877 6427 26943 6430
rect 1117 6354 1183 6357
rect 9765 6354 9831 6357
rect 15101 6354 15167 6357
rect 1117 6352 9831 6354
rect 1117 6296 1122 6352
rect 1178 6296 9770 6352
rect 9826 6296 9831 6352
rect 1117 6294 9831 6296
rect 1117 6291 1183 6294
rect 9765 6291 9831 6294
rect 9998 6352 15167 6354
rect 9998 6296 15106 6352
rect 15162 6296 15167 6352
rect 9998 6294 15167 6296
rect 0 6218 800 6248
rect 1485 6218 1551 6221
rect 3325 6218 3391 6221
rect 0 6216 3391 6218
rect 0 6160 1490 6216
rect 1546 6160 3330 6216
rect 3386 6160 3391 6216
rect 0 6158 3391 6160
rect 0 6128 800 6158
rect 1485 6155 1551 6158
rect 3325 6155 3391 6158
rect 8702 6156 8708 6220
rect 8772 6218 8778 6220
rect 9305 6218 9371 6221
rect 8772 6216 9371 6218
rect 8772 6160 9310 6216
rect 9366 6160 9371 6216
rect 8772 6158 9371 6160
rect 8772 6156 8778 6158
rect 9305 6155 9371 6158
rect 9581 6218 9647 6221
rect 9998 6218 10058 6294
rect 15101 6291 15167 6294
rect 15653 6354 15719 6357
rect 20069 6354 20135 6357
rect 15653 6352 20135 6354
rect 15653 6296 15658 6352
rect 15714 6296 20074 6352
rect 20130 6296 20135 6352
rect 15653 6294 20135 6296
rect 15653 6291 15719 6294
rect 20069 6291 20135 6294
rect 20345 6354 20411 6357
rect 20478 6354 20484 6356
rect 20345 6352 20484 6354
rect 20345 6296 20350 6352
rect 20406 6296 20484 6352
rect 20345 6294 20484 6296
rect 20345 6291 20411 6294
rect 20478 6292 20484 6294
rect 20548 6292 20554 6356
rect 23565 6354 23631 6357
rect 33174 6354 33180 6356
rect 23565 6352 33180 6354
rect 23565 6296 23570 6352
rect 23626 6296 33180 6352
rect 23565 6294 33180 6296
rect 23565 6291 23631 6294
rect 33174 6292 33180 6294
rect 33244 6292 33250 6356
rect 9581 6216 10058 6218
rect 9581 6160 9586 6216
rect 9642 6160 10058 6216
rect 9581 6158 10058 6160
rect 10225 6218 10291 6221
rect 14181 6218 14247 6221
rect 10225 6216 14247 6218
rect 10225 6160 10230 6216
rect 10286 6160 14186 6216
rect 14242 6160 14247 6216
rect 10225 6158 14247 6160
rect 9581 6155 9647 6158
rect 10225 6155 10291 6158
rect 14181 6155 14247 6158
rect 15377 6218 15443 6221
rect 32765 6218 32831 6221
rect 15377 6216 32831 6218
rect 15377 6160 15382 6216
rect 15438 6160 32770 6216
rect 32826 6160 32831 6216
rect 15377 6158 32831 6160
rect 15377 6155 15443 6158
rect 32765 6155 32831 6158
rect 8569 6082 8635 6085
rect 10542 6082 10548 6084
rect 8569 6080 10548 6082
rect 8569 6024 8574 6080
rect 8630 6024 10548 6080
rect 8569 6022 10548 6024
rect 8569 6019 8635 6022
rect 10542 6020 10548 6022
rect 10612 6020 10618 6084
rect 11646 6020 11652 6084
rect 11716 6082 11722 6084
rect 13537 6082 13603 6085
rect 11716 6080 13603 6082
rect 11716 6024 13542 6080
rect 13598 6024 13603 6080
rect 11716 6022 13603 6024
rect 11716 6020 11722 6022
rect 13537 6019 13603 6022
rect 16389 6082 16455 6085
rect 25078 6082 25084 6084
rect 16389 6080 25084 6082
rect 16389 6024 16394 6080
rect 16450 6024 25084 6080
rect 16389 6022 25084 6024
rect 16389 6019 16455 6022
rect 25078 6020 25084 6022
rect 25148 6020 25154 6084
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 4981 5946 5047 5949
rect 9397 5948 9463 5949
rect 9397 5946 9444 5948
rect 4981 5944 9444 5946
rect 4981 5888 4986 5944
rect 5042 5888 9402 5944
rect 4981 5886 9444 5888
rect 4981 5883 5047 5886
rect 9397 5884 9444 5886
rect 9508 5884 9514 5948
rect 11053 5946 11119 5949
rect 16757 5946 16823 5949
rect 27153 5948 27219 5949
rect 11053 5944 16823 5946
rect 11053 5888 11058 5944
rect 11114 5888 16762 5944
rect 16818 5888 16823 5944
rect 11053 5886 16823 5888
rect 9397 5883 9463 5884
rect 11053 5883 11119 5886
rect 16757 5883 16823 5886
rect 16982 5884 16988 5948
rect 17052 5946 17058 5948
rect 20294 5946 20300 5948
rect 17052 5886 20300 5946
rect 17052 5884 17058 5886
rect 20294 5884 20300 5886
rect 20364 5884 20370 5948
rect 27102 5884 27108 5948
rect 27172 5946 27219 5948
rect 27797 5946 27863 5949
rect 28022 5946 28028 5948
rect 27172 5944 27264 5946
rect 27214 5888 27264 5944
rect 27172 5886 27264 5888
rect 27797 5944 28028 5946
rect 27797 5888 27802 5944
rect 27858 5888 28028 5944
rect 27797 5886 28028 5888
rect 27172 5884 27219 5886
rect 27153 5883 27219 5884
rect 27797 5883 27863 5886
rect 28022 5884 28028 5886
rect 28092 5884 28098 5948
rect 11329 5810 11395 5813
rect 11462 5810 11468 5812
rect 11329 5808 11468 5810
rect 11329 5752 11334 5808
rect 11390 5752 11468 5808
rect 11329 5750 11468 5752
rect 11329 5747 11395 5750
rect 11462 5748 11468 5750
rect 11532 5748 11538 5812
rect 12249 5810 12315 5813
rect 17166 5810 17172 5812
rect 12249 5808 17172 5810
rect 12249 5752 12254 5808
rect 12310 5752 17172 5808
rect 12249 5750 17172 5752
rect 12249 5747 12315 5750
rect 17166 5748 17172 5750
rect 17236 5748 17242 5812
rect 17585 5810 17651 5813
rect 17585 5808 19994 5810
rect 17585 5752 17590 5808
rect 17646 5752 19994 5808
rect 17585 5750 19994 5752
rect 17585 5747 17651 5750
rect 4654 5612 4660 5676
rect 4724 5674 4730 5676
rect 10225 5674 10291 5677
rect 4724 5672 10291 5674
rect 4724 5616 10230 5672
rect 10286 5616 10291 5672
rect 4724 5614 10291 5616
rect 4724 5612 4730 5614
rect 10225 5611 10291 5614
rect 10593 5674 10659 5677
rect 11789 5676 11855 5677
rect 10726 5674 10732 5676
rect 10593 5672 10732 5674
rect 10593 5616 10598 5672
rect 10654 5616 10732 5672
rect 10593 5614 10732 5616
rect 10593 5611 10659 5614
rect 10726 5612 10732 5614
rect 10796 5612 10802 5676
rect 11789 5674 11836 5676
rect 11744 5672 11836 5674
rect 11744 5616 11794 5672
rect 11744 5614 11836 5616
rect 11789 5612 11836 5614
rect 11900 5612 11906 5676
rect 13854 5612 13860 5676
rect 13924 5674 13930 5676
rect 14365 5674 14431 5677
rect 17585 5676 17651 5677
rect 13924 5672 14431 5674
rect 13924 5616 14370 5672
rect 14426 5616 14431 5672
rect 13924 5614 14431 5616
rect 13924 5612 13930 5614
rect 11789 5611 11855 5612
rect 14365 5611 14431 5614
rect 17534 5612 17540 5676
rect 17604 5674 17651 5676
rect 17604 5672 17696 5674
rect 17646 5616 17696 5672
rect 17604 5614 17696 5616
rect 17604 5612 17651 5614
rect 19374 5612 19380 5676
rect 19444 5674 19450 5676
rect 19701 5674 19767 5677
rect 19444 5672 19767 5674
rect 19444 5616 19706 5672
rect 19762 5616 19767 5672
rect 19444 5614 19767 5616
rect 19934 5674 19994 5750
rect 20478 5748 20484 5812
rect 20548 5810 20554 5812
rect 22921 5810 22987 5813
rect 20548 5808 22987 5810
rect 20548 5752 22926 5808
rect 22982 5752 22987 5808
rect 20548 5750 22987 5752
rect 20548 5748 20554 5750
rect 22921 5747 22987 5750
rect 22185 5676 22251 5677
rect 20662 5674 20668 5676
rect 19934 5614 20668 5674
rect 19444 5612 19450 5614
rect 17585 5611 17651 5612
rect 19701 5611 19767 5614
rect 20662 5612 20668 5614
rect 20732 5612 20738 5676
rect 22134 5674 22140 5676
rect 22094 5614 22140 5674
rect 22204 5672 22251 5676
rect 22246 5616 22251 5672
rect 22134 5612 22140 5614
rect 22204 5612 22251 5616
rect 22185 5611 22251 5612
rect 0 5538 800 5568
rect 3969 5538 4035 5541
rect 0 5536 4035 5538
rect 0 5480 3974 5536
rect 4030 5480 4035 5536
rect 0 5478 4035 5480
rect 0 5448 800 5478
rect 3969 5475 4035 5478
rect 4613 5538 4679 5541
rect 9673 5538 9739 5541
rect 10961 5538 11027 5541
rect 4613 5536 11027 5538
rect 4613 5480 4618 5536
rect 4674 5480 9678 5536
rect 9734 5480 10966 5536
rect 11022 5480 11027 5536
rect 4613 5478 11027 5480
rect 4613 5475 4679 5478
rect 9673 5475 9739 5478
rect 10961 5475 11027 5478
rect 23422 5476 23428 5540
rect 23492 5538 23498 5540
rect 28533 5538 28599 5541
rect 23492 5536 28599 5538
rect 23492 5480 28538 5536
rect 28594 5480 28599 5536
rect 23492 5478 28599 5480
rect 23492 5476 23498 5478
rect 28533 5475 28599 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 4061 5402 4127 5405
rect 18321 5402 18387 5405
rect 19006 5402 19012 5404
rect 4061 5400 17280 5402
rect 4061 5344 4066 5400
rect 4122 5344 17280 5400
rect 4061 5342 17280 5344
rect 4061 5339 4127 5342
rect 657 5266 723 5269
rect 11145 5266 11211 5269
rect 657 5264 11211 5266
rect 657 5208 662 5264
rect 718 5208 11150 5264
rect 11206 5208 11211 5264
rect 657 5206 11211 5208
rect 657 5203 723 5206
rect 11145 5203 11211 5206
rect 12157 5266 12223 5269
rect 13721 5266 13787 5269
rect 12157 5264 13787 5266
rect 12157 5208 12162 5264
rect 12218 5208 13726 5264
rect 13782 5208 13787 5264
rect 12157 5206 13787 5208
rect 17220 5266 17280 5342
rect 18321 5400 19012 5402
rect 18321 5344 18326 5400
rect 18382 5344 19012 5400
rect 18321 5342 19012 5344
rect 18321 5339 18387 5342
rect 19006 5340 19012 5342
rect 19076 5340 19082 5404
rect 21081 5266 21147 5269
rect 17220 5264 21147 5266
rect 17220 5208 21086 5264
rect 21142 5208 21147 5264
rect 17220 5206 21147 5208
rect 12157 5203 12223 5206
rect 13721 5203 13787 5206
rect 21081 5203 21147 5206
rect 22369 5266 22435 5269
rect 33869 5266 33935 5269
rect 22369 5264 33935 5266
rect 22369 5208 22374 5264
rect 22430 5208 33874 5264
rect 33930 5208 33935 5264
rect 22369 5206 33935 5208
rect 22369 5203 22435 5206
rect 33869 5203 33935 5206
rect 5206 5068 5212 5132
rect 5276 5130 5282 5132
rect 10777 5130 10843 5133
rect 5276 5128 10843 5130
rect 5276 5072 10782 5128
rect 10838 5072 10843 5128
rect 5276 5070 10843 5072
rect 5276 5068 5282 5070
rect 10777 5067 10843 5070
rect 16849 5130 16915 5133
rect 22921 5130 22987 5133
rect 16849 5128 22987 5130
rect 16849 5072 16854 5128
rect 16910 5072 22926 5128
rect 22982 5072 22987 5128
rect 16849 5070 22987 5072
rect 16849 5067 16915 5070
rect 22921 5067 22987 5070
rect 27337 5130 27403 5133
rect 34053 5130 34119 5133
rect 27337 5128 34119 5130
rect 27337 5072 27342 5128
rect 27398 5072 34058 5128
rect 34114 5072 34119 5128
rect 27337 5070 34119 5072
rect 27337 5067 27403 5070
rect 34053 5067 34119 5070
rect 0 4994 800 5024
rect 1485 4994 1551 4997
rect 0 4992 1551 4994
rect 0 4936 1490 4992
rect 1546 4936 1551 4992
rect 0 4934 1551 4936
rect 0 4904 800 4934
rect 1485 4931 1551 4934
rect 4889 4994 4955 4997
rect 23657 4994 23723 4997
rect 4889 4992 23723 4994
rect 4889 4936 4894 4992
rect 4950 4936 23662 4992
rect 23718 4936 23723 4992
rect 4889 4934 23723 4936
rect 4889 4931 4955 4934
rect 23657 4931 23723 4934
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 9121 4860 9187 4861
rect 9070 4796 9076 4860
rect 9140 4858 9187 4860
rect 9140 4856 9232 4858
rect 9182 4800 9232 4856
rect 9140 4798 9232 4800
rect 9140 4796 9187 4798
rect 10726 4796 10732 4860
rect 10796 4858 10802 4860
rect 12157 4858 12223 4861
rect 10796 4856 12223 4858
rect 10796 4800 12162 4856
rect 12218 4800 12223 4856
rect 10796 4798 12223 4800
rect 10796 4796 10802 4798
rect 9121 4795 9187 4796
rect 12157 4795 12223 4798
rect 17166 4796 17172 4860
rect 17236 4858 17242 4860
rect 28901 4858 28967 4861
rect 17236 4856 28967 4858
rect 17236 4800 28906 4856
rect 28962 4800 28967 4856
rect 17236 4798 28967 4800
rect 17236 4796 17242 4798
rect 28901 4795 28967 4798
rect 2037 4722 2103 4725
rect 23565 4722 23631 4725
rect 2037 4720 23631 4722
rect 2037 4664 2042 4720
rect 2098 4664 23570 4720
rect 23626 4664 23631 4720
rect 2037 4662 23631 4664
rect 2037 4659 2103 4662
rect 23565 4659 23631 4662
rect 5533 4586 5599 4589
rect 10133 4586 10199 4589
rect 5533 4584 10199 4586
rect 5533 4528 5538 4584
rect 5594 4528 10138 4584
rect 10194 4528 10199 4584
rect 5533 4526 10199 4528
rect 5533 4523 5599 4526
rect 10133 4523 10199 4526
rect 10777 4586 10843 4589
rect 22093 4586 22159 4589
rect 10777 4584 22159 4586
rect 10777 4528 10782 4584
rect 10838 4528 22098 4584
rect 22154 4528 22159 4584
rect 10777 4526 22159 4528
rect 10777 4523 10843 4526
rect 22093 4523 22159 4526
rect 0 4450 800 4480
rect 4061 4450 4127 4453
rect 0 4448 4127 4450
rect 0 4392 4066 4448
rect 4122 4392 4127 4448
rect 0 4390 4127 4392
rect 0 4360 800 4390
rect 4061 4387 4127 4390
rect 8937 4450 9003 4453
rect 13813 4450 13879 4453
rect 8937 4448 13879 4450
rect 8937 4392 8942 4448
rect 8998 4392 13818 4448
rect 13874 4392 13879 4448
rect 8937 4390 13879 4392
rect 8937 4387 9003 4390
rect 13813 4387 13879 4390
rect 14181 4450 14247 4453
rect 17309 4452 17375 4453
rect 16614 4450 16620 4452
rect 14181 4448 16620 4450
rect 14181 4392 14186 4448
rect 14242 4392 16620 4448
rect 14181 4390 16620 4392
rect 14181 4387 14247 4390
rect 16614 4388 16620 4390
rect 16684 4388 16690 4452
rect 17309 4448 17356 4452
rect 17420 4450 17426 4452
rect 20713 4450 20779 4453
rect 22737 4450 22803 4453
rect 17309 4392 17314 4448
rect 17309 4388 17356 4392
rect 17420 4390 17466 4450
rect 20713 4448 22110 4450
rect 20713 4392 20718 4448
rect 20774 4392 22110 4448
rect 20713 4390 22110 4392
rect 17420 4388 17426 4390
rect 17309 4387 17375 4388
rect 20713 4387 20779 4390
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 12433 4314 12499 4317
rect 17677 4314 17743 4317
rect 22050 4314 22110 4390
rect 22737 4448 35910 4450
rect 22737 4392 22742 4448
rect 22798 4392 35910 4448
rect 22737 4390 35910 4392
rect 22737 4387 22803 4390
rect 35850 4314 35910 4390
rect 39849 4314 39915 4317
rect 12433 4312 17743 4314
rect 12433 4256 12438 4312
rect 12494 4256 17682 4312
rect 17738 4256 17743 4312
rect 12433 4254 17743 4256
rect 12433 4251 12499 4254
rect 17677 4251 17743 4254
rect 19980 4254 21788 4314
rect 22050 4254 31770 4314
rect 35850 4312 39915 4314
rect 35850 4256 39854 4312
rect 39910 4256 39915 4312
rect 35850 4254 39915 4256
rect 10501 4178 10567 4181
rect 16982 4178 16988 4180
rect 10501 4176 16988 4178
rect 10501 4120 10506 4176
rect 10562 4120 16988 4176
rect 10501 4118 16988 4120
rect 10501 4115 10567 4118
rect 16982 4116 16988 4118
rect 17052 4116 17058 4180
rect 17309 4178 17375 4181
rect 19980 4178 20040 4254
rect 17309 4176 20040 4178
rect 17309 4120 17314 4176
rect 17370 4120 20040 4176
rect 17309 4118 20040 4120
rect 17309 4115 17375 4118
rect 20662 4116 20668 4180
rect 20732 4178 20738 4180
rect 21541 4178 21607 4181
rect 20732 4176 21607 4178
rect 20732 4120 21546 4176
rect 21602 4120 21607 4176
rect 20732 4118 21607 4120
rect 21728 4178 21788 4254
rect 23105 4178 23171 4181
rect 21728 4176 23171 4178
rect 21728 4120 23110 4176
rect 23166 4120 23171 4176
rect 21728 4118 23171 4120
rect 20732 4116 20738 4118
rect 21541 4115 21607 4118
rect 23105 4115 23171 4118
rect 23422 4116 23428 4180
rect 23492 4178 23498 4180
rect 24025 4178 24091 4181
rect 24945 4180 25011 4181
rect 24894 4178 24900 4180
rect 23492 4176 24091 4178
rect 23492 4120 24030 4176
rect 24086 4120 24091 4176
rect 23492 4118 24091 4120
rect 24854 4118 24900 4178
rect 24964 4176 25011 4180
rect 25006 4120 25011 4176
rect 23492 4116 23498 4118
rect 24025 4115 24091 4118
rect 24894 4116 24900 4118
rect 24964 4116 25011 4120
rect 31710 4178 31770 4254
rect 39849 4251 39915 4254
rect 39389 4178 39455 4181
rect 31710 4176 39455 4178
rect 31710 4120 39394 4176
rect 39450 4120 39455 4176
rect 31710 4118 39455 4120
rect 24945 4115 25011 4116
rect 39389 4115 39455 4118
rect 14181 4044 14247 4045
rect 15377 4044 15443 4045
rect 14181 4040 14228 4044
rect 14292 4042 14298 4044
rect 14181 3984 14186 4040
rect 14181 3980 14228 3984
rect 14292 3982 14338 4042
rect 14292 3980 14298 3982
rect 15326 3980 15332 4044
rect 15396 4042 15443 4044
rect 15837 4042 15903 4045
rect 20437 4042 20503 4045
rect 15396 4040 15488 4042
rect 15438 3984 15488 4040
rect 15396 3982 15488 3984
rect 15837 4040 20503 4042
rect 15837 3984 15842 4040
rect 15898 3984 20442 4040
rect 20498 3984 20503 4040
rect 15837 3982 20503 3984
rect 15396 3980 15443 3982
rect 14181 3979 14247 3980
rect 15377 3979 15443 3980
rect 15837 3979 15903 3982
rect 20437 3979 20503 3982
rect 4705 3906 4771 3909
rect 25129 3906 25195 3909
rect 4705 3904 25195 3906
rect 4705 3848 4710 3904
rect 4766 3848 25134 3904
rect 25190 3848 25195 3904
rect 4705 3846 25195 3848
rect 4705 3843 4771 3846
rect 25129 3843 25195 3846
rect 4208 3840 4528 3841
rect 0 3770 800 3800
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 1393 3770 1459 3773
rect 0 3768 1459 3770
rect 0 3712 1398 3768
rect 1454 3712 1459 3768
rect 0 3710 1459 3712
rect 0 3680 800 3710
rect 1393 3707 1459 3710
rect 9489 3770 9555 3773
rect 15193 3770 15259 3773
rect 29453 3770 29519 3773
rect 9489 3768 15026 3770
rect 9489 3712 9494 3768
rect 9550 3712 15026 3768
rect 9489 3710 15026 3712
rect 9489 3707 9555 3710
rect 3969 3634 4035 3637
rect 13854 3634 13860 3636
rect 3969 3632 13860 3634
rect 3969 3576 3974 3632
rect 4030 3576 13860 3632
rect 3969 3574 13860 3576
rect 3969 3571 4035 3574
rect 13854 3572 13860 3574
rect 13924 3572 13930 3636
rect 14966 3634 15026 3710
rect 15193 3768 29519 3770
rect 15193 3712 15198 3768
rect 15254 3712 29458 3768
rect 29514 3712 29519 3768
rect 15193 3710 29519 3712
rect 15193 3707 15259 3710
rect 29453 3707 29519 3710
rect 15837 3634 15903 3637
rect 14966 3632 15903 3634
rect 14966 3576 15842 3632
rect 15898 3576 15903 3632
rect 14966 3574 15903 3576
rect 15837 3571 15903 3574
rect 18689 3634 18755 3637
rect 31937 3634 32003 3637
rect 18689 3632 32003 3634
rect 18689 3576 18694 3632
rect 18750 3576 31942 3632
rect 31998 3576 32003 3632
rect 18689 3574 32003 3576
rect 18689 3571 18755 3574
rect 31937 3571 32003 3574
rect 4613 3498 4679 3501
rect 15929 3498 15995 3501
rect 4613 3496 15995 3498
rect 4613 3440 4618 3496
rect 4674 3440 15934 3496
rect 15990 3440 15995 3496
rect 4613 3438 15995 3440
rect 4613 3435 4679 3438
rect 15929 3435 15995 3438
rect 19333 3498 19399 3501
rect 24577 3498 24643 3501
rect 19333 3496 24643 3498
rect 19333 3440 19338 3496
rect 19394 3440 24582 3496
rect 24638 3440 24643 3496
rect 19333 3438 24643 3440
rect 19333 3435 19399 3438
rect 24577 3435 24643 3438
rect 6729 3362 6795 3365
rect 11789 3362 11855 3365
rect 6729 3360 11855 3362
rect 6729 3304 6734 3360
rect 6790 3304 11794 3360
rect 11850 3304 11855 3360
rect 6729 3302 11855 3304
rect 6729 3299 6795 3302
rect 11789 3299 11855 3302
rect 14774 3300 14780 3364
rect 14844 3362 14850 3364
rect 15101 3362 15167 3365
rect 16573 3362 16639 3365
rect 14844 3360 16639 3362
rect 14844 3304 15106 3360
rect 15162 3304 16578 3360
rect 16634 3304 16639 3360
rect 14844 3302 16639 3304
rect 14844 3300 14850 3302
rect 15101 3299 15167 3302
rect 16573 3299 16639 3302
rect 19568 3296 19888 3297
rect 0 3226 800 3256
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 3877 3226 3943 3229
rect 0 3224 3943 3226
rect 0 3168 3882 3224
rect 3938 3168 3943 3224
rect 0 3166 3943 3168
rect 0 3136 800 3166
rect 3877 3163 3943 3166
rect 4061 3226 4127 3229
rect 9990 3226 9996 3228
rect 4061 3224 9996 3226
rect 4061 3168 4066 3224
rect 4122 3168 9996 3224
rect 4061 3166 9996 3168
rect 4061 3163 4127 3166
rect 9990 3164 9996 3166
rect 10060 3164 10066 3228
rect 11145 3226 11211 3229
rect 12934 3226 12940 3228
rect 11145 3224 12940 3226
rect 11145 3168 11150 3224
rect 11206 3168 12940 3224
rect 11145 3166 12940 3168
rect 11145 3163 11211 3166
rect 12934 3164 12940 3166
rect 13004 3164 13010 3228
rect 13670 3164 13676 3228
rect 13740 3226 13746 3228
rect 14365 3226 14431 3229
rect 17033 3226 17099 3229
rect 13740 3224 14431 3226
rect 13740 3168 14370 3224
rect 14426 3168 14431 3224
rect 13740 3166 14431 3168
rect 13740 3164 13746 3166
rect 14365 3163 14431 3166
rect 16438 3224 17099 3226
rect 16438 3168 17038 3224
rect 17094 3168 17099 3224
rect 16438 3166 17099 3168
rect 3417 3090 3483 3093
rect 16438 3090 16498 3166
rect 17033 3163 17099 3166
rect 23054 3164 23060 3228
rect 23124 3226 23130 3228
rect 40217 3226 40283 3229
rect 23124 3224 40283 3226
rect 23124 3168 40222 3224
rect 40278 3168 40283 3224
rect 23124 3166 40283 3168
rect 23124 3164 23130 3166
rect 40217 3163 40283 3166
rect 3417 3088 16498 3090
rect 3417 3032 3422 3088
rect 3478 3032 16498 3088
rect 3417 3030 16498 3032
rect 3417 3027 3483 3030
rect 16614 3028 16620 3092
rect 16684 3090 16690 3092
rect 34513 3090 34579 3093
rect 16684 3088 34579 3090
rect 16684 3032 34518 3088
rect 34574 3032 34579 3088
rect 16684 3030 34579 3032
rect 16684 3028 16690 3030
rect 34513 3027 34579 3030
rect 13721 2954 13787 2957
rect 33225 2954 33291 2957
rect 13721 2952 33291 2954
rect 13721 2896 13726 2952
rect 13782 2896 33230 2952
rect 33286 2896 33291 2952
rect 13721 2894 33291 2896
rect 13721 2891 13787 2894
rect 33225 2891 33291 2894
rect 5165 2818 5231 2821
rect 21909 2818 21975 2821
rect 5165 2816 21975 2818
rect 5165 2760 5170 2816
rect 5226 2760 21914 2816
rect 21970 2760 21975 2816
rect 5165 2758 21975 2760
rect 5165 2755 5231 2758
rect 21909 2755 21975 2758
rect 4208 2752 4528 2753
rect 0 2682 800 2712
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 3049 2682 3115 2685
rect 0 2680 3115 2682
rect 0 2624 3054 2680
rect 3110 2624 3115 2680
rect 0 2622 3115 2624
rect 0 2592 800 2622
rect 3049 2619 3115 2622
rect 7005 2682 7071 2685
rect 15510 2682 15516 2684
rect 7005 2680 15516 2682
rect 7005 2624 7010 2680
rect 7066 2624 15516 2680
rect 7005 2622 15516 2624
rect 7005 2619 7071 2622
rect 15510 2620 15516 2622
rect 15580 2620 15586 2684
rect 17769 2682 17835 2685
rect 17902 2682 17908 2684
rect 17769 2680 17908 2682
rect 17769 2624 17774 2680
rect 17830 2624 17908 2680
rect 17769 2622 17908 2624
rect 17769 2619 17835 2622
rect 17902 2620 17908 2622
rect 17972 2620 17978 2684
rect 18229 2682 18295 2685
rect 18229 2680 31034 2682
rect 18229 2624 18234 2680
rect 18290 2624 31034 2680
rect 18229 2622 31034 2624
rect 18229 2619 18295 2622
rect 933 2546 999 2549
rect 9765 2546 9831 2549
rect 933 2544 9831 2546
rect 933 2488 938 2544
rect 994 2488 9770 2544
rect 9826 2488 9831 2544
rect 933 2486 9831 2488
rect 933 2483 999 2486
rect 9765 2483 9831 2486
rect 10133 2546 10199 2549
rect 19374 2546 19380 2548
rect 10133 2544 19380 2546
rect 10133 2488 10138 2544
rect 10194 2488 19380 2544
rect 10133 2486 19380 2488
rect 10133 2483 10199 2486
rect 19374 2484 19380 2486
rect 19444 2484 19450 2548
rect 24894 2546 24900 2548
rect 19566 2486 24900 2546
rect 15837 2410 15903 2413
rect 19190 2410 19196 2412
rect 15837 2408 19196 2410
rect 15837 2352 15842 2408
rect 15898 2352 19196 2408
rect 15837 2350 19196 2352
rect 15837 2347 15903 2350
rect 19190 2348 19196 2350
rect 19260 2348 19266 2412
rect 19566 2410 19626 2486
rect 24894 2484 24900 2486
rect 24964 2484 24970 2548
rect 25957 2546 26023 2549
rect 28574 2546 28580 2548
rect 25957 2544 28580 2546
rect 25957 2488 25962 2544
rect 26018 2488 28580 2544
rect 25957 2486 28580 2488
rect 25957 2483 26023 2486
rect 28574 2484 28580 2486
rect 28644 2484 28650 2548
rect 30974 2546 31034 2622
rect 35065 2546 35131 2549
rect 30974 2544 35131 2546
rect 30974 2488 35070 2544
rect 35126 2488 35131 2544
rect 30974 2486 35131 2488
rect 35065 2483 35131 2486
rect 19382 2350 19626 2410
rect 9581 2274 9647 2277
rect 19382 2274 19442 2350
rect 23606 2348 23612 2412
rect 23676 2410 23682 2412
rect 42885 2410 42951 2413
rect 23676 2408 42951 2410
rect 23676 2352 42890 2408
rect 42946 2352 42951 2408
rect 23676 2350 42951 2352
rect 23676 2348 23682 2350
rect 42885 2347 42951 2350
rect 9581 2272 19442 2274
rect 9581 2216 9586 2272
rect 9642 2216 19442 2272
rect 9581 2214 19442 2216
rect 9581 2211 9647 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 3049 2138 3115 2141
rect 15142 2138 15148 2140
rect 3049 2136 15148 2138
rect 3049 2080 3054 2136
rect 3110 2080 15148 2136
rect 3049 2078 15148 2080
rect 3049 2075 3115 2078
rect 15142 2076 15148 2078
rect 15212 2076 15218 2140
rect 0 2002 800 2032
rect 4061 2002 4127 2005
rect 0 2000 4127 2002
rect 0 1944 4066 2000
rect 4122 1944 4127 2000
rect 0 1942 4127 1944
rect 0 1912 800 1942
rect 4061 1939 4127 1942
rect 18505 2002 18571 2005
rect 27981 2002 28047 2005
rect 18505 2000 28047 2002
rect 18505 1944 18510 2000
rect 18566 1944 27986 2000
rect 28042 1944 28047 2000
rect 18505 1942 28047 1944
rect 18505 1939 18571 1942
rect 27981 1939 28047 1942
rect 6545 1866 6611 1869
rect 26417 1866 26483 1869
rect 6545 1864 26483 1866
rect 6545 1808 6550 1864
rect 6606 1808 26422 1864
rect 26478 1808 26483 1864
rect 6545 1806 26483 1808
rect 6545 1803 6611 1806
rect 26417 1803 26483 1806
rect 17861 1730 17927 1733
rect 6870 1728 17927 1730
rect 6870 1672 17866 1728
rect 17922 1672 17927 1728
rect 6870 1670 17927 1672
rect 2957 1594 3023 1597
rect 6870 1594 6930 1670
rect 17861 1667 17927 1670
rect 2957 1592 6930 1594
rect 2957 1536 2962 1592
rect 3018 1536 6930 1592
rect 2957 1534 6930 1536
rect 12433 1594 12499 1597
rect 17309 1594 17375 1597
rect 12433 1592 17375 1594
rect 12433 1536 12438 1592
rect 12494 1536 17314 1592
rect 17370 1536 17375 1592
rect 12433 1534 17375 1536
rect 2957 1531 3023 1534
rect 12433 1531 12499 1534
rect 17309 1531 17375 1534
rect 17534 1532 17540 1596
rect 17604 1594 17610 1596
rect 20713 1594 20779 1597
rect 17604 1592 20779 1594
rect 17604 1536 20718 1592
rect 20774 1536 20779 1592
rect 17604 1534 20779 1536
rect 17604 1532 17610 1534
rect 20713 1531 20779 1534
rect 0 1458 800 1488
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1368 800 1398
rect 2865 1395 2931 1398
rect 17350 1396 17356 1460
rect 17420 1458 17426 1460
rect 30373 1458 30439 1461
rect 17420 1456 30439 1458
rect 17420 1400 30378 1456
rect 30434 1400 30439 1456
rect 17420 1398 30439 1400
rect 17420 1396 17426 1398
rect 30373 1395 30439 1398
rect 3325 1322 3391 1325
rect 20478 1322 20484 1324
rect 3325 1320 20484 1322
rect 3325 1264 3330 1320
rect 3386 1264 20484 1320
rect 3325 1262 20484 1264
rect 3325 1259 3391 1262
rect 20478 1260 20484 1262
rect 20548 1260 20554 1324
rect 22185 1322 22251 1325
rect 23790 1322 23796 1324
rect 22185 1320 23796 1322
rect 22185 1264 22190 1320
rect 22246 1264 23796 1320
rect 22185 1262 23796 1264
rect 22185 1259 22251 1262
rect 23790 1260 23796 1262
rect 23860 1260 23866 1324
rect 4613 1186 4679 1189
rect 24393 1186 24459 1189
rect 4613 1184 24459 1186
rect 4613 1128 4618 1184
rect 4674 1128 24398 1184
rect 24454 1128 24459 1184
rect 4613 1126 24459 1128
rect 4613 1123 4679 1126
rect 24393 1123 24459 1126
rect 20161 1050 20227 1053
rect 27102 1050 27108 1052
rect 20161 1048 27108 1050
rect 20161 992 20166 1048
rect 20222 992 27108 1048
rect 20161 990 27108 992
rect 20161 987 20227 990
rect 27102 988 27108 990
rect 27172 988 27178 1052
rect 0 914 800 944
rect 2773 914 2839 917
rect 0 912 2839 914
rect 0 856 2778 912
rect 2834 856 2839 912
rect 0 854 2839 856
rect 0 824 800 854
rect 2773 851 2839 854
rect 3141 914 3207 917
rect 25262 914 25268 916
rect 3141 912 25268 914
rect 3141 856 3146 912
rect 3202 856 25268 912
rect 3141 854 25268 856
rect 3141 851 3207 854
rect 25262 852 25268 854
rect 25332 852 25338 916
rect 11605 778 11671 781
rect 23422 778 23428 780
rect 11605 776 23428 778
rect 11605 720 11610 776
rect 11666 720 23428 776
rect 11605 718 23428 720
rect 11605 715 11671 718
rect 23422 716 23428 718
rect 23492 716 23498 780
rect 21766 580 21772 644
rect 21836 642 21842 644
rect 40125 642 40191 645
rect 21836 640 40191 642
rect 21836 584 40130 640
rect 40186 584 40191 640
rect 21836 582 40191 584
rect 21836 580 21842 582
rect 40125 579 40191 582
rect 0 370 800 400
rect 933 370 999 373
rect 0 368 999 370
rect 0 312 938 368
rect 994 312 999 368
rect 0 310 999 312
rect 0 280 800 310
rect 933 307 999 310
rect 6177 234 6243 237
rect 20662 234 20668 236
rect 6177 232 20668 234
rect 6177 176 6182 232
rect 6238 176 20668 232
rect 6177 174 20668 176
rect 6177 171 6243 174
rect 20662 172 20668 174
rect 20732 172 20738 236
rect 4245 98 4311 101
rect 22134 98 22140 100
rect 4245 96 22140 98
rect 4245 40 4250 96
rect 4306 40 22140 96
rect 4245 38 22140 40
rect 4245 35 4311 38
rect 22134 36 22140 38
rect 22204 36 22210 100
<< via3 >>
rect 27476 37844 27540 37908
rect 22508 37572 22572 37636
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 18092 37436 18156 37500
rect 28396 37436 28460 37500
rect 15884 37300 15948 37364
rect 23980 37300 24044 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 16988 36544 17052 36548
rect 16988 36488 17038 36544
rect 17038 36488 17052 36544
rect 16988 36484 17052 36488
rect 17724 36544 17788 36548
rect 17724 36488 17774 36544
rect 17774 36488 17788 36544
rect 17724 36484 17788 36488
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19380 36076 19444 36140
rect 5580 35940 5644 36004
rect 14412 36000 14476 36004
rect 14412 35944 14426 36000
rect 14426 35944 14476 36000
rect 14412 35940 14476 35944
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4660 34640 4724 34644
rect 4660 34584 4710 34640
rect 4710 34584 4724 34640
rect 4660 34580 4724 34584
rect 14964 34580 15028 34644
rect 17540 34580 17604 34644
rect 26740 34580 26804 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 22692 32404 22756 32468
rect 26004 32404 26068 32468
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 17908 30500 17972 30564
rect 27292 30500 27356 30564
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 14780 30364 14844 30428
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 25452 29276 25516 29340
rect 5948 29140 6012 29204
rect 33180 29140 33244 29204
rect 3556 29004 3620 29068
rect 3924 29064 3988 29068
rect 3924 29008 3938 29064
rect 3938 29008 3988 29064
rect 3924 29004 3988 29008
rect 5212 29004 5276 29068
rect 15148 28868 15212 28932
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 18460 28460 18524 28524
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 1348 28052 1412 28116
rect 23428 28052 23492 28116
rect 6868 27916 6932 27980
rect 20484 27916 20548 27980
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 7604 27100 7668 27164
rect 16068 26964 16132 27028
rect 7052 26828 7116 26892
rect 7236 26692 7300 26756
rect 24900 26828 24964 26892
rect 11836 26692 11900 26756
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 13308 26556 13372 26620
rect 9444 26480 9508 26484
rect 9444 26424 9494 26480
rect 9494 26424 9508 26480
rect 9444 26420 9508 26424
rect 12756 26420 12820 26484
rect 14044 26420 14108 26484
rect 1164 26284 1228 26348
rect 21036 26284 21100 26348
rect 6868 26208 6932 26212
rect 6868 26152 6918 26208
rect 6918 26152 6932 26208
rect 6868 26148 6932 26152
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 11100 25604 11164 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 9076 25468 9140 25532
rect 29316 25468 29380 25532
rect 10364 25060 10428 25124
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 8708 24848 8772 24852
rect 8708 24792 8722 24848
rect 8722 24792 8772 24848
rect 8708 24788 8772 24792
rect 15700 24848 15764 24852
rect 15700 24792 15750 24848
rect 15750 24792 15764 24848
rect 15700 24788 15764 24792
rect 20668 24788 20732 24852
rect 32260 24788 32324 24852
rect 1716 24516 1780 24580
rect 5396 24516 5460 24580
rect 20852 24516 20916 24580
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 10916 24380 10980 24444
rect 21772 24380 21836 24444
rect 20300 24108 20364 24172
rect 2268 23972 2332 24036
rect 10180 24032 10244 24036
rect 10180 23976 10194 24032
rect 10194 23976 10244 24032
rect 10180 23972 10244 23976
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 2820 23896 2884 23900
rect 2820 23840 2870 23896
rect 2870 23840 2884 23896
rect 2820 23836 2884 23840
rect 5764 23836 5828 23900
rect 10548 23836 10612 23900
rect 17172 23700 17236 23764
rect 6684 23624 6748 23628
rect 6684 23568 6698 23624
rect 6698 23568 6748 23624
rect 6684 23564 6748 23568
rect 7788 23564 7852 23628
rect 25084 23564 25148 23628
rect 1532 23428 1596 23492
rect 4844 23428 4908 23492
rect 7604 23428 7668 23492
rect 9260 23428 9324 23492
rect 12572 23428 12636 23492
rect 16804 23488 16868 23492
rect 16804 23432 16854 23488
rect 16854 23432 16868 23488
rect 16804 23428 16868 23432
rect 17540 23428 17604 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 3924 23156 3988 23220
rect 18092 23216 18156 23220
rect 18092 23160 18106 23216
rect 18106 23160 18156 23216
rect 18092 23156 18156 23160
rect 10732 23020 10796 23084
rect 13124 23020 13188 23084
rect 3924 22944 3988 22948
rect 3924 22888 3974 22944
rect 3974 22888 3988 22944
rect 3924 22884 3988 22888
rect 9444 22884 9508 22948
rect 10364 22884 10428 22948
rect 13492 22884 13556 22948
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 7420 22748 7484 22812
rect 15884 22808 15948 22812
rect 15884 22752 15898 22808
rect 15898 22752 15948 22808
rect 15884 22748 15948 22752
rect 9076 22612 9140 22676
rect 11100 22612 11164 22676
rect 11284 22672 11348 22676
rect 11284 22616 11334 22672
rect 11334 22616 11348 22672
rect 11284 22612 11348 22616
rect 10364 22536 10428 22540
rect 10364 22480 10378 22536
rect 10378 22480 10428 22536
rect 10364 22476 10428 22480
rect 8892 22340 8956 22404
rect 9260 22340 9324 22404
rect 9444 22340 9508 22404
rect 17356 22476 17420 22540
rect 18276 22340 18340 22404
rect 30420 22340 30484 22404
rect 30788 22340 30852 22404
rect 31524 22340 31588 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 3556 21856 3620 21860
rect 3556 21800 3606 21856
rect 3606 21800 3620 21856
rect 3556 21796 3620 21800
rect 6500 21796 6564 21860
rect 7052 21932 7116 21996
rect 10180 21932 10244 21996
rect 10732 21932 10796 21996
rect 27660 22068 27724 22132
rect 16988 21932 17052 21996
rect 17724 21796 17788 21860
rect 18644 21796 18708 21860
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 13308 21660 13372 21724
rect 5028 21524 5092 21588
rect 14780 21524 14844 21588
rect 31892 21524 31956 21588
rect 15884 21388 15948 21452
rect 16252 21388 16316 21452
rect 12756 21252 12820 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 4660 20980 4724 21044
rect 12020 20980 12084 21044
rect 24532 21388 24596 21452
rect 27108 21116 27172 21180
rect 15884 20980 15948 21044
rect 16252 20980 16316 21044
rect 24164 20980 24228 21044
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 3924 20844 3988 20908
rect 12756 20844 12820 20908
rect 980 20708 1044 20772
rect 12204 20708 12268 20772
rect 16988 20844 17052 20908
rect 21404 20844 21468 20908
rect 16252 20708 16316 20772
rect 18460 20768 18524 20772
rect 18460 20712 18474 20768
rect 18474 20712 18524 20768
rect 18460 20708 18524 20712
rect 20300 20708 20364 20772
rect 22140 20768 22204 20772
rect 22140 20712 22190 20768
rect 22190 20712 22204 20768
rect 22140 20708 22204 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 5580 20632 5644 20636
rect 5580 20576 5594 20632
rect 5594 20576 5644 20632
rect 5580 20572 5644 20576
rect 10180 20572 10244 20636
rect 14412 20632 14476 20636
rect 14412 20576 14426 20632
rect 14426 20576 14476 20632
rect 14412 20572 14476 20576
rect 14964 20632 15028 20636
rect 14964 20576 15014 20632
rect 15014 20576 15028 20632
rect 14964 20572 15028 20576
rect 15148 20632 15212 20636
rect 15148 20576 15198 20632
rect 15198 20576 15212 20632
rect 15148 20572 15212 20576
rect 16436 20572 16500 20636
rect 22692 20632 22756 20636
rect 22692 20576 22706 20632
rect 22706 20576 22756 20632
rect 22692 20572 22756 20576
rect 28396 20632 28460 20636
rect 28396 20576 28410 20632
rect 28410 20576 28460 20632
rect 28396 20572 28460 20576
rect 8708 20436 8772 20500
rect 4844 20300 4908 20364
rect 6684 20360 6748 20364
rect 6684 20304 6698 20360
rect 6698 20304 6748 20360
rect 6684 20300 6748 20304
rect 9260 20300 9324 20364
rect 12572 20300 12636 20364
rect 11836 20164 11900 20228
rect 29132 20224 29196 20228
rect 29132 20168 29146 20224
rect 29146 20168 29196 20224
rect 29132 20164 29196 20168
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 3740 20088 3804 20092
rect 3740 20032 3754 20088
rect 3754 20032 3804 20088
rect 3740 20028 3804 20032
rect 13308 20028 13372 20092
rect 25268 19892 25332 19956
rect 5580 19620 5644 19684
rect 13676 19756 13740 19820
rect 14964 19756 15028 19820
rect 25820 19756 25884 19820
rect 32076 19756 32140 19820
rect 8156 19620 8220 19684
rect 16620 19620 16684 19684
rect 22324 19620 22388 19684
rect 28948 19620 29012 19684
rect 31340 19680 31404 19684
rect 31340 19624 31390 19680
rect 31390 19624 31404 19680
rect 31340 19620 31404 19624
rect 33916 19620 33980 19684
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 3188 19348 3252 19412
rect 5028 19348 5092 19412
rect 5764 19348 5828 19412
rect 6684 19348 6748 19412
rect 9628 19484 9692 19548
rect 10364 19544 10428 19548
rect 10364 19488 10378 19544
rect 10378 19488 10428 19544
rect 10364 19484 10428 19488
rect 21220 19544 21284 19548
rect 21220 19488 21270 19544
rect 21270 19488 21284 19544
rect 13860 19348 13924 19412
rect 14596 19348 14660 19412
rect 21220 19484 21284 19488
rect 21956 19544 22020 19548
rect 21956 19488 22006 19544
rect 22006 19488 22020 19544
rect 21956 19484 22020 19488
rect 30236 19544 30300 19548
rect 30236 19488 30250 19544
rect 30250 19488 30300 19544
rect 30236 19484 30300 19488
rect 25084 19348 25148 19412
rect 26004 19408 26068 19412
rect 26004 19352 26054 19408
rect 26054 19352 26068 19408
rect 26004 19348 26068 19352
rect 27844 19348 27908 19412
rect 28580 19348 28644 19412
rect 2268 19212 2332 19276
rect 16068 19212 16132 19276
rect 16804 19212 16868 19276
rect 18092 19272 18156 19276
rect 18092 19216 18142 19272
rect 18142 19216 18156 19272
rect 18092 19212 18156 19216
rect 19380 19212 19444 19276
rect 22140 19212 22204 19276
rect 25452 19272 25516 19276
rect 25452 19216 25502 19272
rect 25502 19216 25516 19272
rect 25452 19212 25516 19216
rect 27292 19272 27356 19276
rect 27292 19216 27306 19272
rect 27306 19216 27356 19272
rect 27292 19212 27356 19216
rect 11652 19076 11716 19140
rect 19380 19076 19444 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 12572 18940 12636 19004
rect 2820 18804 2884 18868
rect 22508 18940 22572 19004
rect 20668 18804 20732 18868
rect 3004 18668 3068 18732
rect 5948 18668 6012 18732
rect 20300 18668 20364 18732
rect 28028 18668 28092 18732
rect 11284 18532 11348 18596
rect 15516 18532 15580 18596
rect 16804 18532 16868 18596
rect 26556 18592 26620 18596
rect 26556 18536 26606 18592
rect 26606 18536 26620 18592
rect 26556 18532 26620 18536
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 5212 18396 5276 18460
rect 24900 18396 24964 18460
rect 24900 18260 24964 18324
rect 26740 18260 26804 18324
rect 32260 18260 32324 18324
rect 3556 17988 3620 18052
rect 12940 17988 13004 18052
rect 18092 18048 18156 18052
rect 18092 17992 18142 18048
rect 18142 17992 18156 18048
rect 18092 17988 18156 17992
rect 20116 17988 20180 18052
rect 22692 17988 22756 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 15516 17852 15580 17916
rect 17172 17912 17236 17916
rect 17172 17856 17186 17912
rect 17186 17856 17236 17912
rect 17172 17852 17236 17856
rect 17908 17852 17972 17916
rect 8708 17580 8772 17644
rect 17724 17580 17788 17644
rect 20300 17852 20364 17916
rect 20668 17852 20732 17916
rect 21036 17852 21100 17916
rect 22508 17852 22572 17916
rect 32444 18124 32508 18188
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 27660 17852 27724 17916
rect 19012 17640 19076 17644
rect 19012 17584 19026 17640
rect 19026 17584 19076 17640
rect 19012 17580 19076 17584
rect 20668 17580 20732 17644
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 19196 17308 19260 17372
rect 27660 17308 27724 17372
rect 1164 17036 1228 17100
rect 12388 16900 12452 16964
rect 18460 16900 18524 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 10548 16764 10612 16828
rect 19380 16764 19444 16828
rect 20300 16764 20364 16828
rect 22140 16824 22204 16828
rect 22140 16768 22154 16824
rect 22154 16768 22204 16824
rect 22140 16764 22204 16768
rect 7604 16688 7668 16692
rect 7604 16632 7618 16688
rect 7618 16632 7668 16688
rect 7604 16628 7668 16632
rect 13676 16628 13740 16692
rect 19012 16688 19076 16692
rect 19012 16632 19062 16688
rect 19062 16632 19076 16688
rect 19012 16628 19076 16632
rect 19380 16628 19444 16692
rect 20852 16628 20916 16692
rect 5580 16492 5644 16556
rect 6500 16492 6564 16556
rect 7236 16552 7300 16556
rect 7236 16496 7250 16552
rect 7250 16496 7300 16552
rect 7236 16492 7300 16496
rect 9628 16492 9692 16556
rect 18828 16492 18892 16556
rect 21220 16492 21284 16556
rect 10916 16356 10980 16420
rect 19012 16356 19076 16420
rect 20852 16356 20916 16420
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 1716 16280 1780 16284
rect 1716 16224 1730 16280
rect 1730 16224 1780 16280
rect 1716 16220 1780 16224
rect 18092 16220 18156 16284
rect 1532 16008 1596 16012
rect 1532 15952 1582 16008
rect 1582 15952 1596 16008
rect 1532 15948 1596 15952
rect 6684 16008 6748 16012
rect 6684 15952 6734 16008
rect 6734 15952 6748 16008
rect 6684 15948 6748 15952
rect 16068 15812 16132 15876
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 8156 15676 8220 15740
rect 18092 15676 18156 15740
rect 30420 15676 30484 15740
rect 2268 15404 2332 15468
rect 16804 15268 16868 15332
rect 20300 15268 20364 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 5028 15132 5092 15196
rect 17908 15132 17972 15196
rect 19196 15132 19260 15196
rect 20852 15192 20916 15196
rect 20852 15136 20866 15192
rect 20866 15136 20916 15192
rect 20852 15132 20916 15136
rect 21588 15132 21652 15196
rect 24900 15132 24964 15196
rect 25084 15132 25148 15196
rect 27844 15132 27908 15196
rect 23980 14920 24044 14924
rect 23980 14864 24030 14920
rect 24030 14864 24044 14920
rect 23980 14860 24044 14864
rect 30236 14860 30300 14924
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 17172 14724 17236 14788
rect 19380 14724 19444 14788
rect 20300 14724 20364 14788
rect 13492 14588 13556 14652
rect 18460 14588 18524 14652
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 27476 14648 27540 14652
rect 27476 14592 27490 14648
rect 27490 14592 27540 14648
rect 13124 14512 13188 14516
rect 13124 14456 13138 14512
rect 13138 14456 13188 14512
rect 13124 14452 13188 14456
rect 27476 14588 27540 14592
rect 1164 14316 1228 14380
rect 5396 14316 5460 14380
rect 28948 14316 29012 14380
rect 3924 14240 3988 14244
rect 3924 14184 3938 14240
rect 3938 14184 3988 14240
rect 3924 14180 3988 14184
rect 28948 14180 29012 14244
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 12204 14044 12268 14108
rect 15700 14104 15764 14108
rect 15700 14048 15750 14104
rect 15750 14048 15764 14104
rect 15700 14044 15764 14048
rect 16988 14044 17052 14108
rect 18644 14044 18708 14108
rect 23428 14104 23492 14108
rect 23428 14048 23442 14104
rect 23442 14048 23492 14104
rect 23428 14044 23492 14048
rect 29316 14104 29380 14108
rect 29316 14048 29330 14104
rect 29330 14048 29380 14104
rect 29316 14044 29380 14048
rect 2636 13908 2700 13972
rect 7236 13908 7300 13972
rect 12756 13772 12820 13836
rect 13676 13772 13740 13836
rect 14228 13908 14292 13972
rect 20852 13908 20916 13972
rect 23428 13908 23492 13972
rect 1900 13636 1964 13700
rect 5948 13636 6012 13700
rect 8340 13636 8404 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 5396 13500 5460 13564
rect 8156 13500 8220 13564
rect 9444 13500 9508 13564
rect 22140 13560 22204 13564
rect 22140 13504 22154 13560
rect 22154 13504 22204 13560
rect 22140 13500 22204 13504
rect 7420 13364 7484 13428
rect 22508 13424 22572 13428
rect 22508 13368 22558 13424
rect 22558 13368 22572 13424
rect 22508 13364 22572 13368
rect 3004 13228 3068 13292
rect 5212 13228 5276 13292
rect 7604 13228 7668 13292
rect 18460 13228 18524 13292
rect 3556 13152 3620 13156
rect 3556 13096 3570 13152
rect 3570 13096 3620 13152
rect 3556 13092 3620 13096
rect 9260 13092 9324 13156
rect 10364 13092 10428 13156
rect 18460 13092 18524 13156
rect 19380 13092 19444 13156
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 10548 13016 10612 13020
rect 10548 12960 10598 13016
rect 10598 12960 10612 13016
rect 10548 12956 10612 12960
rect 16804 12820 16868 12884
rect 18092 12820 18156 12884
rect 4660 12548 4724 12612
rect 5580 12548 5644 12612
rect 13860 12548 13924 12612
rect 22324 12548 22388 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 5396 12412 5460 12476
rect 6684 12412 6748 12476
rect 18644 12412 18708 12476
rect 31708 12472 31772 12476
rect 31708 12416 31722 12472
rect 31722 12416 31772 12472
rect 31708 12412 31772 12416
rect 16988 12276 17052 12340
rect 17908 12276 17972 12340
rect 20668 12276 20732 12340
rect 17540 12140 17604 12204
rect 20484 12140 20548 12204
rect 27660 12276 27724 12340
rect 31708 12336 31772 12340
rect 31708 12280 31722 12336
rect 31722 12280 31772 12336
rect 31708 12276 31772 12280
rect 1348 12004 1412 12068
rect 10548 12004 10612 12068
rect 18644 12064 18708 12068
rect 18644 12008 18658 12064
rect 18658 12008 18708 12064
rect 18644 12004 18708 12008
rect 20668 12004 20732 12068
rect 21036 12004 21100 12068
rect 5580 11868 5644 11932
rect 7788 11868 7852 11932
rect 19012 11868 19076 11932
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 20484 11868 20548 11932
rect 13860 11732 13924 11796
rect 20300 11732 20364 11796
rect 4844 11460 4908 11524
rect 29132 11732 29196 11796
rect 31340 11596 31404 11660
rect 23612 11520 23676 11524
rect 23612 11464 23626 11520
rect 23626 11464 23676 11520
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 23612 11460 23676 11464
rect 23796 11460 23860 11524
rect 33916 11460 33980 11524
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4844 11384 4908 11388
rect 4844 11328 4894 11384
rect 4894 11328 4908 11384
rect 4844 11324 4908 11328
rect 5028 11052 5092 11116
rect 11284 11324 11348 11388
rect 10180 11188 10244 11252
rect 17356 11324 17420 11388
rect 12940 11248 13004 11252
rect 12940 11192 12954 11248
rect 12954 11192 13004 11248
rect 12940 11188 13004 11192
rect 14228 11188 14292 11252
rect 14412 11188 14476 11252
rect 21404 11324 21468 11388
rect 24532 11324 24596 11388
rect 2636 10916 2700 10980
rect 4660 10780 4724 10844
rect 6132 10780 6196 10844
rect 6500 10840 6564 10844
rect 6500 10784 6514 10840
rect 6514 10784 6564 10840
rect 6500 10780 6564 10784
rect 7052 10780 7116 10844
rect 17540 10780 17604 10844
rect 19196 10840 19260 10844
rect 19196 10784 19246 10840
rect 19246 10784 19260 10840
rect 19196 10780 19260 10784
rect 11100 10644 11164 10708
rect 30788 11052 30852 11116
rect 23428 10916 23492 10980
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 7972 10508 8036 10572
rect 12940 10508 13004 10572
rect 14044 10568 14108 10572
rect 14044 10512 14058 10568
rect 14058 10512 14108 10568
rect 14044 10508 14108 10512
rect 14780 10508 14844 10572
rect 21588 10372 21652 10436
rect 21772 10372 21836 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 7420 10236 7484 10300
rect 9260 10236 9324 10300
rect 9812 10236 9876 10300
rect 2452 10100 2516 10164
rect 4660 9964 4724 10028
rect 8156 9964 8220 10028
rect 17356 10236 17420 10300
rect 20484 10236 20548 10300
rect 31524 10236 31588 10300
rect 12388 9964 12452 10028
rect 28948 10160 29012 10164
rect 28948 10104 28998 10160
rect 28998 10104 29012 10160
rect 28948 10100 29012 10104
rect 5212 9828 5276 9892
rect 8708 9828 8772 9892
rect 9444 9828 9508 9892
rect 3188 9692 3252 9756
rect 3556 9752 3620 9756
rect 3556 9696 3606 9752
rect 3606 9696 3620 9752
rect 3556 9692 3620 9696
rect 13308 9828 13372 9892
rect 14412 9888 14476 9892
rect 14412 9832 14462 9888
rect 14462 9832 14476 9888
rect 14412 9828 14476 9832
rect 19012 9828 19076 9892
rect 20300 9828 20364 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 1164 9556 1228 9620
rect 7788 9556 7852 9620
rect 12020 9616 12084 9620
rect 20484 9692 20548 9756
rect 21036 9692 21100 9756
rect 12020 9560 12034 9616
rect 12034 9560 12084 9616
rect 12020 9556 12084 9560
rect 17172 9556 17236 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 5948 9148 6012 9212
rect 1348 8936 1412 8940
rect 1348 8880 1398 8936
rect 1398 8880 1412 8936
rect 1348 8876 1412 8880
rect 980 8740 1044 8804
rect 5580 8876 5644 8940
rect 7972 9148 8036 9212
rect 16620 9420 16684 9484
rect 18828 9556 18892 9620
rect 19012 9556 19076 9620
rect 23428 9556 23492 9620
rect 24164 9616 24228 9620
rect 24164 9560 24214 9616
rect 24214 9560 24228 9616
rect 24164 9556 24228 9560
rect 25820 9556 25884 9620
rect 18276 9420 18340 9484
rect 18644 9480 18708 9484
rect 18644 9424 18658 9480
rect 18658 9424 18708 9480
rect 18644 9420 18708 9424
rect 8708 9208 8772 9212
rect 17724 9284 17788 9348
rect 23060 9284 23124 9348
rect 32076 9420 32140 9484
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 8708 9152 8722 9208
rect 8722 9152 8772 9208
rect 8708 9148 8772 9152
rect 12756 9148 12820 9212
rect 16252 9148 16316 9212
rect 17540 9148 17604 9212
rect 18092 9208 18156 9212
rect 18092 9152 18106 9208
rect 18106 9152 18156 9208
rect 18092 9148 18156 9152
rect 25268 9148 25332 9212
rect 26188 9148 26252 9212
rect 10548 9012 10612 9076
rect 7420 8936 7484 8940
rect 7420 8880 7434 8936
rect 7434 8880 7484 8936
rect 7420 8876 7484 8880
rect 16804 8876 16868 8940
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 3004 8604 3068 8668
rect 1900 8332 1964 8396
rect 2268 8196 2332 8260
rect 2636 8120 2700 8124
rect 2636 8064 2686 8120
rect 2686 8064 2700 8120
rect 2636 8060 2700 8064
rect 6684 8468 6748 8532
rect 9812 8332 9876 8396
rect 15332 8392 15396 8396
rect 15332 8336 15346 8392
rect 15346 8336 15396 8392
rect 15332 8332 15396 8336
rect 7420 8196 7484 8260
rect 13860 8196 13924 8260
rect 14964 8256 15028 8260
rect 14964 8200 15014 8256
rect 15014 8200 15028 8256
rect 14964 8196 15028 8200
rect 15516 8256 15580 8260
rect 15516 8200 15566 8256
rect 15566 8200 15580 8256
rect 15516 8196 15580 8200
rect 25268 8332 25332 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 5396 8060 5460 8124
rect 11468 8060 11532 8124
rect 19380 8196 19444 8260
rect 31892 8196 31956 8260
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 16068 8060 16132 8124
rect 18460 8060 18524 8124
rect 20852 8060 20916 8124
rect 22692 8060 22756 8124
rect 7052 7924 7116 7988
rect 8156 7788 8220 7852
rect 7236 7652 7300 7716
rect 8892 7848 8956 7852
rect 9444 7984 9508 7988
rect 9444 7928 9494 7984
rect 9494 7928 9508 7984
rect 9444 7924 9508 7928
rect 8892 7792 8942 7848
rect 8942 7792 8956 7848
rect 8892 7788 8956 7792
rect 16436 7788 16500 7852
rect 17356 7788 17420 7852
rect 8524 7652 8588 7716
rect 796 7516 860 7580
rect 2452 7516 2516 7580
rect 26556 7652 26620 7716
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 11836 7516 11900 7580
rect 14596 7516 14660 7580
rect 15148 7516 15212 7580
rect 9996 7380 10060 7444
rect 5212 7244 5276 7308
rect 17908 7380 17972 7444
rect 12572 7244 12636 7308
rect 20116 7380 20180 7444
rect 11284 7108 11348 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4844 6972 4908 7036
rect 5764 6972 5828 7036
rect 9076 6972 9140 7036
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4660 6836 4724 6900
rect 5580 6836 5644 6900
rect 10364 6836 10428 6900
rect 5028 6760 5092 6764
rect 5028 6704 5078 6760
rect 5078 6704 5092 6760
rect 5028 6700 5092 6704
rect 6132 6700 6196 6764
rect 7604 6700 7668 6764
rect 10732 6700 10796 6764
rect 16988 6972 17052 7036
rect 17908 6972 17972 7036
rect 26188 6972 26252 7036
rect 32444 6836 32508 6900
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 3924 6488 3988 6492
rect 3924 6432 3938 6488
rect 3938 6432 3988 6488
rect 3924 6428 3988 6432
rect 8708 6156 8772 6220
rect 20484 6292 20548 6356
rect 33180 6292 33244 6356
rect 10548 6020 10612 6084
rect 11652 6020 11716 6084
rect 25084 6020 25148 6084
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 9444 5944 9508 5948
rect 9444 5888 9458 5944
rect 9458 5888 9508 5944
rect 9444 5884 9508 5888
rect 16988 5884 17052 5948
rect 20300 5884 20364 5948
rect 27108 5944 27172 5948
rect 27108 5888 27158 5944
rect 27158 5888 27172 5944
rect 27108 5884 27172 5888
rect 28028 5884 28092 5948
rect 11468 5748 11532 5812
rect 17172 5748 17236 5812
rect 4660 5612 4724 5676
rect 10732 5612 10796 5676
rect 11836 5672 11900 5676
rect 11836 5616 11850 5672
rect 11850 5616 11900 5672
rect 11836 5612 11900 5616
rect 13860 5612 13924 5676
rect 17540 5672 17604 5676
rect 17540 5616 17590 5672
rect 17590 5616 17604 5672
rect 17540 5612 17604 5616
rect 19380 5612 19444 5676
rect 20484 5748 20548 5812
rect 20668 5612 20732 5676
rect 22140 5672 22204 5676
rect 22140 5616 22190 5672
rect 22190 5616 22204 5672
rect 22140 5612 22204 5616
rect 23428 5476 23492 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 19012 5340 19076 5404
rect 5212 5068 5276 5132
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 9076 4856 9140 4860
rect 9076 4800 9126 4856
rect 9126 4800 9140 4856
rect 9076 4796 9140 4800
rect 10732 4796 10796 4860
rect 17172 4796 17236 4860
rect 16620 4388 16684 4452
rect 17356 4448 17420 4452
rect 17356 4392 17370 4448
rect 17370 4392 17420 4448
rect 17356 4388 17420 4392
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 16988 4116 17052 4180
rect 20668 4116 20732 4180
rect 23428 4116 23492 4180
rect 24900 4176 24964 4180
rect 24900 4120 24950 4176
rect 24950 4120 24964 4176
rect 24900 4116 24964 4120
rect 14228 4040 14292 4044
rect 14228 3984 14242 4040
rect 14242 3984 14292 4040
rect 14228 3980 14292 3984
rect 15332 4040 15396 4044
rect 15332 3984 15382 4040
rect 15382 3984 15396 4040
rect 15332 3980 15396 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 13860 3572 13924 3636
rect 14780 3300 14844 3364
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 9996 3164 10060 3228
rect 12940 3164 13004 3228
rect 13676 3164 13740 3228
rect 23060 3164 23124 3228
rect 16620 3028 16684 3092
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 15516 2620 15580 2684
rect 17908 2620 17972 2684
rect 19380 2484 19444 2548
rect 19196 2348 19260 2412
rect 24900 2484 24964 2548
rect 28580 2484 28644 2548
rect 23612 2348 23676 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 15148 2076 15212 2140
rect 17540 1532 17604 1596
rect 17356 1396 17420 1460
rect 20484 1260 20548 1324
rect 23796 1260 23860 1324
rect 27108 988 27172 1052
rect 25268 852 25332 916
rect 23428 716 23492 780
rect 21772 580 21836 644
rect 20668 172 20732 236
rect 22140 36 22204 100
<< metal4 >>
rect 27475 37908 27541 37909
rect 27475 37844 27476 37908
rect 27540 37844 27541 37908
rect 27475 37843 27541 37844
rect 22507 37636 22573 37637
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 18091 37500 18157 37501
rect 18091 37436 18092 37500
rect 18156 37436 18157 37500
rect 18091 37435 18157 37436
rect 15883 37364 15949 37365
rect 15883 37300 15884 37364
rect 15948 37300 15949 37364
rect 15883 37299 15949 37300
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 5579 36004 5645 36005
rect 5579 35940 5580 36004
rect 5644 35940 5645 36004
rect 5579 35939 5645 35940
rect 14411 36004 14477 36005
rect 14411 35940 14412 36004
rect 14476 35940 14477 36004
rect 14411 35939 14477 35940
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4659 34644 4725 34645
rect 4659 34580 4660 34644
rect 4724 34580 4725 34644
rect 4659 34579 4725 34580
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 3555 29068 3621 29069
rect 3555 29004 3556 29068
rect 3620 29004 3621 29068
rect 3555 29003 3621 29004
rect 3923 29068 3989 29069
rect 3923 29004 3924 29068
rect 3988 29004 3989 29068
rect 3923 29003 3989 29004
rect 1347 28116 1413 28117
rect 1347 28052 1348 28116
rect 1412 28052 1413 28116
rect 1347 28051 1413 28052
rect 1163 26348 1229 26349
rect 1163 26284 1164 26348
rect 1228 26284 1229 26348
rect 1163 26283 1229 26284
rect 979 20772 1045 20773
rect 979 20770 980 20772
rect 798 20710 980 20770
rect 798 7581 858 20710
rect 979 20708 980 20710
rect 1044 20708 1045 20772
rect 979 20707 1045 20708
rect 1166 17101 1226 26283
rect 1163 17100 1229 17101
rect 1163 17036 1164 17100
rect 1228 17036 1229 17100
rect 1163 17035 1229 17036
rect 1350 16590 1410 28051
rect 1715 24580 1781 24581
rect 1715 24516 1716 24580
rect 1780 24516 1781 24580
rect 1715 24515 1781 24516
rect 1531 23492 1597 23493
rect 1531 23428 1532 23492
rect 1596 23428 1597 23492
rect 1531 23427 1597 23428
rect 982 16530 1410 16590
rect 982 8805 1042 16530
rect 1534 16013 1594 23427
rect 1718 16285 1778 24515
rect 2267 24036 2333 24037
rect 2267 23972 2268 24036
rect 2332 23972 2333 24036
rect 2267 23971 2333 23972
rect 2270 19277 2330 23971
rect 2819 23900 2885 23901
rect 2819 23836 2820 23900
rect 2884 23836 2885 23900
rect 2819 23835 2885 23836
rect 2267 19276 2333 19277
rect 2267 19212 2268 19276
rect 2332 19212 2333 19276
rect 2267 19211 2333 19212
rect 2822 18869 2882 23835
rect 3558 22110 3618 29003
rect 3926 23221 3986 29003
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 3923 23220 3989 23221
rect 3923 23156 3924 23220
rect 3988 23156 3989 23220
rect 3923 23155 3989 23156
rect 3923 22948 3989 22949
rect 3923 22884 3924 22948
rect 3988 22884 3989 22948
rect 3923 22883 3989 22884
rect 3558 22050 3802 22110
rect 3555 21860 3621 21861
rect 3555 21796 3556 21860
rect 3620 21796 3621 21860
rect 3555 21795 3621 21796
rect 3187 19412 3253 19413
rect 3187 19348 3188 19412
rect 3252 19348 3253 19412
rect 3187 19347 3253 19348
rect 2819 18868 2885 18869
rect 2819 18804 2820 18868
rect 2884 18804 2885 18868
rect 2819 18803 2885 18804
rect 3003 18732 3069 18733
rect 3003 18668 3004 18732
rect 3068 18668 3069 18732
rect 3003 18667 3069 18668
rect 1715 16284 1781 16285
rect 1715 16220 1716 16284
rect 1780 16220 1781 16284
rect 1715 16219 1781 16220
rect 1531 16012 1597 16013
rect 1531 15948 1532 16012
rect 1596 15948 1597 16012
rect 1531 15947 1597 15948
rect 2267 15468 2333 15469
rect 2267 15404 2268 15468
rect 2332 15404 2333 15468
rect 2267 15403 2333 15404
rect 1163 14380 1229 14381
rect 1163 14316 1164 14380
rect 1228 14316 1229 14380
rect 1163 14315 1229 14316
rect 1166 9621 1226 14315
rect 1899 13700 1965 13701
rect 1899 13636 1900 13700
rect 1964 13636 1965 13700
rect 1899 13635 1965 13636
rect 1347 12068 1413 12069
rect 1347 12004 1348 12068
rect 1412 12004 1413 12068
rect 1347 12003 1413 12004
rect 1163 9620 1229 9621
rect 1163 9556 1164 9620
rect 1228 9556 1229 9620
rect 1163 9555 1229 9556
rect 1350 8941 1410 12003
rect 1347 8940 1413 8941
rect 1347 8876 1348 8940
rect 1412 8876 1413 8940
rect 1347 8875 1413 8876
rect 979 8804 1045 8805
rect 979 8740 980 8804
rect 1044 8740 1045 8804
rect 979 8739 1045 8740
rect 1902 8397 1962 13635
rect 1899 8396 1965 8397
rect 1899 8332 1900 8396
rect 1964 8332 1965 8396
rect 1899 8331 1965 8332
rect 2270 8261 2330 15403
rect 2635 13972 2701 13973
rect 2635 13908 2636 13972
rect 2700 13908 2701 13972
rect 2635 13907 2701 13908
rect 2638 10981 2698 13907
rect 3006 13293 3066 18667
rect 3003 13292 3069 13293
rect 3003 13228 3004 13292
rect 3068 13228 3069 13292
rect 3003 13227 3069 13228
rect 2635 10980 2701 10981
rect 2635 10916 2636 10980
rect 2700 10916 2701 10980
rect 2635 10915 2701 10916
rect 2451 10164 2517 10165
rect 2451 10100 2452 10164
rect 2516 10100 2517 10164
rect 2451 10099 2517 10100
rect 2267 8260 2333 8261
rect 2267 8196 2268 8260
rect 2332 8196 2333 8260
rect 2267 8195 2333 8196
rect 2454 7581 2514 10099
rect 2638 8125 2698 10915
rect 3006 8669 3066 13227
rect 3190 9757 3250 19347
rect 3558 18053 3618 21795
rect 3742 20093 3802 22050
rect 3926 20909 3986 22883
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 3923 20908 3989 20909
rect 3923 20844 3924 20908
rect 3988 20844 3989 20908
rect 3923 20843 3989 20844
rect 4208 20160 4528 21184
rect 4662 21045 4722 34579
rect 5211 29068 5277 29069
rect 5211 29004 5212 29068
rect 5276 29004 5277 29068
rect 5211 29003 5277 29004
rect 4843 23492 4909 23493
rect 4843 23428 4844 23492
rect 4908 23428 4909 23492
rect 4843 23427 4909 23428
rect 4659 21044 4725 21045
rect 4659 20980 4660 21044
rect 4724 20980 4725 21044
rect 4659 20979 4725 20980
rect 4846 20365 4906 23427
rect 5027 21588 5093 21589
rect 5027 21524 5028 21588
rect 5092 21524 5093 21588
rect 5027 21523 5093 21524
rect 4843 20364 4909 20365
rect 4843 20300 4844 20364
rect 4908 20300 4909 20364
rect 4843 20299 4909 20300
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 3739 20092 3805 20093
rect 3739 20028 3740 20092
rect 3804 20028 3805 20092
rect 3739 20027 3805 20028
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 3555 18052 3621 18053
rect 3555 17988 3556 18052
rect 3620 17988 3621 18052
rect 3555 17987 3621 17988
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 3923 14244 3989 14245
rect 3923 14180 3924 14244
rect 3988 14180 3989 14244
rect 3923 14179 3989 14180
rect 3555 13156 3621 13157
rect 3555 13092 3556 13156
rect 3620 13092 3621 13156
rect 3555 13091 3621 13092
rect 3558 9757 3618 13091
rect 3187 9756 3253 9757
rect 3187 9692 3188 9756
rect 3252 9692 3253 9756
rect 3187 9691 3253 9692
rect 3555 9756 3621 9757
rect 3555 9692 3556 9756
rect 3620 9692 3621 9756
rect 3555 9691 3621 9692
rect 3003 8668 3069 8669
rect 3003 8604 3004 8668
rect 3068 8604 3069 8668
rect 3003 8603 3069 8604
rect 2635 8124 2701 8125
rect 2635 8060 2636 8124
rect 2700 8060 2701 8124
rect 2635 8059 2701 8060
rect 795 7580 861 7581
rect 795 7516 796 7580
rect 860 7516 861 7580
rect 795 7515 861 7516
rect 2451 7580 2517 7581
rect 2451 7516 2452 7580
rect 2516 7516 2517 7580
rect 2451 7515 2517 7516
rect 3926 6493 3986 14179
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4659 12612 4725 12613
rect 4659 12548 4660 12612
rect 4724 12548 4725 12612
rect 4659 12547 4725 12548
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4662 10845 4722 12547
rect 4846 11525 4906 20299
rect 5030 19413 5090 21523
rect 5027 19412 5093 19413
rect 5027 19348 5028 19412
rect 5092 19348 5093 19412
rect 5027 19347 5093 19348
rect 5030 15197 5090 19347
rect 5214 18461 5274 29003
rect 5395 24580 5461 24581
rect 5395 24516 5396 24580
rect 5460 24516 5461 24580
rect 5395 24515 5461 24516
rect 5211 18460 5277 18461
rect 5211 18396 5212 18460
rect 5276 18396 5277 18460
rect 5211 18395 5277 18396
rect 5027 15196 5093 15197
rect 5027 15132 5028 15196
rect 5092 15132 5093 15196
rect 5027 15131 5093 15132
rect 5398 14381 5458 24515
rect 5582 20637 5642 35939
rect 5947 29204 6013 29205
rect 5947 29140 5948 29204
rect 6012 29140 6013 29204
rect 5947 29139 6013 29140
rect 5763 23900 5829 23901
rect 5763 23836 5764 23900
rect 5828 23836 5829 23900
rect 5763 23835 5829 23836
rect 5579 20636 5645 20637
rect 5579 20572 5580 20636
rect 5644 20572 5645 20636
rect 5579 20571 5645 20572
rect 5579 19684 5645 19685
rect 5579 19620 5580 19684
rect 5644 19620 5645 19684
rect 5579 19619 5645 19620
rect 5582 16557 5642 19619
rect 5766 19413 5826 23835
rect 5763 19412 5829 19413
rect 5763 19348 5764 19412
rect 5828 19348 5829 19412
rect 5763 19347 5829 19348
rect 5950 18733 6010 29139
rect 6867 27980 6933 27981
rect 6867 27916 6868 27980
rect 6932 27916 6933 27980
rect 6867 27915 6933 27916
rect 6870 26213 6930 27915
rect 7603 27164 7669 27165
rect 7603 27100 7604 27164
rect 7668 27100 7669 27164
rect 7603 27099 7669 27100
rect 7051 26892 7117 26893
rect 7051 26828 7052 26892
rect 7116 26828 7117 26892
rect 7051 26827 7117 26828
rect 6867 26212 6933 26213
rect 6867 26210 6868 26212
rect 6502 26150 6868 26210
rect 6502 21861 6562 26150
rect 6867 26148 6868 26150
rect 6932 26148 6933 26212
rect 6867 26147 6933 26148
rect 6683 23628 6749 23629
rect 6683 23564 6684 23628
rect 6748 23564 6749 23628
rect 6683 23563 6749 23564
rect 6499 21860 6565 21861
rect 6499 21796 6500 21860
rect 6564 21796 6565 21860
rect 6499 21795 6565 21796
rect 6686 20365 6746 23563
rect 7054 21997 7114 26827
rect 7235 26756 7301 26757
rect 7235 26692 7236 26756
rect 7300 26692 7301 26756
rect 7235 26691 7301 26692
rect 7051 21996 7117 21997
rect 7051 21932 7052 21996
rect 7116 21932 7117 21996
rect 7051 21931 7117 21932
rect 6683 20364 6749 20365
rect 6683 20300 6684 20364
rect 6748 20300 6749 20364
rect 6683 20299 6749 20300
rect 6683 19412 6749 19413
rect 6683 19348 6684 19412
rect 6748 19348 6749 19412
rect 6683 19347 6749 19348
rect 5947 18732 6013 18733
rect 5947 18668 5948 18732
rect 6012 18668 6013 18732
rect 5947 18667 6013 18668
rect 5579 16556 5645 16557
rect 5579 16492 5580 16556
rect 5644 16492 5645 16556
rect 5579 16491 5645 16492
rect 6499 16556 6565 16557
rect 6499 16492 6500 16556
rect 6564 16492 6565 16556
rect 6499 16491 6565 16492
rect 5395 14380 5461 14381
rect 5395 14316 5396 14380
rect 5460 14316 5461 14380
rect 5395 14315 5461 14316
rect 5398 13565 5458 14315
rect 5947 13700 6013 13701
rect 5947 13636 5948 13700
rect 6012 13636 6013 13700
rect 5947 13635 6013 13636
rect 5395 13564 5461 13565
rect 5395 13500 5396 13564
rect 5460 13500 5461 13564
rect 5395 13499 5461 13500
rect 5211 13292 5277 13293
rect 5211 13228 5212 13292
rect 5276 13228 5277 13292
rect 5211 13227 5277 13228
rect 4843 11524 4909 11525
rect 4843 11460 4844 11524
rect 4908 11460 4909 11524
rect 4843 11459 4909 11460
rect 4843 11388 4909 11389
rect 4843 11324 4844 11388
rect 4908 11324 4909 11388
rect 4843 11323 4909 11324
rect 4659 10844 4725 10845
rect 4659 10780 4660 10844
rect 4724 10780 4725 10844
rect 4659 10779 4725 10780
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4659 10028 4725 10029
rect 4659 9964 4660 10028
rect 4724 9964 4725 10028
rect 4659 9963 4725 9964
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 3923 6492 3989 6493
rect 3923 6428 3924 6492
rect 3988 6428 3989 6492
rect 3923 6427 3989 6428
rect 4208 6016 4528 7040
rect 4662 6901 4722 9963
rect 4846 7037 4906 11323
rect 5027 11116 5093 11117
rect 5027 11052 5028 11116
rect 5092 11052 5093 11116
rect 5027 11051 5093 11052
rect 4843 7036 4909 7037
rect 4843 6972 4844 7036
rect 4908 6972 4909 7036
rect 4843 6971 4909 6972
rect 4659 6900 4725 6901
rect 4659 6836 4660 6900
rect 4724 6836 4725 6900
rect 4659 6835 4725 6836
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4662 5677 4722 6835
rect 5030 6765 5090 11051
rect 5214 9893 5274 13227
rect 5579 12612 5645 12613
rect 5579 12548 5580 12612
rect 5644 12548 5645 12612
rect 5579 12547 5645 12548
rect 5395 12476 5461 12477
rect 5395 12412 5396 12476
rect 5460 12412 5461 12476
rect 5395 12411 5461 12412
rect 5211 9892 5277 9893
rect 5211 9828 5212 9892
rect 5276 9828 5277 9892
rect 5211 9827 5277 9828
rect 5214 7309 5274 9827
rect 5398 8125 5458 12411
rect 5582 11933 5642 12547
rect 5579 11932 5645 11933
rect 5579 11868 5580 11932
rect 5644 11930 5645 11932
rect 5644 11870 5826 11930
rect 5644 11868 5645 11870
rect 5579 11867 5645 11868
rect 5579 8940 5645 8941
rect 5579 8876 5580 8940
rect 5644 8876 5645 8940
rect 5579 8875 5645 8876
rect 5395 8124 5461 8125
rect 5395 8060 5396 8124
rect 5460 8060 5461 8124
rect 5395 8059 5461 8060
rect 5211 7308 5277 7309
rect 5211 7244 5212 7308
rect 5276 7244 5277 7308
rect 5211 7243 5277 7244
rect 5027 6764 5093 6765
rect 5027 6700 5028 6764
rect 5092 6700 5093 6764
rect 5027 6699 5093 6700
rect 4659 5676 4725 5677
rect 4659 5612 4660 5676
rect 4724 5612 4725 5676
rect 4659 5611 4725 5612
rect 5214 5133 5274 7243
rect 5582 6901 5642 8875
rect 5766 7037 5826 11870
rect 5950 9213 6010 13635
rect 6502 10845 6562 16491
rect 6686 16013 6746 19347
rect 7238 16557 7298 26691
rect 7606 23493 7666 27099
rect 11835 26756 11901 26757
rect 11835 26692 11836 26756
rect 11900 26692 11901 26756
rect 11835 26691 11901 26692
rect 9443 26484 9509 26485
rect 9443 26420 9444 26484
rect 9508 26420 9509 26484
rect 9443 26419 9509 26420
rect 9075 25532 9141 25533
rect 9075 25468 9076 25532
rect 9140 25468 9141 25532
rect 9075 25467 9141 25468
rect 8707 24852 8773 24853
rect 8707 24788 8708 24852
rect 8772 24788 8773 24852
rect 8707 24787 8773 24788
rect 7787 23628 7853 23629
rect 7787 23564 7788 23628
rect 7852 23564 7853 23628
rect 7787 23563 7853 23564
rect 7603 23492 7669 23493
rect 7603 23428 7604 23492
rect 7668 23428 7669 23492
rect 7603 23427 7669 23428
rect 7419 22812 7485 22813
rect 7419 22748 7420 22812
rect 7484 22748 7485 22812
rect 7419 22747 7485 22748
rect 7235 16556 7301 16557
rect 7235 16492 7236 16556
rect 7300 16492 7301 16556
rect 7235 16491 7301 16492
rect 6683 16012 6749 16013
rect 6683 15948 6684 16012
rect 6748 15948 6749 16012
rect 6683 15947 6749 15948
rect 7235 13972 7301 13973
rect 7235 13908 7236 13972
rect 7300 13908 7301 13972
rect 7235 13907 7301 13908
rect 6683 12476 6749 12477
rect 6683 12412 6684 12476
rect 6748 12412 6749 12476
rect 6683 12411 6749 12412
rect 6131 10844 6197 10845
rect 6131 10780 6132 10844
rect 6196 10780 6197 10844
rect 6131 10779 6197 10780
rect 6499 10844 6565 10845
rect 6499 10780 6500 10844
rect 6564 10780 6565 10844
rect 6499 10779 6565 10780
rect 5947 9212 6013 9213
rect 5947 9148 5948 9212
rect 6012 9148 6013 9212
rect 5947 9147 6013 9148
rect 5763 7036 5829 7037
rect 5763 6972 5764 7036
rect 5828 6972 5829 7036
rect 5763 6971 5829 6972
rect 5579 6900 5645 6901
rect 5579 6836 5580 6900
rect 5644 6836 5645 6900
rect 5579 6835 5645 6836
rect 6134 6765 6194 10779
rect 6686 8533 6746 12411
rect 7051 10844 7117 10845
rect 7051 10780 7052 10844
rect 7116 10780 7117 10844
rect 7051 10779 7117 10780
rect 6683 8532 6749 8533
rect 6683 8468 6684 8532
rect 6748 8468 6749 8532
rect 6683 8467 6749 8468
rect 7054 7989 7114 10779
rect 7051 7988 7117 7989
rect 7051 7924 7052 7988
rect 7116 7924 7117 7988
rect 7051 7923 7117 7924
rect 7238 7717 7298 13907
rect 7422 13429 7482 22747
rect 7790 22110 7850 23563
rect 7606 22050 7850 22110
rect 7606 16693 7666 22050
rect 8710 20501 8770 24787
rect 9078 22677 9138 25467
rect 9259 23492 9325 23493
rect 9259 23428 9260 23492
rect 9324 23428 9325 23492
rect 9259 23427 9325 23428
rect 9075 22676 9141 22677
rect 9075 22612 9076 22676
rect 9140 22612 9141 22676
rect 9075 22611 9141 22612
rect 8891 22404 8957 22405
rect 8891 22340 8892 22404
rect 8956 22340 8957 22404
rect 8891 22339 8957 22340
rect 8707 20500 8773 20501
rect 8707 20436 8708 20500
rect 8772 20436 8773 20500
rect 8707 20435 8773 20436
rect 8155 19684 8221 19685
rect 8155 19620 8156 19684
rect 8220 19620 8221 19684
rect 8155 19619 8221 19620
rect 7603 16692 7669 16693
rect 7603 16628 7604 16692
rect 7668 16628 7669 16692
rect 7603 16627 7669 16628
rect 8158 15741 8218 19619
rect 8707 17644 8773 17645
rect 8707 17580 8708 17644
rect 8772 17580 8773 17644
rect 8707 17579 8773 17580
rect 8155 15740 8221 15741
rect 8155 15676 8156 15740
rect 8220 15676 8221 15740
rect 8155 15675 8221 15676
rect 8339 13700 8405 13701
rect 8339 13636 8340 13700
rect 8404 13636 8405 13700
rect 8339 13635 8405 13636
rect 8155 13564 8221 13565
rect 8155 13500 8156 13564
rect 8220 13500 8221 13564
rect 8155 13499 8221 13500
rect 7419 13428 7485 13429
rect 7419 13364 7420 13428
rect 7484 13364 7485 13428
rect 7419 13363 7485 13364
rect 7422 10301 7482 13363
rect 7603 13292 7669 13293
rect 7603 13228 7604 13292
rect 7668 13228 7669 13292
rect 7603 13227 7669 13228
rect 7419 10300 7485 10301
rect 7419 10236 7420 10300
rect 7484 10236 7485 10300
rect 7419 10235 7485 10236
rect 7419 8940 7485 8941
rect 7419 8876 7420 8940
rect 7484 8876 7485 8940
rect 7419 8875 7485 8876
rect 7422 8261 7482 8875
rect 7419 8260 7485 8261
rect 7419 8196 7420 8260
rect 7484 8196 7485 8260
rect 7419 8195 7485 8196
rect 7235 7716 7301 7717
rect 7235 7652 7236 7716
rect 7300 7652 7301 7716
rect 7235 7651 7301 7652
rect 7606 6765 7666 13227
rect 7787 11932 7853 11933
rect 7787 11868 7788 11932
rect 7852 11868 7853 11932
rect 7787 11867 7853 11868
rect 7790 9621 7850 11867
rect 7971 10572 8037 10573
rect 7971 10508 7972 10572
rect 8036 10508 8037 10572
rect 7971 10507 8037 10508
rect 7787 9620 7853 9621
rect 7787 9556 7788 9620
rect 7852 9556 7853 9620
rect 7787 9555 7853 9556
rect 7974 9213 8034 10507
rect 8158 10029 8218 13499
rect 8342 12450 8402 13635
rect 8342 12390 8586 12450
rect 8155 10028 8221 10029
rect 8155 9964 8156 10028
rect 8220 9964 8221 10028
rect 8155 9963 8221 9964
rect 7971 9212 8037 9213
rect 7971 9148 7972 9212
rect 8036 9148 8037 9212
rect 7971 9147 8037 9148
rect 8158 7853 8218 9963
rect 8155 7852 8221 7853
rect 8155 7788 8156 7852
rect 8220 7788 8221 7852
rect 8155 7787 8221 7788
rect 8526 7717 8586 12390
rect 8710 9893 8770 17579
rect 8707 9892 8773 9893
rect 8707 9828 8708 9892
rect 8772 9828 8773 9892
rect 8707 9827 8773 9828
rect 8707 9212 8773 9213
rect 8707 9148 8708 9212
rect 8772 9148 8773 9212
rect 8707 9147 8773 9148
rect 8523 7716 8589 7717
rect 8523 7652 8524 7716
rect 8588 7652 8589 7716
rect 8523 7651 8589 7652
rect 6131 6764 6197 6765
rect 6131 6700 6132 6764
rect 6196 6700 6197 6764
rect 6131 6699 6197 6700
rect 7603 6764 7669 6765
rect 7603 6700 7604 6764
rect 7668 6700 7669 6764
rect 7603 6699 7669 6700
rect 8710 6221 8770 9147
rect 8894 7853 8954 22339
rect 8891 7852 8957 7853
rect 8891 7788 8892 7852
rect 8956 7788 8957 7852
rect 8891 7787 8957 7788
rect 9078 7037 9138 22611
rect 9262 22405 9322 23427
rect 9446 22949 9506 26419
rect 11099 25668 11165 25669
rect 11099 25604 11100 25668
rect 11164 25604 11165 25668
rect 11099 25603 11165 25604
rect 10363 25124 10429 25125
rect 10363 25060 10364 25124
rect 10428 25060 10429 25124
rect 10363 25059 10429 25060
rect 10179 24036 10245 24037
rect 10179 23972 10180 24036
rect 10244 23972 10245 24036
rect 10179 23971 10245 23972
rect 9443 22948 9509 22949
rect 9443 22884 9444 22948
rect 9508 22884 9509 22948
rect 9443 22883 9509 22884
rect 9259 22404 9325 22405
rect 9259 22340 9260 22404
rect 9324 22340 9325 22404
rect 9259 22339 9325 22340
rect 9443 22404 9509 22405
rect 9443 22340 9444 22404
rect 9508 22340 9509 22404
rect 9443 22339 9509 22340
rect 9259 20364 9325 20365
rect 9259 20300 9260 20364
rect 9324 20300 9325 20364
rect 9259 20299 9325 20300
rect 9262 13157 9322 20299
rect 9446 13565 9506 22339
rect 10182 21997 10242 23971
rect 10366 22949 10426 25059
rect 10915 24444 10981 24445
rect 10915 24380 10916 24444
rect 10980 24380 10981 24444
rect 10915 24379 10981 24380
rect 10547 23900 10613 23901
rect 10547 23836 10548 23900
rect 10612 23836 10613 23900
rect 10547 23835 10613 23836
rect 10363 22948 10429 22949
rect 10363 22884 10364 22948
rect 10428 22884 10429 22948
rect 10363 22883 10429 22884
rect 10363 22540 10429 22541
rect 10363 22476 10364 22540
rect 10428 22476 10429 22540
rect 10363 22475 10429 22476
rect 10179 21996 10245 21997
rect 10179 21932 10180 21996
rect 10244 21932 10245 21996
rect 10179 21931 10245 21932
rect 10179 20636 10245 20637
rect 10179 20572 10180 20636
rect 10244 20572 10245 20636
rect 10179 20571 10245 20572
rect 9627 19548 9693 19549
rect 9627 19484 9628 19548
rect 9692 19484 9693 19548
rect 9627 19483 9693 19484
rect 9630 16557 9690 19483
rect 9627 16556 9693 16557
rect 9627 16492 9628 16556
rect 9692 16492 9693 16556
rect 9627 16491 9693 16492
rect 9443 13564 9509 13565
rect 9443 13500 9444 13564
rect 9508 13500 9509 13564
rect 9443 13499 9509 13500
rect 9259 13156 9325 13157
rect 9259 13092 9260 13156
rect 9324 13092 9325 13156
rect 9259 13091 9325 13092
rect 9262 10301 9322 13091
rect 10182 11253 10242 20571
rect 10366 19549 10426 22475
rect 10363 19548 10429 19549
rect 10363 19484 10364 19548
rect 10428 19484 10429 19548
rect 10363 19483 10429 19484
rect 10550 16829 10610 23835
rect 10731 23084 10797 23085
rect 10731 23020 10732 23084
rect 10796 23020 10797 23084
rect 10731 23019 10797 23020
rect 10734 21997 10794 23019
rect 10731 21996 10797 21997
rect 10731 21932 10732 21996
rect 10796 21932 10797 21996
rect 10731 21931 10797 21932
rect 10547 16828 10613 16829
rect 10547 16764 10548 16828
rect 10612 16764 10613 16828
rect 10547 16763 10613 16764
rect 10363 13156 10429 13157
rect 10363 13092 10364 13156
rect 10428 13092 10429 13156
rect 10363 13091 10429 13092
rect 10179 11252 10245 11253
rect 10179 11188 10180 11252
rect 10244 11188 10245 11252
rect 10179 11187 10245 11188
rect 9259 10300 9325 10301
rect 9259 10236 9260 10300
rect 9324 10236 9325 10300
rect 9259 10235 9325 10236
rect 9811 10300 9877 10301
rect 9811 10236 9812 10300
rect 9876 10236 9877 10300
rect 9811 10235 9877 10236
rect 9262 7850 9322 10235
rect 9443 9892 9509 9893
rect 9443 9828 9444 9892
rect 9508 9828 9509 9892
rect 9443 9827 9509 9828
rect 9446 7989 9506 9827
rect 9814 8397 9874 10235
rect 9811 8396 9877 8397
rect 9811 8332 9812 8396
rect 9876 8332 9877 8396
rect 9811 8331 9877 8332
rect 9443 7988 9509 7989
rect 9443 7924 9444 7988
rect 9508 7924 9509 7988
rect 9443 7923 9509 7924
rect 9262 7790 9506 7850
rect 9075 7036 9141 7037
rect 9075 6972 9076 7036
rect 9140 6972 9141 7036
rect 9075 6971 9141 6972
rect 8707 6220 8773 6221
rect 8707 6156 8708 6220
rect 8772 6156 8773 6220
rect 8707 6155 8773 6156
rect 5211 5132 5277 5133
rect 5211 5068 5212 5132
rect 5276 5068 5277 5132
rect 5211 5067 5277 5068
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 9078 4861 9138 6971
rect 9446 5949 9506 7790
rect 9995 7444 10061 7445
rect 9995 7380 9996 7444
rect 10060 7380 10061 7444
rect 9995 7379 10061 7380
rect 9443 5948 9509 5949
rect 9443 5884 9444 5948
rect 9508 5884 9509 5948
rect 9443 5883 9509 5884
rect 9075 4860 9141 4861
rect 9075 4796 9076 4860
rect 9140 4796 9141 4860
rect 9075 4795 9141 4796
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 9998 3229 10058 7379
rect 10366 6901 10426 13091
rect 10550 13021 10610 16763
rect 10918 16421 10978 24379
rect 11102 22677 11162 25603
rect 11099 22676 11165 22677
rect 11099 22612 11100 22676
rect 11164 22612 11165 22676
rect 11099 22611 11165 22612
rect 11283 22676 11349 22677
rect 11283 22612 11284 22676
rect 11348 22612 11349 22676
rect 11283 22611 11349 22612
rect 11286 18597 11346 22611
rect 11838 20229 11898 26691
rect 13307 26620 13373 26621
rect 13307 26556 13308 26620
rect 13372 26556 13373 26620
rect 13307 26555 13373 26556
rect 12755 26484 12821 26485
rect 12755 26420 12756 26484
rect 12820 26420 12821 26484
rect 12755 26419 12821 26420
rect 12571 23492 12637 23493
rect 12571 23428 12572 23492
rect 12636 23428 12637 23492
rect 12571 23427 12637 23428
rect 12019 21044 12085 21045
rect 12019 20980 12020 21044
rect 12084 20980 12085 21044
rect 12019 20979 12085 20980
rect 11835 20228 11901 20229
rect 11835 20164 11836 20228
rect 11900 20164 11901 20228
rect 11835 20163 11901 20164
rect 11651 19140 11717 19141
rect 11651 19076 11652 19140
rect 11716 19076 11717 19140
rect 11651 19075 11717 19076
rect 11283 18596 11349 18597
rect 11283 18532 11284 18596
rect 11348 18532 11349 18596
rect 11283 18531 11349 18532
rect 10915 16420 10981 16421
rect 10915 16356 10916 16420
rect 10980 16356 10981 16420
rect 10915 16355 10981 16356
rect 10918 16010 10978 16355
rect 10918 15950 11162 16010
rect 10547 13020 10613 13021
rect 10547 12956 10548 13020
rect 10612 12956 10613 13020
rect 10547 12955 10613 12956
rect 10550 12069 10610 12955
rect 10547 12068 10613 12069
rect 10547 12004 10548 12068
rect 10612 12004 10613 12068
rect 10547 12003 10613 12004
rect 10550 9210 10610 12003
rect 11102 10709 11162 15950
rect 11283 11388 11349 11389
rect 11283 11324 11284 11388
rect 11348 11324 11349 11388
rect 11283 11323 11349 11324
rect 11099 10708 11165 10709
rect 11099 10644 11100 10708
rect 11164 10644 11165 10708
rect 11099 10643 11165 10644
rect 10550 9150 10794 9210
rect 10547 9076 10613 9077
rect 10547 9012 10548 9076
rect 10612 9012 10613 9076
rect 10547 9011 10613 9012
rect 10363 6900 10429 6901
rect 10363 6836 10364 6900
rect 10428 6836 10429 6900
rect 10363 6835 10429 6836
rect 10550 6085 10610 9011
rect 10734 6765 10794 9150
rect 11286 7173 11346 11323
rect 11467 8124 11533 8125
rect 11467 8060 11468 8124
rect 11532 8060 11533 8124
rect 11467 8059 11533 8060
rect 11283 7172 11349 7173
rect 11283 7108 11284 7172
rect 11348 7108 11349 7172
rect 11283 7107 11349 7108
rect 10731 6764 10797 6765
rect 10731 6700 10732 6764
rect 10796 6700 10797 6764
rect 10731 6699 10797 6700
rect 10547 6084 10613 6085
rect 10547 6020 10548 6084
rect 10612 6020 10613 6084
rect 10547 6019 10613 6020
rect 11470 5813 11530 8059
rect 11654 6085 11714 19075
rect 12022 9621 12082 20979
rect 12203 20772 12269 20773
rect 12203 20708 12204 20772
rect 12268 20708 12269 20772
rect 12203 20707 12269 20708
rect 12206 14109 12266 20707
rect 12574 20365 12634 23427
rect 12758 21317 12818 26419
rect 13123 23084 13189 23085
rect 13123 23020 13124 23084
rect 13188 23020 13189 23084
rect 13123 23019 13189 23020
rect 12755 21316 12821 21317
rect 12755 21252 12756 21316
rect 12820 21252 12821 21316
rect 12755 21251 12821 21252
rect 12758 20909 12818 21251
rect 12755 20908 12821 20909
rect 12755 20844 12756 20908
rect 12820 20844 12821 20908
rect 12755 20843 12821 20844
rect 12571 20364 12637 20365
rect 12571 20300 12572 20364
rect 12636 20300 12637 20364
rect 12571 20299 12637 20300
rect 12571 19004 12637 19005
rect 12571 18940 12572 19004
rect 12636 18940 12637 19004
rect 12571 18939 12637 18940
rect 12387 16964 12453 16965
rect 12387 16900 12388 16964
rect 12452 16900 12453 16964
rect 12387 16899 12453 16900
rect 12203 14108 12269 14109
rect 12203 14044 12204 14108
rect 12268 14044 12269 14108
rect 12203 14043 12269 14044
rect 12390 10029 12450 16899
rect 12387 10028 12453 10029
rect 12387 9964 12388 10028
rect 12452 9964 12453 10028
rect 12387 9963 12453 9964
rect 12019 9620 12085 9621
rect 12019 9556 12020 9620
rect 12084 9556 12085 9620
rect 12019 9555 12085 9556
rect 11835 7580 11901 7581
rect 11835 7516 11836 7580
rect 11900 7516 11901 7580
rect 11835 7515 11901 7516
rect 11651 6084 11717 6085
rect 11651 6020 11652 6084
rect 11716 6020 11717 6084
rect 11651 6019 11717 6020
rect 11467 5812 11533 5813
rect 11467 5748 11468 5812
rect 11532 5748 11533 5812
rect 11467 5747 11533 5748
rect 11838 5677 11898 7515
rect 12574 7309 12634 18939
rect 12939 18052 13005 18053
rect 12939 17988 12940 18052
rect 13004 17988 13005 18052
rect 12939 17987 13005 17988
rect 12755 13836 12821 13837
rect 12755 13772 12756 13836
rect 12820 13772 12821 13836
rect 12755 13771 12821 13772
rect 12758 9213 12818 13771
rect 12942 11253 13002 17987
rect 13126 14517 13186 23019
rect 13310 21725 13370 26555
rect 14043 26484 14109 26485
rect 14043 26420 14044 26484
rect 14108 26420 14109 26484
rect 14043 26419 14109 26420
rect 13491 22948 13557 22949
rect 13491 22884 13492 22948
rect 13556 22884 13557 22948
rect 13491 22883 13557 22884
rect 13307 21724 13373 21725
rect 13307 21660 13308 21724
rect 13372 21660 13373 21724
rect 13307 21659 13373 21660
rect 13307 20092 13373 20093
rect 13307 20028 13308 20092
rect 13372 20028 13373 20092
rect 13307 20027 13373 20028
rect 13123 14516 13189 14517
rect 13123 14452 13124 14516
rect 13188 14452 13189 14516
rect 13123 14451 13189 14452
rect 12939 11252 13005 11253
rect 12939 11188 12940 11252
rect 13004 11188 13005 11252
rect 12939 11187 13005 11188
rect 12939 10572 13005 10573
rect 12939 10508 12940 10572
rect 13004 10508 13005 10572
rect 12939 10507 13005 10508
rect 12755 9212 12821 9213
rect 12755 9148 12756 9212
rect 12820 9148 12821 9212
rect 12755 9147 12821 9148
rect 12571 7308 12637 7309
rect 12571 7244 12572 7308
rect 12636 7244 12637 7308
rect 12571 7243 12637 7244
rect 10731 5676 10797 5677
rect 10731 5612 10732 5676
rect 10796 5612 10797 5676
rect 10731 5611 10797 5612
rect 11835 5676 11901 5677
rect 11835 5612 11836 5676
rect 11900 5612 11901 5676
rect 11835 5611 11901 5612
rect 10734 4861 10794 5611
rect 10731 4860 10797 4861
rect 10731 4796 10732 4860
rect 10796 4796 10797 4860
rect 10731 4795 10797 4796
rect 12942 3229 13002 10507
rect 13310 9893 13370 20027
rect 13494 14653 13554 22883
rect 13675 19820 13741 19821
rect 13675 19756 13676 19820
rect 13740 19756 13741 19820
rect 13675 19755 13741 19756
rect 13678 16693 13738 19755
rect 13859 19412 13925 19413
rect 13859 19348 13860 19412
rect 13924 19348 13925 19412
rect 13859 19347 13925 19348
rect 13675 16692 13741 16693
rect 13675 16628 13676 16692
rect 13740 16628 13741 16692
rect 13675 16627 13741 16628
rect 13491 14652 13557 14653
rect 13491 14588 13492 14652
rect 13556 14588 13557 14652
rect 13491 14587 13557 14588
rect 13675 13836 13741 13837
rect 13675 13772 13676 13836
rect 13740 13772 13741 13836
rect 13675 13771 13741 13772
rect 13307 9892 13373 9893
rect 13307 9828 13308 9892
rect 13372 9828 13373 9892
rect 13307 9827 13373 9828
rect 13678 3229 13738 13771
rect 13862 12613 13922 19347
rect 13859 12612 13925 12613
rect 13859 12548 13860 12612
rect 13924 12548 13925 12612
rect 13859 12547 13925 12548
rect 13859 11796 13925 11797
rect 13859 11732 13860 11796
rect 13924 11732 13925 11796
rect 13859 11731 13925 11732
rect 13862 8261 13922 11731
rect 14046 10573 14106 26419
rect 14414 20637 14474 35939
rect 14963 34644 15029 34645
rect 14963 34580 14964 34644
rect 15028 34580 15029 34644
rect 14963 34579 15029 34580
rect 14779 30428 14845 30429
rect 14779 30364 14780 30428
rect 14844 30364 14845 30428
rect 14779 30363 14845 30364
rect 14782 21589 14842 30363
rect 14779 21588 14845 21589
rect 14779 21524 14780 21588
rect 14844 21524 14845 21588
rect 14779 21523 14845 21524
rect 14966 20637 15026 34579
rect 15147 28932 15213 28933
rect 15147 28868 15148 28932
rect 15212 28868 15213 28932
rect 15147 28867 15213 28868
rect 15150 20637 15210 28867
rect 15699 24852 15765 24853
rect 15699 24788 15700 24852
rect 15764 24788 15765 24852
rect 15699 24787 15765 24788
rect 14411 20636 14477 20637
rect 14411 20572 14412 20636
rect 14476 20572 14477 20636
rect 14411 20571 14477 20572
rect 14963 20636 15029 20637
rect 14963 20572 14964 20636
rect 15028 20572 15029 20636
rect 14963 20571 15029 20572
rect 15147 20636 15213 20637
rect 15147 20572 15148 20636
rect 15212 20572 15213 20636
rect 15147 20571 15213 20572
rect 14963 19820 15029 19821
rect 14963 19756 14964 19820
rect 15028 19756 15029 19820
rect 14963 19755 15029 19756
rect 14595 19412 14661 19413
rect 14595 19348 14596 19412
rect 14660 19348 14661 19412
rect 14595 19347 14661 19348
rect 14227 13972 14293 13973
rect 14227 13908 14228 13972
rect 14292 13908 14293 13972
rect 14227 13907 14293 13908
rect 14230 11253 14290 13907
rect 14227 11252 14293 11253
rect 14227 11188 14228 11252
rect 14292 11188 14293 11252
rect 14227 11187 14293 11188
rect 14411 11252 14477 11253
rect 14411 11188 14412 11252
rect 14476 11188 14477 11252
rect 14411 11187 14477 11188
rect 14043 10572 14109 10573
rect 14043 10508 14044 10572
rect 14108 10508 14109 10572
rect 14043 10507 14109 10508
rect 13859 8260 13925 8261
rect 13859 8196 13860 8260
rect 13924 8196 13925 8260
rect 13859 8195 13925 8196
rect 13859 5676 13925 5677
rect 13859 5612 13860 5676
rect 13924 5612 13925 5676
rect 13859 5611 13925 5612
rect 13862 3637 13922 5611
rect 14230 4045 14290 11187
rect 14414 9893 14474 11187
rect 14411 9892 14477 9893
rect 14411 9828 14412 9892
rect 14476 9828 14477 9892
rect 14411 9827 14477 9828
rect 14598 7581 14658 19347
rect 14779 10572 14845 10573
rect 14779 10508 14780 10572
rect 14844 10508 14845 10572
rect 14779 10507 14845 10508
rect 14595 7580 14661 7581
rect 14595 7516 14596 7580
rect 14660 7516 14661 7580
rect 14595 7515 14661 7516
rect 14227 4044 14293 4045
rect 14227 3980 14228 4044
rect 14292 3980 14293 4044
rect 14227 3979 14293 3980
rect 13859 3636 13925 3637
rect 13859 3572 13860 3636
rect 13924 3572 13925 3636
rect 13859 3571 13925 3572
rect 14782 3365 14842 10507
rect 14966 8261 15026 19755
rect 15702 19350 15762 24787
rect 15886 22813 15946 37299
rect 16987 36548 17053 36549
rect 16987 36484 16988 36548
rect 17052 36484 17053 36548
rect 16987 36483 17053 36484
rect 17723 36548 17789 36549
rect 17723 36484 17724 36548
rect 17788 36484 17789 36548
rect 17723 36483 17789 36484
rect 16067 27028 16133 27029
rect 16067 26964 16068 27028
rect 16132 26964 16133 27028
rect 16067 26963 16133 26964
rect 15883 22812 15949 22813
rect 15883 22748 15884 22812
rect 15948 22748 15949 22812
rect 15883 22747 15949 22748
rect 15886 21453 15946 22747
rect 15883 21452 15949 21453
rect 15883 21388 15884 21452
rect 15948 21388 15949 21452
rect 15883 21387 15949 21388
rect 15883 21044 15949 21045
rect 15883 20980 15884 21044
rect 15948 20980 15949 21044
rect 15883 20979 15949 20980
rect 15518 19290 15762 19350
rect 15518 18597 15578 19290
rect 15515 18596 15581 18597
rect 15515 18532 15516 18596
rect 15580 18532 15581 18596
rect 15515 18531 15581 18532
rect 15518 17917 15578 18531
rect 15515 17916 15581 17917
rect 15515 17852 15516 17916
rect 15580 17852 15581 17916
rect 15515 17851 15581 17852
rect 15886 15330 15946 20979
rect 16070 19277 16130 26963
rect 16803 23492 16869 23493
rect 16803 23428 16804 23492
rect 16868 23428 16869 23492
rect 16803 23427 16869 23428
rect 16251 21452 16317 21453
rect 16251 21388 16252 21452
rect 16316 21388 16317 21452
rect 16251 21387 16317 21388
rect 16254 21045 16314 21387
rect 16251 21044 16317 21045
rect 16251 20980 16252 21044
rect 16316 20980 16317 21044
rect 16251 20979 16317 20980
rect 16251 20772 16317 20773
rect 16251 20708 16252 20772
rect 16316 20708 16317 20772
rect 16251 20707 16317 20708
rect 16067 19276 16133 19277
rect 16067 19212 16068 19276
rect 16132 19212 16133 19276
rect 16067 19211 16133 19212
rect 16067 15876 16133 15877
rect 16067 15812 16068 15876
rect 16132 15812 16133 15876
rect 16067 15811 16133 15812
rect 15702 15270 15946 15330
rect 15702 14109 15762 15270
rect 15699 14108 15765 14109
rect 15699 14044 15700 14108
rect 15764 14044 15765 14108
rect 15699 14043 15765 14044
rect 15331 8396 15397 8397
rect 15331 8332 15332 8396
rect 15396 8332 15397 8396
rect 15331 8331 15397 8332
rect 14963 8260 15029 8261
rect 14963 8196 14964 8260
rect 15028 8196 15029 8260
rect 14963 8195 15029 8196
rect 15147 7580 15213 7581
rect 15147 7516 15148 7580
rect 15212 7516 15213 7580
rect 15147 7515 15213 7516
rect 14779 3364 14845 3365
rect 14779 3300 14780 3364
rect 14844 3300 14845 3364
rect 14779 3299 14845 3300
rect 9995 3228 10061 3229
rect 9995 3164 9996 3228
rect 10060 3164 10061 3228
rect 9995 3163 10061 3164
rect 12939 3228 13005 3229
rect 12939 3164 12940 3228
rect 13004 3164 13005 3228
rect 12939 3163 13005 3164
rect 13675 3228 13741 3229
rect 13675 3164 13676 3228
rect 13740 3164 13741 3228
rect 13675 3163 13741 3164
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 15150 2141 15210 7515
rect 15334 4045 15394 8331
rect 15515 8260 15581 8261
rect 15515 8196 15516 8260
rect 15580 8196 15581 8260
rect 15515 8195 15581 8196
rect 15331 4044 15397 4045
rect 15331 3980 15332 4044
rect 15396 3980 15397 4044
rect 15331 3979 15397 3980
rect 15518 2685 15578 8195
rect 16070 8125 16130 15811
rect 16254 9213 16314 20707
rect 16435 20636 16501 20637
rect 16435 20572 16436 20636
rect 16500 20572 16501 20636
rect 16435 20571 16501 20572
rect 16251 9212 16317 9213
rect 16251 9148 16252 9212
rect 16316 9148 16317 9212
rect 16251 9147 16317 9148
rect 16067 8124 16133 8125
rect 16067 8060 16068 8124
rect 16132 8060 16133 8124
rect 16067 8059 16133 8060
rect 16438 7853 16498 20571
rect 16619 19684 16685 19685
rect 16619 19620 16620 19684
rect 16684 19620 16685 19684
rect 16619 19619 16685 19620
rect 16622 9485 16682 19619
rect 16806 19277 16866 23427
rect 16990 21997 17050 36483
rect 17539 34644 17605 34645
rect 17539 34580 17540 34644
rect 17604 34580 17605 34644
rect 17539 34579 17605 34580
rect 17171 23764 17237 23765
rect 17171 23700 17172 23764
rect 17236 23700 17237 23764
rect 17171 23699 17237 23700
rect 16987 21996 17053 21997
rect 16987 21932 16988 21996
rect 17052 21932 17053 21996
rect 16987 21931 17053 21932
rect 16987 20908 17053 20909
rect 16987 20844 16988 20908
rect 17052 20844 17053 20908
rect 16987 20843 17053 20844
rect 16803 19276 16869 19277
rect 16803 19212 16804 19276
rect 16868 19212 16869 19276
rect 16803 19211 16869 19212
rect 16803 18596 16869 18597
rect 16803 18532 16804 18596
rect 16868 18532 16869 18596
rect 16803 18531 16869 18532
rect 16806 15333 16866 18531
rect 16803 15332 16869 15333
rect 16803 15268 16804 15332
rect 16868 15268 16869 15332
rect 16803 15267 16869 15268
rect 16990 14109 17050 20843
rect 17174 17917 17234 23699
rect 17542 23493 17602 34579
rect 17539 23492 17605 23493
rect 17539 23428 17540 23492
rect 17604 23428 17605 23492
rect 17539 23427 17605 23428
rect 17355 22540 17421 22541
rect 17355 22476 17356 22540
rect 17420 22476 17421 22540
rect 17355 22475 17421 22476
rect 17171 17916 17237 17917
rect 17171 17852 17172 17916
rect 17236 17852 17237 17916
rect 17171 17851 17237 17852
rect 17171 14788 17237 14789
rect 17171 14724 17172 14788
rect 17236 14724 17237 14788
rect 17171 14723 17237 14724
rect 16987 14108 17053 14109
rect 16987 14044 16988 14108
rect 17052 14044 17053 14108
rect 16987 14043 17053 14044
rect 16803 12884 16869 12885
rect 16803 12820 16804 12884
rect 16868 12820 16869 12884
rect 16803 12819 16869 12820
rect 16619 9484 16685 9485
rect 16619 9420 16620 9484
rect 16684 9420 16685 9484
rect 16619 9419 16685 9420
rect 16806 8941 16866 12819
rect 16987 12340 17053 12341
rect 16987 12276 16988 12340
rect 17052 12276 17053 12340
rect 16987 12275 17053 12276
rect 16803 8940 16869 8941
rect 16803 8876 16804 8940
rect 16868 8876 16869 8940
rect 16803 8875 16869 8876
rect 16435 7852 16501 7853
rect 16435 7788 16436 7852
rect 16500 7788 16501 7852
rect 16435 7787 16501 7788
rect 16990 7037 17050 12275
rect 17174 9621 17234 14723
rect 17358 11389 17418 22475
rect 17726 21861 17786 36483
rect 17907 30564 17973 30565
rect 17907 30500 17908 30564
rect 17972 30500 17973 30564
rect 17907 30499 17973 30500
rect 17723 21860 17789 21861
rect 17723 21796 17724 21860
rect 17788 21796 17789 21860
rect 17723 21795 17789 21796
rect 17910 17917 17970 30499
rect 18094 23221 18154 37435
rect 19568 37024 19888 37584
rect 22507 37572 22508 37636
rect 22572 37572 22573 37636
rect 22507 37571 22573 37572
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19379 36140 19445 36141
rect 19379 36076 19380 36140
rect 19444 36076 19445 36140
rect 19379 36075 19445 36076
rect 18459 28524 18525 28525
rect 18459 28460 18460 28524
rect 18524 28460 18525 28524
rect 18459 28459 18525 28460
rect 18091 23220 18157 23221
rect 18091 23156 18092 23220
rect 18156 23156 18157 23220
rect 18091 23155 18157 23156
rect 18094 19277 18154 23155
rect 18275 22404 18341 22405
rect 18275 22340 18276 22404
rect 18340 22340 18341 22404
rect 18275 22339 18341 22340
rect 18091 19276 18157 19277
rect 18091 19212 18092 19276
rect 18156 19212 18157 19276
rect 18091 19211 18157 19212
rect 18091 18052 18157 18053
rect 18091 17988 18092 18052
rect 18156 17988 18157 18052
rect 18091 17987 18157 17988
rect 17907 17916 17973 17917
rect 17907 17852 17908 17916
rect 17972 17852 17973 17916
rect 17907 17851 17973 17852
rect 17723 17644 17789 17645
rect 17723 17580 17724 17644
rect 17788 17580 17789 17644
rect 17723 17579 17789 17580
rect 17539 12204 17605 12205
rect 17539 12140 17540 12204
rect 17604 12140 17605 12204
rect 17539 12139 17605 12140
rect 17355 11388 17421 11389
rect 17355 11324 17356 11388
rect 17420 11324 17421 11388
rect 17355 11323 17421 11324
rect 17542 10845 17602 12139
rect 17539 10844 17605 10845
rect 17539 10780 17540 10844
rect 17604 10780 17605 10844
rect 17539 10779 17605 10780
rect 17355 10300 17421 10301
rect 17355 10236 17356 10300
rect 17420 10236 17421 10300
rect 17355 10235 17421 10236
rect 17171 9620 17237 9621
rect 17171 9556 17172 9620
rect 17236 9556 17237 9620
rect 17171 9555 17237 9556
rect 17358 7853 17418 10235
rect 17726 9349 17786 17579
rect 18094 16285 18154 17987
rect 18091 16284 18157 16285
rect 18091 16220 18092 16284
rect 18156 16220 18157 16284
rect 18091 16219 18157 16220
rect 18091 15740 18157 15741
rect 18091 15676 18092 15740
rect 18156 15676 18157 15740
rect 18091 15675 18157 15676
rect 17907 15196 17973 15197
rect 17907 15132 17908 15196
rect 17972 15132 17973 15196
rect 17907 15131 17973 15132
rect 17910 12341 17970 15131
rect 18094 12885 18154 15675
rect 18091 12884 18157 12885
rect 18091 12820 18092 12884
rect 18156 12820 18157 12884
rect 18091 12819 18157 12820
rect 17907 12340 17973 12341
rect 17907 12276 17908 12340
rect 17972 12276 17973 12340
rect 17907 12275 17973 12276
rect 18278 9485 18338 22339
rect 18462 20773 18522 28459
rect 18643 21860 18709 21861
rect 18643 21796 18644 21860
rect 18708 21796 18709 21860
rect 18643 21795 18709 21796
rect 18459 20772 18525 20773
rect 18459 20708 18460 20772
rect 18524 20708 18525 20772
rect 18459 20707 18525 20708
rect 18646 19350 18706 21795
rect 18462 19290 18706 19350
rect 18462 16965 18522 19290
rect 19382 19277 19442 36075
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 20483 27980 20549 27981
rect 20483 27916 20484 27980
rect 20548 27916 20549 27980
rect 20483 27915 20549 27916
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 20299 24172 20365 24173
rect 20299 24108 20300 24172
rect 20364 24108 20365 24172
rect 20299 24107 20365 24108
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 20302 20773 20362 24107
rect 20299 20772 20365 20773
rect 20299 20708 20300 20772
rect 20364 20708 20365 20772
rect 20299 20707 20365 20708
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19379 19276 19445 19277
rect 19379 19212 19380 19276
rect 19444 19212 19445 19276
rect 19379 19211 19445 19212
rect 19379 19140 19445 19141
rect 19379 19076 19380 19140
rect 19444 19076 19445 19140
rect 19379 19075 19445 19076
rect 19011 17644 19077 17645
rect 19011 17580 19012 17644
rect 19076 17580 19077 17644
rect 19011 17579 19077 17580
rect 18459 16964 18525 16965
rect 18459 16900 18460 16964
rect 18524 16900 18525 16964
rect 18459 16899 18525 16900
rect 19014 16693 19074 17579
rect 19195 17372 19261 17373
rect 19195 17308 19196 17372
rect 19260 17308 19261 17372
rect 19195 17307 19261 17308
rect 19011 16692 19077 16693
rect 19011 16628 19012 16692
rect 19076 16628 19077 16692
rect 19011 16627 19077 16628
rect 18827 16556 18893 16557
rect 18827 16492 18828 16556
rect 18892 16492 18893 16556
rect 18827 16491 18893 16492
rect 18459 14652 18525 14653
rect 18459 14588 18460 14652
rect 18524 14588 18525 14652
rect 18459 14587 18525 14588
rect 18462 13293 18522 14587
rect 18643 14108 18709 14109
rect 18643 14044 18644 14108
rect 18708 14044 18709 14108
rect 18643 14043 18709 14044
rect 18459 13292 18525 13293
rect 18459 13228 18460 13292
rect 18524 13228 18525 13292
rect 18459 13227 18525 13228
rect 18459 13156 18525 13157
rect 18459 13092 18460 13156
rect 18524 13092 18525 13156
rect 18459 13091 18525 13092
rect 18275 9484 18341 9485
rect 18275 9420 18276 9484
rect 18340 9420 18341 9484
rect 18275 9419 18341 9420
rect 17723 9348 17789 9349
rect 17723 9284 17724 9348
rect 17788 9284 17789 9348
rect 17723 9283 17789 9284
rect 17539 9212 17605 9213
rect 17539 9148 17540 9212
rect 17604 9148 17605 9212
rect 17539 9147 17605 9148
rect 18091 9212 18157 9213
rect 18091 9148 18092 9212
rect 18156 9148 18157 9212
rect 18091 9147 18157 9148
rect 17355 7852 17421 7853
rect 17355 7788 17356 7852
rect 17420 7788 17421 7852
rect 17355 7787 17421 7788
rect 16987 7036 17053 7037
rect 16987 6972 16988 7036
rect 17052 6972 17053 7036
rect 16987 6971 17053 6972
rect 16987 5948 17053 5949
rect 16987 5884 16988 5948
rect 17052 5884 17053 5948
rect 16987 5883 17053 5884
rect 16619 4452 16685 4453
rect 16619 4388 16620 4452
rect 16684 4388 16685 4452
rect 16619 4387 16685 4388
rect 16622 3093 16682 4387
rect 16990 4181 17050 5883
rect 17171 5812 17237 5813
rect 17171 5748 17172 5812
rect 17236 5748 17237 5812
rect 17171 5747 17237 5748
rect 17174 4861 17234 5747
rect 17542 5677 17602 9147
rect 18094 8310 18154 9147
rect 17910 8250 18154 8310
rect 17910 7445 17970 8250
rect 18462 8125 18522 13091
rect 18646 12477 18706 14043
rect 18643 12476 18709 12477
rect 18643 12412 18644 12476
rect 18708 12412 18709 12476
rect 18643 12411 18709 12412
rect 18643 12068 18709 12069
rect 18643 12004 18644 12068
rect 18708 12004 18709 12068
rect 18643 12003 18709 12004
rect 18646 9485 18706 12003
rect 18830 9621 18890 16491
rect 19011 16420 19077 16421
rect 19011 16356 19012 16420
rect 19076 16356 19077 16420
rect 19011 16355 19077 16356
rect 19014 11933 19074 16355
rect 19198 15197 19258 17307
rect 19382 16829 19442 19075
rect 19568 18528 19888 19552
rect 20299 18732 20365 18733
rect 20299 18668 20300 18732
rect 20364 18668 20365 18732
rect 20299 18667 20365 18668
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 20115 18052 20181 18053
rect 20115 17988 20116 18052
rect 20180 17988 20181 18052
rect 20115 17987 20181 17988
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19379 16828 19445 16829
rect 19379 16764 19380 16828
rect 19444 16764 19445 16828
rect 19379 16763 19445 16764
rect 19379 16692 19445 16693
rect 19379 16628 19380 16692
rect 19444 16628 19445 16692
rect 19379 16627 19445 16628
rect 19195 15196 19261 15197
rect 19195 15132 19196 15196
rect 19260 15132 19261 15196
rect 19195 15131 19261 15132
rect 19382 14789 19442 16627
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19379 14788 19445 14789
rect 19379 14724 19380 14788
rect 19444 14724 19445 14788
rect 19379 14723 19445 14724
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19379 13156 19445 13157
rect 19379 13092 19380 13156
rect 19444 13092 19445 13156
rect 19379 13091 19445 13092
rect 19011 11932 19077 11933
rect 19011 11868 19012 11932
rect 19076 11868 19077 11932
rect 19011 11867 19077 11868
rect 19195 10844 19261 10845
rect 19195 10780 19196 10844
rect 19260 10780 19261 10844
rect 19195 10779 19261 10780
rect 19011 9892 19077 9893
rect 19011 9828 19012 9892
rect 19076 9828 19077 9892
rect 19011 9827 19077 9828
rect 19014 9621 19074 9827
rect 18827 9620 18893 9621
rect 18827 9556 18828 9620
rect 18892 9556 18893 9620
rect 18827 9555 18893 9556
rect 19011 9620 19077 9621
rect 19011 9556 19012 9620
rect 19076 9556 19077 9620
rect 19011 9555 19077 9556
rect 18643 9484 18709 9485
rect 18643 9420 18644 9484
rect 18708 9420 18709 9484
rect 18643 9419 18709 9420
rect 18459 8124 18525 8125
rect 18459 8060 18460 8124
rect 18524 8060 18525 8124
rect 18459 8059 18525 8060
rect 17907 7444 17973 7445
rect 17907 7380 17908 7444
rect 17972 7380 17973 7444
rect 17907 7379 17973 7380
rect 17907 7036 17973 7037
rect 17907 6972 17908 7036
rect 17972 6972 17973 7036
rect 17907 6971 17973 6972
rect 17539 5676 17605 5677
rect 17539 5612 17540 5676
rect 17604 5612 17605 5676
rect 17539 5611 17605 5612
rect 17171 4860 17237 4861
rect 17171 4796 17172 4860
rect 17236 4796 17237 4860
rect 17171 4795 17237 4796
rect 17355 4452 17421 4453
rect 17355 4388 17356 4452
rect 17420 4388 17421 4452
rect 17355 4387 17421 4388
rect 16987 4180 17053 4181
rect 16987 4116 16988 4180
rect 17052 4116 17053 4180
rect 16987 4115 17053 4116
rect 16619 3092 16685 3093
rect 16619 3028 16620 3092
rect 16684 3028 16685 3092
rect 16619 3027 16685 3028
rect 15515 2684 15581 2685
rect 15515 2620 15516 2684
rect 15580 2620 15581 2684
rect 15515 2619 15581 2620
rect 15147 2140 15213 2141
rect 15147 2076 15148 2140
rect 15212 2076 15213 2140
rect 15147 2075 15213 2076
rect 17358 1461 17418 4387
rect 17542 1597 17602 5611
rect 17910 2685 17970 6971
rect 19014 5405 19074 9555
rect 19011 5404 19077 5405
rect 19011 5340 19012 5404
rect 19076 5340 19077 5404
rect 19011 5339 19077 5340
rect 17907 2684 17973 2685
rect 17907 2620 17908 2684
rect 17972 2620 17973 2684
rect 17907 2619 17973 2620
rect 19198 2413 19258 10779
rect 19382 8261 19442 13091
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19379 8260 19445 8261
rect 19379 8196 19380 8260
rect 19444 8196 19445 8260
rect 19379 8195 19445 8196
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 20118 7445 20178 17987
rect 20302 17917 20362 18667
rect 20299 17916 20365 17917
rect 20299 17852 20300 17916
rect 20364 17852 20365 17916
rect 20299 17851 20365 17852
rect 20299 16828 20365 16829
rect 20299 16764 20300 16828
rect 20364 16764 20365 16828
rect 20299 16763 20365 16764
rect 20302 15333 20362 16763
rect 20299 15332 20365 15333
rect 20299 15268 20300 15332
rect 20364 15268 20365 15332
rect 20299 15267 20365 15268
rect 20299 14788 20365 14789
rect 20299 14724 20300 14788
rect 20364 14724 20365 14788
rect 20299 14723 20365 14724
rect 20302 11797 20362 14723
rect 20486 12205 20546 27915
rect 21035 26348 21101 26349
rect 21035 26284 21036 26348
rect 21100 26284 21101 26348
rect 21035 26283 21101 26284
rect 20667 24852 20733 24853
rect 20667 24788 20668 24852
rect 20732 24788 20733 24852
rect 20667 24787 20733 24788
rect 20670 18869 20730 24787
rect 20851 24580 20917 24581
rect 20851 24516 20852 24580
rect 20916 24516 20917 24580
rect 20851 24515 20917 24516
rect 20667 18868 20733 18869
rect 20667 18804 20668 18868
rect 20732 18804 20733 18868
rect 20667 18803 20733 18804
rect 20670 17917 20730 18803
rect 20667 17916 20733 17917
rect 20667 17852 20668 17916
rect 20732 17852 20733 17916
rect 20667 17851 20733 17852
rect 20667 17644 20733 17645
rect 20667 17580 20668 17644
rect 20732 17580 20733 17644
rect 20667 17579 20733 17580
rect 20670 12341 20730 17579
rect 20854 16693 20914 24515
rect 21038 17917 21098 26283
rect 21771 24444 21837 24445
rect 21771 24380 21772 24444
rect 21836 24380 21837 24444
rect 21771 24379 21837 24380
rect 21774 22110 21834 24379
rect 21774 22050 22018 22110
rect 21403 20908 21469 20909
rect 21403 20844 21404 20908
rect 21468 20844 21469 20908
rect 21403 20843 21469 20844
rect 21219 19548 21285 19549
rect 21219 19484 21220 19548
rect 21284 19484 21285 19548
rect 21219 19483 21285 19484
rect 21035 17916 21101 17917
rect 21035 17852 21036 17916
rect 21100 17852 21101 17916
rect 21035 17851 21101 17852
rect 20851 16692 20917 16693
rect 20851 16628 20852 16692
rect 20916 16628 20917 16692
rect 20851 16627 20917 16628
rect 21222 16557 21282 19483
rect 21219 16556 21285 16557
rect 21219 16492 21220 16556
rect 21284 16492 21285 16556
rect 21219 16491 21285 16492
rect 20851 16420 20917 16421
rect 20851 16356 20852 16420
rect 20916 16356 20917 16420
rect 20851 16355 20917 16356
rect 20854 15197 20914 16355
rect 20851 15196 20917 15197
rect 20851 15132 20852 15196
rect 20916 15132 20917 15196
rect 20851 15131 20917 15132
rect 20851 13972 20917 13973
rect 20851 13908 20852 13972
rect 20916 13908 20917 13972
rect 20851 13907 20917 13908
rect 20667 12340 20733 12341
rect 20667 12276 20668 12340
rect 20732 12276 20733 12340
rect 20667 12275 20733 12276
rect 20483 12204 20549 12205
rect 20483 12140 20484 12204
rect 20548 12140 20549 12204
rect 20483 12139 20549 12140
rect 20667 12068 20733 12069
rect 20667 12004 20668 12068
rect 20732 12004 20733 12068
rect 20667 12003 20733 12004
rect 20483 11932 20549 11933
rect 20483 11868 20484 11932
rect 20548 11868 20549 11932
rect 20483 11867 20549 11868
rect 20299 11796 20365 11797
rect 20299 11732 20300 11796
rect 20364 11732 20365 11796
rect 20299 11731 20365 11732
rect 20486 10301 20546 11867
rect 20483 10300 20549 10301
rect 20483 10236 20484 10300
rect 20548 10236 20549 10300
rect 20483 10235 20549 10236
rect 20299 9892 20365 9893
rect 20299 9828 20300 9892
rect 20364 9828 20365 9892
rect 20299 9827 20365 9828
rect 20115 7444 20181 7445
rect 20115 7380 20116 7444
rect 20180 7380 20181 7444
rect 20115 7379 20181 7380
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19379 5676 19445 5677
rect 19379 5612 19380 5676
rect 19444 5612 19445 5676
rect 19379 5611 19445 5612
rect 19382 2549 19442 5611
rect 19568 5472 19888 6496
rect 20302 5949 20362 9827
rect 20483 9756 20549 9757
rect 20483 9692 20484 9756
rect 20548 9692 20549 9756
rect 20483 9691 20549 9692
rect 20486 6357 20546 9691
rect 20483 6356 20549 6357
rect 20483 6292 20484 6356
rect 20548 6292 20549 6356
rect 20483 6291 20549 6292
rect 20299 5948 20365 5949
rect 20299 5884 20300 5948
rect 20364 5884 20365 5948
rect 20299 5883 20365 5884
rect 20483 5812 20549 5813
rect 20483 5748 20484 5812
rect 20548 5748 20549 5812
rect 20483 5747 20549 5748
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19379 2548 19445 2549
rect 19379 2484 19380 2548
rect 19444 2484 19445 2548
rect 19379 2483 19445 2484
rect 19195 2412 19261 2413
rect 19195 2348 19196 2412
rect 19260 2348 19261 2412
rect 19195 2347 19261 2348
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 17539 1596 17605 1597
rect 17539 1532 17540 1596
rect 17604 1532 17605 1596
rect 17539 1531 17605 1532
rect 17355 1460 17421 1461
rect 17355 1396 17356 1460
rect 17420 1396 17421 1460
rect 17355 1395 17421 1396
rect 20486 1325 20546 5747
rect 20670 5677 20730 12003
rect 20854 8125 20914 13907
rect 21035 12068 21101 12069
rect 21035 12004 21036 12068
rect 21100 12004 21101 12068
rect 21035 12003 21101 12004
rect 21038 9757 21098 12003
rect 21406 11389 21466 20843
rect 21958 19549 22018 22050
rect 22139 20772 22205 20773
rect 22139 20708 22140 20772
rect 22204 20708 22205 20772
rect 22139 20707 22205 20708
rect 21955 19548 22021 19549
rect 21955 19484 21956 19548
rect 22020 19484 22021 19548
rect 21955 19483 22021 19484
rect 22142 19277 22202 20707
rect 22323 19684 22389 19685
rect 22323 19620 22324 19684
rect 22388 19620 22389 19684
rect 22323 19619 22389 19620
rect 22139 19276 22205 19277
rect 22139 19212 22140 19276
rect 22204 19212 22205 19276
rect 22139 19211 22205 19212
rect 22139 16828 22205 16829
rect 22139 16764 22140 16828
rect 22204 16764 22205 16828
rect 22139 16763 22205 16764
rect 21587 15196 21653 15197
rect 21587 15132 21588 15196
rect 21652 15132 21653 15196
rect 21587 15131 21653 15132
rect 21403 11388 21469 11389
rect 21403 11324 21404 11388
rect 21468 11324 21469 11388
rect 21403 11323 21469 11324
rect 21590 10437 21650 15131
rect 22142 13565 22202 16763
rect 22139 13564 22205 13565
rect 22139 13500 22140 13564
rect 22204 13500 22205 13564
rect 22139 13499 22205 13500
rect 22326 12613 22386 19619
rect 22510 19005 22570 37571
rect 23979 37364 24045 37365
rect 23979 37300 23980 37364
rect 24044 37300 24045 37364
rect 23979 37299 24045 37300
rect 22691 32468 22757 32469
rect 22691 32404 22692 32468
rect 22756 32404 22757 32468
rect 22691 32403 22757 32404
rect 22694 20637 22754 32403
rect 23427 28116 23493 28117
rect 23427 28052 23428 28116
rect 23492 28052 23493 28116
rect 23427 28051 23493 28052
rect 22691 20636 22757 20637
rect 22691 20572 22692 20636
rect 22756 20572 22757 20636
rect 22691 20571 22757 20572
rect 22507 19004 22573 19005
rect 22507 18940 22508 19004
rect 22572 18940 22573 19004
rect 22507 18939 22573 18940
rect 22691 18052 22757 18053
rect 22691 17988 22692 18052
rect 22756 17988 22757 18052
rect 22691 17987 22757 17988
rect 22507 17916 22573 17917
rect 22507 17852 22508 17916
rect 22572 17852 22573 17916
rect 22507 17851 22573 17852
rect 22510 13429 22570 17851
rect 22507 13428 22573 13429
rect 22507 13364 22508 13428
rect 22572 13364 22573 13428
rect 22507 13363 22573 13364
rect 22323 12612 22389 12613
rect 22323 12548 22324 12612
rect 22388 12548 22389 12612
rect 22323 12547 22389 12548
rect 21587 10436 21653 10437
rect 21587 10372 21588 10436
rect 21652 10372 21653 10436
rect 21587 10371 21653 10372
rect 21771 10436 21837 10437
rect 21771 10372 21772 10436
rect 21836 10372 21837 10436
rect 21771 10371 21837 10372
rect 21035 9756 21101 9757
rect 21035 9692 21036 9756
rect 21100 9692 21101 9756
rect 21035 9691 21101 9692
rect 20851 8124 20917 8125
rect 20851 8060 20852 8124
rect 20916 8060 20917 8124
rect 20851 8059 20917 8060
rect 20667 5676 20733 5677
rect 20667 5612 20668 5676
rect 20732 5612 20733 5676
rect 20667 5611 20733 5612
rect 20667 4180 20733 4181
rect 20667 4116 20668 4180
rect 20732 4116 20733 4180
rect 20667 4115 20733 4116
rect 20483 1324 20549 1325
rect 20483 1260 20484 1324
rect 20548 1260 20549 1324
rect 20483 1259 20549 1260
rect 20670 237 20730 4115
rect 21774 645 21834 10371
rect 22694 8125 22754 17987
rect 23430 14109 23490 28051
rect 23982 14925 24042 37299
rect 26739 34644 26805 34645
rect 26739 34580 26740 34644
rect 26804 34580 26805 34644
rect 26739 34579 26805 34580
rect 26003 32468 26069 32469
rect 26003 32404 26004 32468
rect 26068 32404 26069 32468
rect 26003 32403 26069 32404
rect 25451 29340 25517 29341
rect 25451 29276 25452 29340
rect 25516 29276 25517 29340
rect 25451 29275 25517 29276
rect 24899 26892 24965 26893
rect 24899 26828 24900 26892
rect 24964 26828 24965 26892
rect 24899 26827 24965 26828
rect 24531 21452 24597 21453
rect 24531 21388 24532 21452
rect 24596 21388 24597 21452
rect 24531 21387 24597 21388
rect 24163 21044 24229 21045
rect 24163 20980 24164 21044
rect 24228 20980 24229 21044
rect 24163 20979 24229 20980
rect 23979 14924 24045 14925
rect 23979 14860 23980 14924
rect 24044 14860 24045 14924
rect 23979 14859 24045 14860
rect 23427 14108 23493 14109
rect 23427 14044 23428 14108
rect 23492 14044 23493 14108
rect 23427 14043 23493 14044
rect 23427 13972 23493 13973
rect 23427 13908 23428 13972
rect 23492 13908 23493 13972
rect 23427 13907 23493 13908
rect 23430 10981 23490 13907
rect 23611 11524 23677 11525
rect 23611 11460 23612 11524
rect 23676 11460 23677 11524
rect 23611 11459 23677 11460
rect 23795 11524 23861 11525
rect 23795 11460 23796 11524
rect 23860 11460 23861 11524
rect 23795 11459 23861 11460
rect 23427 10980 23493 10981
rect 23427 10916 23428 10980
rect 23492 10916 23493 10980
rect 23427 10915 23493 10916
rect 23427 9620 23493 9621
rect 23427 9556 23428 9620
rect 23492 9556 23493 9620
rect 23427 9555 23493 9556
rect 23059 9348 23125 9349
rect 23059 9284 23060 9348
rect 23124 9284 23125 9348
rect 23059 9283 23125 9284
rect 22691 8124 22757 8125
rect 22691 8060 22692 8124
rect 22756 8060 22757 8124
rect 22691 8059 22757 8060
rect 22139 5676 22205 5677
rect 22139 5612 22140 5676
rect 22204 5612 22205 5676
rect 22139 5611 22205 5612
rect 21771 644 21837 645
rect 21771 580 21772 644
rect 21836 580 21837 644
rect 21771 579 21837 580
rect 20667 236 20733 237
rect 20667 172 20668 236
rect 20732 172 20733 236
rect 20667 171 20733 172
rect 22142 101 22202 5611
rect 23062 3229 23122 9283
rect 23430 5541 23490 9555
rect 23427 5540 23493 5541
rect 23427 5476 23428 5540
rect 23492 5476 23493 5540
rect 23427 5475 23493 5476
rect 23427 4180 23493 4181
rect 23427 4116 23428 4180
rect 23492 4116 23493 4180
rect 23427 4115 23493 4116
rect 23059 3228 23125 3229
rect 23059 3164 23060 3228
rect 23124 3164 23125 3228
rect 23059 3163 23125 3164
rect 23430 781 23490 4115
rect 23614 2413 23674 11459
rect 23611 2412 23677 2413
rect 23611 2348 23612 2412
rect 23676 2348 23677 2412
rect 23611 2347 23677 2348
rect 23798 1325 23858 11459
rect 24166 9621 24226 20979
rect 24534 11389 24594 21387
rect 24902 18461 24962 26827
rect 25083 23628 25149 23629
rect 25083 23564 25084 23628
rect 25148 23564 25149 23628
rect 25083 23563 25149 23564
rect 25086 19413 25146 23563
rect 25267 19956 25333 19957
rect 25267 19892 25268 19956
rect 25332 19892 25333 19956
rect 25267 19891 25333 19892
rect 25083 19412 25149 19413
rect 25083 19348 25084 19412
rect 25148 19348 25149 19412
rect 25083 19347 25149 19348
rect 24899 18460 24965 18461
rect 24899 18396 24900 18460
rect 24964 18396 24965 18460
rect 24899 18395 24965 18396
rect 24899 18324 24965 18325
rect 24899 18260 24900 18324
rect 24964 18260 24965 18324
rect 24899 18259 24965 18260
rect 24902 15197 24962 18259
rect 24899 15196 24965 15197
rect 24899 15132 24900 15196
rect 24964 15132 24965 15196
rect 24899 15131 24965 15132
rect 25083 15196 25149 15197
rect 25083 15132 25084 15196
rect 25148 15132 25149 15196
rect 25083 15131 25149 15132
rect 24531 11388 24597 11389
rect 24531 11324 24532 11388
rect 24596 11324 24597 11388
rect 24531 11323 24597 11324
rect 24163 9620 24229 9621
rect 24163 9556 24164 9620
rect 24228 9556 24229 9620
rect 24163 9555 24229 9556
rect 25086 6085 25146 15131
rect 25270 9213 25330 19891
rect 25454 19277 25514 29275
rect 25819 19820 25885 19821
rect 25819 19756 25820 19820
rect 25884 19756 25885 19820
rect 25819 19755 25885 19756
rect 25451 19276 25517 19277
rect 25451 19212 25452 19276
rect 25516 19212 25517 19276
rect 25451 19211 25517 19212
rect 25822 9621 25882 19755
rect 26006 19413 26066 32403
rect 26003 19412 26069 19413
rect 26003 19348 26004 19412
rect 26068 19348 26069 19412
rect 26003 19347 26069 19348
rect 26555 18596 26621 18597
rect 26555 18532 26556 18596
rect 26620 18532 26621 18596
rect 26555 18531 26621 18532
rect 25819 9620 25885 9621
rect 25819 9556 25820 9620
rect 25884 9556 25885 9620
rect 25819 9555 25885 9556
rect 25267 9212 25333 9213
rect 25267 9148 25268 9212
rect 25332 9148 25333 9212
rect 25267 9147 25333 9148
rect 26187 9212 26253 9213
rect 26187 9148 26188 9212
rect 26252 9148 26253 9212
rect 26187 9147 26253 9148
rect 25267 8396 25333 8397
rect 25267 8332 25268 8396
rect 25332 8332 25333 8396
rect 25267 8331 25333 8332
rect 25083 6084 25149 6085
rect 25083 6020 25084 6084
rect 25148 6020 25149 6084
rect 25083 6019 25149 6020
rect 24899 4180 24965 4181
rect 24899 4116 24900 4180
rect 24964 4116 24965 4180
rect 24899 4115 24965 4116
rect 24902 2549 24962 4115
rect 24899 2548 24965 2549
rect 24899 2484 24900 2548
rect 24964 2484 24965 2548
rect 24899 2483 24965 2484
rect 23795 1324 23861 1325
rect 23795 1260 23796 1324
rect 23860 1260 23861 1324
rect 23795 1259 23861 1260
rect 25270 917 25330 8331
rect 26190 7037 26250 9147
rect 26558 7717 26618 18531
rect 26742 18325 26802 34579
rect 27291 30564 27357 30565
rect 27291 30500 27292 30564
rect 27356 30500 27357 30564
rect 27291 30499 27357 30500
rect 27107 21180 27173 21181
rect 27107 21116 27108 21180
rect 27172 21116 27173 21180
rect 27107 21115 27173 21116
rect 26739 18324 26805 18325
rect 26739 18260 26740 18324
rect 26804 18260 26805 18324
rect 26739 18259 26805 18260
rect 26555 7716 26621 7717
rect 26555 7652 26556 7716
rect 26620 7652 26621 7716
rect 26555 7651 26621 7652
rect 26187 7036 26253 7037
rect 26187 6972 26188 7036
rect 26252 6972 26253 7036
rect 26187 6971 26253 6972
rect 27110 5949 27170 21115
rect 27294 19277 27354 30499
rect 27291 19276 27357 19277
rect 27291 19212 27292 19276
rect 27356 19212 27357 19276
rect 27291 19211 27357 19212
rect 27478 14653 27538 37843
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 28395 37500 28461 37501
rect 28395 37436 28396 37500
rect 28460 37436 28461 37500
rect 28395 37435 28461 37436
rect 27659 22132 27725 22133
rect 27659 22068 27660 22132
rect 27724 22068 27725 22132
rect 27659 22067 27725 22068
rect 27662 17917 27722 22067
rect 28398 20637 28458 37435
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 33179 29204 33245 29205
rect 33179 29140 33180 29204
rect 33244 29140 33245 29204
rect 33179 29139 33245 29140
rect 29315 25532 29381 25533
rect 29315 25468 29316 25532
rect 29380 25468 29381 25532
rect 29315 25467 29381 25468
rect 28395 20636 28461 20637
rect 28395 20572 28396 20636
rect 28460 20572 28461 20636
rect 28395 20571 28461 20572
rect 29131 20228 29197 20229
rect 29131 20164 29132 20228
rect 29196 20164 29197 20228
rect 29131 20163 29197 20164
rect 28947 19684 29013 19685
rect 28947 19620 28948 19684
rect 29012 19620 29013 19684
rect 28947 19619 29013 19620
rect 27843 19412 27909 19413
rect 27843 19348 27844 19412
rect 27908 19348 27909 19412
rect 27843 19347 27909 19348
rect 28579 19412 28645 19413
rect 28579 19348 28580 19412
rect 28644 19348 28645 19412
rect 28579 19347 28645 19348
rect 27659 17916 27725 17917
rect 27659 17852 27660 17916
rect 27724 17852 27725 17916
rect 27659 17851 27725 17852
rect 27659 17372 27725 17373
rect 27659 17308 27660 17372
rect 27724 17308 27725 17372
rect 27659 17307 27725 17308
rect 27475 14652 27541 14653
rect 27475 14588 27476 14652
rect 27540 14588 27541 14652
rect 27475 14587 27541 14588
rect 27662 12341 27722 17307
rect 27846 15197 27906 19347
rect 28027 18732 28093 18733
rect 28027 18668 28028 18732
rect 28092 18668 28093 18732
rect 28027 18667 28093 18668
rect 27843 15196 27909 15197
rect 27843 15132 27844 15196
rect 27908 15132 27909 15196
rect 27843 15131 27909 15132
rect 27659 12340 27725 12341
rect 27659 12276 27660 12340
rect 27724 12276 27725 12340
rect 27659 12275 27725 12276
rect 28030 5949 28090 18667
rect 27107 5948 27173 5949
rect 27107 5884 27108 5948
rect 27172 5884 27173 5948
rect 27107 5883 27173 5884
rect 28027 5948 28093 5949
rect 28027 5884 28028 5948
rect 28092 5884 28093 5948
rect 28027 5883 28093 5884
rect 27110 1053 27170 5883
rect 28582 2549 28642 19347
rect 28950 14381 29010 19619
rect 28947 14380 29013 14381
rect 28947 14316 28948 14380
rect 29012 14316 29013 14380
rect 28947 14315 29013 14316
rect 28947 14244 29013 14245
rect 28947 14180 28948 14244
rect 29012 14180 29013 14244
rect 28947 14179 29013 14180
rect 28950 10165 29010 14179
rect 29134 11797 29194 20163
rect 29318 14109 29378 25467
rect 32259 24852 32325 24853
rect 32259 24788 32260 24852
rect 32324 24788 32325 24852
rect 32259 24787 32325 24788
rect 30419 22404 30485 22405
rect 30419 22340 30420 22404
rect 30484 22340 30485 22404
rect 30419 22339 30485 22340
rect 30787 22404 30853 22405
rect 30787 22340 30788 22404
rect 30852 22340 30853 22404
rect 30787 22339 30853 22340
rect 31523 22404 31589 22405
rect 31523 22340 31524 22404
rect 31588 22340 31589 22404
rect 31523 22339 31589 22340
rect 30235 19548 30301 19549
rect 30235 19484 30236 19548
rect 30300 19484 30301 19548
rect 30235 19483 30301 19484
rect 30238 14925 30298 19483
rect 30422 15741 30482 22339
rect 30419 15740 30485 15741
rect 30419 15676 30420 15740
rect 30484 15676 30485 15740
rect 30419 15675 30485 15676
rect 30235 14924 30301 14925
rect 30235 14860 30236 14924
rect 30300 14860 30301 14924
rect 30235 14859 30301 14860
rect 29315 14108 29381 14109
rect 29315 14044 29316 14108
rect 29380 14044 29381 14108
rect 29315 14043 29381 14044
rect 29131 11796 29197 11797
rect 29131 11732 29132 11796
rect 29196 11732 29197 11796
rect 29131 11731 29197 11732
rect 30790 11117 30850 22339
rect 31339 19684 31405 19685
rect 31339 19620 31340 19684
rect 31404 19620 31405 19684
rect 31339 19619 31405 19620
rect 31342 11661 31402 19619
rect 31339 11660 31405 11661
rect 31339 11596 31340 11660
rect 31404 11596 31405 11660
rect 31339 11595 31405 11596
rect 30787 11116 30853 11117
rect 30787 11052 30788 11116
rect 30852 11052 30853 11116
rect 30787 11051 30853 11052
rect 31526 10301 31586 22339
rect 31891 21588 31957 21589
rect 31891 21524 31892 21588
rect 31956 21524 31957 21588
rect 31891 21523 31957 21524
rect 31707 12476 31773 12477
rect 31707 12412 31708 12476
rect 31772 12412 31773 12476
rect 31707 12411 31773 12412
rect 31710 12341 31770 12411
rect 31707 12340 31773 12341
rect 31707 12276 31708 12340
rect 31772 12276 31773 12340
rect 31707 12275 31773 12276
rect 31523 10300 31589 10301
rect 31523 10236 31524 10300
rect 31588 10236 31589 10300
rect 31523 10235 31589 10236
rect 28947 10164 29013 10165
rect 28947 10100 28948 10164
rect 29012 10100 29013 10164
rect 28947 10099 29013 10100
rect 31894 8261 31954 21523
rect 32075 19820 32141 19821
rect 32075 19756 32076 19820
rect 32140 19756 32141 19820
rect 32075 19755 32141 19756
rect 32078 9485 32138 19755
rect 32262 18325 32322 24787
rect 32259 18324 32325 18325
rect 32259 18260 32260 18324
rect 32324 18260 32325 18324
rect 32259 18259 32325 18260
rect 32443 18188 32509 18189
rect 32443 18124 32444 18188
rect 32508 18124 32509 18188
rect 32443 18123 32509 18124
rect 32075 9484 32141 9485
rect 32075 9420 32076 9484
rect 32140 9420 32141 9484
rect 32075 9419 32141 9420
rect 31891 8260 31957 8261
rect 31891 8196 31892 8260
rect 31956 8196 31957 8260
rect 31891 8195 31957 8196
rect 32446 6901 32506 18123
rect 32443 6900 32509 6901
rect 32443 6836 32444 6900
rect 32508 6836 32509 6900
rect 32443 6835 32509 6836
rect 33182 6357 33242 29139
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 33915 19684 33981 19685
rect 33915 19620 33916 19684
rect 33980 19620 33981 19684
rect 33915 19619 33981 19620
rect 33918 11525 33978 19619
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 33915 11524 33981 11525
rect 33915 11460 33916 11524
rect 33980 11460 33981 11524
rect 33915 11459 33981 11460
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 33179 6356 33245 6357
rect 33179 6292 33180 6356
rect 33244 6292 33245 6356
rect 33179 6291 33245 6292
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 28579 2548 28645 2549
rect 28579 2484 28580 2548
rect 28644 2484 28645 2548
rect 28579 2483 28645 2484
rect 34928 2128 35248 2688
rect 27107 1052 27173 1053
rect 27107 988 27108 1052
rect 27172 988 27173 1052
rect 27107 987 27173 988
rect 25267 916 25333 917
rect 25267 852 25268 916
rect 25332 852 25333 916
rect 25267 851 25333 852
rect 23427 780 23493 781
rect 23427 716 23428 780
rect 23492 716 23493 780
rect 23427 715 23493 716
rect 22139 100 22205 101
rect 22139 36 22140 100
rect 22204 36 22205 100
rect 22139 35 22205 36
use sky130_fd_sc_hd__diode_2  ANTENNA__0398__A PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14352 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0400__A
timestamp 1644511149
transform -1 0 1564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0401__A
timestamp 1644511149
transform 1 0 11960 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0407__A
timestamp 1644511149
transform 1 0 2024 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0408__A
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0415__A
timestamp 1644511149
transform 1 0 2024 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0416__A
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0416__B
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0416__C
timestamp 1644511149
transform 1 0 10856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0416__D
timestamp 1644511149
transform 1 0 16008 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0418__A
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0418__B
timestamp 1644511149
transform 1 0 4416 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0418__C
timestamp 1644511149
transform -1 0 4876 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0418__D
timestamp 1644511149
transform 1 0 3496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0420__A
timestamp 1644511149
transform -1 0 2760 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0420__B
timestamp 1644511149
transform -1 0 2392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0420__C
timestamp 1644511149
transform 1 0 3128 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0420__D
timestamp 1644511149
transform -1 0 2944 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0422__A
timestamp 1644511149
transform -1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0422__B
timestamp 1644511149
transform -1 0 24196 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0422__C
timestamp 1644511149
transform 1 0 17940 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0422__D
timestamp 1644511149
transform -1 0 20056 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0424__A
timestamp 1644511149
transform -1 0 2208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0424__B
timestamp 1644511149
transform -1 0 2760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0424__C
timestamp 1644511149
transform -1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0424__D
timestamp 1644511149
transform -1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0426__A
timestamp 1644511149
transform -1 0 23736 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0427__A
timestamp 1644511149
transform -1 0 8372 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0428__A
timestamp 1644511149
transform -1 0 6624 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0429__A
timestamp 1644511149
transform -1 0 5612 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0430__A
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0430__B
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0430__C
timestamp 1644511149
transform -1 0 24564 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0430__D
timestamp 1644511149
transform -1 0 25760 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0432__A
timestamp 1644511149
transform 1 0 10212 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0432__B
timestamp 1644511149
transform -1 0 8924 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0432__C
timestamp 1644511149
transform -1 0 9476 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0432__D
timestamp 1644511149
transform -1 0 6716 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0434__A
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0434__B
timestamp 1644511149
transform 1 0 2300 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0434__C
timestamp 1644511149
transform 1 0 3312 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0434__D
timestamp 1644511149
transform 1 0 2852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0436__A
timestamp 1644511149
transform -1 0 25116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0436__B
timestamp 1644511149
transform -1 0 26036 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0436__C
timestamp 1644511149
transform 1 0 20424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0436__D
timestamp 1644511149
transform 1 0 24104 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__A
timestamp 1644511149
transform -1 0 9108 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__B
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__C
timestamp 1644511149
transform 1 0 7176 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__D
timestamp 1644511149
transform 1 0 4140 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0440__A
timestamp 1644511149
transform -1 0 10028 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0441__A
timestamp 1644511149
transform -1 0 12696 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0442__A
timestamp 1644511149
transform 1 0 14720 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0443__A
timestamp 1644511149
transform -1 0 15456 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0444__A
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0444__B
timestamp 1644511149
transform -1 0 9292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0444__C
timestamp 1644511149
transform -1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0444__D
timestamp 1644511149
transform -1 0 10948 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__A
timestamp 1644511149
transform 1 0 4324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__B
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__C
timestamp 1644511149
transform 1 0 5428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__D
timestamp 1644511149
transform 1 0 4876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__A
timestamp 1644511149
transform 1 0 25484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__B
timestamp 1644511149
transform -1 0 26220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__C
timestamp 1644511149
transform -1 0 25852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__D
timestamp 1644511149
transform -1 0 26404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0450__A
timestamp 1644511149
transform -1 0 2208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0450__B
timestamp 1644511149
transform -1 0 1656 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0450__C
timestamp 1644511149
transform 1 0 2576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0450__D
timestamp 1644511149
transform 1 0 3128 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0451__A
timestamp 1644511149
transform -1 0 21160 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0452__A
timestamp 1644511149
transform -1 0 26956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0452__B
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0452__C
timestamp 1644511149
transform 1 0 24748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0452__D
timestamp 1644511149
transform 1 0 25668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__A
timestamp 1644511149
transform -1 0 26496 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0456__A
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__A
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__B
timestamp 1644511149
transform -1 0 27508 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__C
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__D
timestamp 1644511149
transform -1 0 25484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__A
timestamp 1644511149
transform -1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__B
timestamp 1644511149
transform 1 0 20608 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__C
timestamp 1644511149
transform 1 0 14628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__D
timestamp 1644511149
transform -1 0 14352 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0462__A
timestamp 1644511149
transform -1 0 23644 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0462__B
timestamp 1644511149
transform -1 0 25116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0462__C
timestamp 1644511149
transform 1 0 26404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0462__D
timestamp 1644511149
transform -1 0 19964 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__A
timestamp 1644511149
transform -1 0 26404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__B
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__C
timestamp 1644511149
transform -1 0 28060 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__D
timestamp 1644511149
transform 1 0 24932 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__A
timestamp 1644511149
transform -1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__B
timestamp 1644511149
transform -1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__C
timestamp 1644511149
transform -1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__D
timestamp 1644511149
transform -1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0467__A
timestamp 1644511149
transform -1 0 26036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__A
timestamp 1644511149
transform 1 0 6716 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0470__A
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__A
timestamp 1644511149
transform -1 0 7360 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__A
timestamp 1644511149
transform 1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__A
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__B
timestamp 1644511149
transform 1 0 3036 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__C
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__D
timestamp 1644511149
transform 1 0 2668 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__A
timestamp 1644511149
transform -1 0 2208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__B
timestamp 1644511149
transform -1 0 2760 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__C
timestamp 1644511149
transform -1 0 3404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__D
timestamp 1644511149
transform -1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__A
timestamp 1644511149
transform -1 0 21344 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__B
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__A
timestamp 1644511149
transform 1 0 22356 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__B
timestamp 1644511149
transform 1 0 23460 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0504__A
timestamp 1644511149
transform -1 0 24196 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0504__B
timestamp 1644511149
transform 1 0 24564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__A
timestamp 1644511149
transform -1 0 23460 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__B
timestamp 1644511149
transform 1 0 23920 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__A
timestamp 1644511149
transform 1 0 17572 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0511__A
timestamp 1644511149
transform -1 0 24472 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__A
timestamp 1644511149
transform -1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__A
timestamp 1644511149
transform -1 0 25024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__A
timestamp 1644511149
transform 1 0 21528 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__A
timestamp 1644511149
transform -1 0 24564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__A
timestamp 1644511149
transform 1 0 22080 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A
timestamp 1644511149
transform -1 0 28060 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__A
timestamp 1644511149
transform 1 0 22632 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__A
timestamp 1644511149
transform 1 0 29716 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__A
timestamp 1644511149
transform 1 0 23184 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__A
timestamp 1644511149
transform 1 0 30452 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__A
timestamp 1644511149
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__A
timestamp 1644511149
transform 1 0 32292 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__A_N
timestamp 1644511149
transform -1 0 26312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__B
timestamp 1644511149
transform 1 0 23092 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__A_N
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__B
timestamp 1644511149
transform 1 0 17572 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__A_N
timestamp 1644511149
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__B
timestamp 1644511149
transform 1 0 19044 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__A_N
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__B
timestamp 1644511149
transform 1 0 20884 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__B
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__A
timestamp 1644511149
transform 1 0 24932 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__B
timestamp 1644511149
transform 1 0 24656 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__B
timestamp 1644511149
transform -1 0 25668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__B
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__B
timestamp 1644511149
transform 1 0 26036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__A_N
timestamp 1644511149
transform -1 0 26956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__B
timestamp 1644511149
transform 1 0 27508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A_N
timestamp 1644511149
transform -1 0 28244 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__B
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A_N
timestamp 1644511149
transform -1 0 26220 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__B
timestamp 1644511149
transform 1 0 27324 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__A_N
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__B
timestamp 1644511149
transform -1 0 28244 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__A_N
timestamp 1644511149
transform -1 0 12236 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__B
timestamp 1644511149
transform 1 0 11040 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__A
timestamp 1644511149
transform -1 0 21988 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A_N
timestamp 1644511149
transform -1 0 13248 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__B
timestamp 1644511149
transform -1 0 10580 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__A
timestamp 1644511149
transform -1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__A_N
timestamp 1644511149
transform -1 0 23828 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__B
timestamp 1644511149
transform 1 0 18032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__A_N
timestamp 1644511149
transform 1 0 25208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__B
timestamp 1644511149
transform -1 0 25116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A_N
timestamp 1644511149
transform -1 0 14352 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B
timestamp 1644511149
transform -1 0 16008 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__A
timestamp 1644511149
transform -1 0 21344 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__B
timestamp 1644511149
transform -1 0 21620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__B
timestamp 1644511149
transform -1 0 25944 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__B
timestamp 1644511149
transform -1 0 22172 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__A
timestamp 1644511149
transform -1 0 26128 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__A_N
timestamp 1644511149
transform -1 0 16376 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__B
timestamp 1644511149
transform 1 0 15456 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A
timestamp 1644511149
transform -1 0 23828 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A_N
timestamp 1644511149
transform 1 0 15180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__A
timestamp 1644511149
transform 1 0 22448 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__A_N
timestamp 1644511149
transform 1 0 16744 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A
timestamp 1644511149
transform 1 0 23000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__A_N
timestamp 1644511149
transform 1 0 17020 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A
timestamp 1644511149
transform -1 0 24288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__A_N
timestamp 1644511149
transform 1 0 17572 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__B
timestamp 1644511149
transform 1 0 18584 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__A
timestamp 1644511149
transform -1 0 25852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A_N
timestamp 1644511149
transform -1 0 22724 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__A
timestamp 1644511149
transform 1 0 26956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__A_N
timestamp 1644511149
transform 1 0 16652 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__B
timestamp 1644511149
transform 1 0 22632 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A
timestamp 1644511149
transform -1 0 6808 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A0
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__S
timestamp 1644511149
transform 1 0 11684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__A0
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__S
timestamp 1644511149
transform 1 0 12328 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A0
timestamp 1644511149
transform 1 0 12880 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__S
timestamp 1644511149
transform 1 0 14720 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__A
timestamp 1644511149
transform -1 0 5888 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__A0
timestamp 1644511149
transform 1 0 13432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__S
timestamp 1644511149
transform 1 0 15732 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A0
timestamp 1644511149
transform 1 0 15272 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__S
timestamp 1644511149
transform 1 0 15824 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__A
timestamp 1644511149
transform -1 0 9660 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__A0
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__B
timestamp 1644511149
transform -1 0 23368 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__A0
timestamp 1644511149
transform 1 0 15456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__A_N
timestamp 1644511149
transform 1 0 23184 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__B
timestamp 1644511149
transform 1 0 23736 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A0
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__S
timestamp 1644511149
transform -1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A0
timestamp 1644511149
transform 1 0 17204 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__S
timestamp 1644511149
transform -1 0 17112 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A0
timestamp 1644511149
transform 1 0 17480 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__S
timestamp 1644511149
transform -1 0 16836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A0
timestamp 1644511149
transform -1 0 23920 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__S
timestamp 1644511149
transform -1 0 18216 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__A0
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__S
timestamp 1644511149
transform -1 0 18768 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__A0
timestamp 1644511149
transform -1 0 25760 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__A1
timestamp 1644511149
transform 1 0 24472 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__S
timestamp 1644511149
transform -1 0 25208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__A_N
timestamp 1644511149
transform -1 0 16284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__S
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A
timestamp 1644511149
transform -1 0 23460 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__S
timestamp 1644511149
transform -1 0 11316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__A
timestamp 1644511149
transform -1 0 18308 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__S
timestamp 1644511149
transform -1 0 12788 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__A
timestamp 1644511149
transform -1 0 21436 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__S
timestamp 1644511149
transform -1 0 13340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A
timestamp 1644511149
transform 1 0 21988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A
timestamp 1644511149
transform -1 0 22172 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__A
timestamp 1644511149
transform -1 0 27140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A
timestamp 1644511149
transform -1 0 27692 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A1
timestamp 1644511149
transform 1 0 17204 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A
timestamp 1644511149
transform -1 0 26680 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__S
timestamp 1644511149
transform -1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A
timestamp 1644511149
transform 1 0 27508 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__S
timestamp 1644511149
transform -1 0 19412 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A
timestamp 1644511149
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__S
timestamp 1644511149
transform -1 0 19964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A
timestamp 1644511149
transform 1 0 29716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__S
timestamp 1644511149
transform 1 0 25024 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A
timestamp 1644511149
transform 1 0 31188 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A_N
timestamp 1644511149
transform -1 0 25760 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B
timestamp 1644511149
transform 1 0 25576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A
timestamp 1644511149
transform -1 0 6992 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__B
timestamp 1644511149
transform 1 0 20700 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A_N
timestamp 1644511149
transform -1 0 26312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__B
timestamp 1644511149
transform -1 0 25300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A_N
timestamp 1644511149
transform -1 0 17388 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A
timestamp 1644511149
transform -1 0 13892 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__B
timestamp 1644511149
transform -1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__D
timestamp 1644511149
transform -1 0 14444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 1644511149
transform 1 0 10396 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__D
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__C
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1644511149
transform 1 0 25668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1644511149
transform 1 0 28612 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__B
timestamp 1644511149
transform 1 0 27876 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__C
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1644511149
transform -1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 1644511149
transform 1 0 26036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A1
timestamp 1644511149
transform 1 0 27508 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B1
timestamp 1644511149
transform 1 0 27508 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A1
timestamp 1644511149
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__B1
timestamp 1644511149
transform 1 0 27140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1644511149
transform -1 0 16836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__B
timestamp 1644511149
transform 1 0 18308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1644511149
transform -1 0 4508 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A
timestamp 1644511149
transform -1 0 15364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__B
timestamp 1644511149
transform 1 0 15364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A
timestamp 1644511149
transform -1 0 5060 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1644511149
transform -1 0 16100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__B
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1644511149
transform -1 0 4784 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A
timestamp 1644511149
transform -1 0 14996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__B
timestamp 1644511149
transform 1 0 17756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A
timestamp 1644511149
transform 1 0 26128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__B
timestamp 1644511149
transform 1 0 24932 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A
timestamp 1644511149
transform -1 0 11776 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__B
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B
timestamp 1644511149
transform 1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B
timestamp 1644511149
transform -1 0 26312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1644511149
transform 1 0 24288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__B
timestamp 1644511149
transform 1 0 24840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A
timestamp 1644511149
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A1
timestamp 1644511149
transform -1 0 26864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B1
timestamp 1644511149
transform 1 0 27508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A
timestamp 1644511149
transform -1 0 28244 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__B
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A
timestamp 1644511149
transform -1 0 3956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A1
timestamp 1644511149
transform -1 0 25668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B1
timestamp 1644511149
transform -1 0 26496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A1
timestamp 1644511149
transform -1 0 27416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A1
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1644511149
transform -1 0 27876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1644511149
transform 1 0 9016 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1644511149
transform 1 0 27508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B
timestamp 1644511149
transform -1 0 28796 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A1
timestamp 1644511149
transform -1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A1
timestamp 1644511149
transform -1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A2
timestamp 1644511149
transform -1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B1
timestamp 1644511149
transform -1 0 8648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A1
timestamp 1644511149
transform -1 0 27324 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A2
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B
timestamp 1644511149
transform -1 0 11684 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A1
timestamp 1644511149
transform -1 0 10488 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A2
timestamp 1644511149
transform -1 0 12328 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1644511149
transform -1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B
timestamp 1644511149
transform -1 0 9292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__C
timestamp 1644511149
transform -1 0 7912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A
timestamp 1644511149
transform -1 0 11868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__C
timestamp 1644511149
transform -1 0 28244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A
timestamp 1644511149
transform -1 0 29716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A2
timestamp 1644511149
transform -1 0 29348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__B
timestamp 1644511149
transform -1 0 12236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B
timestamp 1644511149
transform -1 0 8096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A2
timestamp 1644511149
transform 1 0 28612 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A1
timestamp 1644511149
transform -1 0 6348 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A2
timestamp 1644511149
transform -1 0 7360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B1
timestamp 1644511149
transform -1 0 6808 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A1
timestamp 1644511149
transform 1 0 28244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A2
timestamp 1644511149
transform 1 0 27508 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__B
timestamp 1644511149
transform -1 0 29900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A1
timestamp 1644511149
transform -1 0 30452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A2
timestamp 1644511149
transform -1 0 29716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1644511149
transform 1 0 5612 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__B
timestamp 1644511149
transform -1 0 6808 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__C
timestamp 1644511149
transform -1 0 5244 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1644511149
transform -1 0 13524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__B
timestamp 1644511149
transform -1 0 14904 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2
timestamp 1644511149
transform -1 0 28244 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A
timestamp 1644511149
transform -1 0 29348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B
timestamp 1644511149
transform -1 0 30268 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A
timestamp 1644511149
transform 1 0 4324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__B
timestamp 1644511149
transform 1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1
timestamp 1644511149
transform -1 0 10120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1644511149
transform -1 0 2944 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1644511149
transform -1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__C
timestamp 1644511149
transform -1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A
timestamp 1644511149
transform -1 0 2208 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A2
timestamp 1644511149
transform -1 0 17388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B
timestamp 1644511149
transform 1 0 19412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 1644511149
transform -1 0 28980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B
timestamp 1644511149
transform -1 0 27968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1
timestamp 1644511149
transform -1 0 13340 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A2
timestamp 1644511149
transform -1 0 12880 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B1
timestamp 1644511149
transform -1 0 14260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A1
timestamp 1644511149
transform -1 0 28796 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A2
timestamp 1644511149
transform -1 0 28520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A
timestamp 1644511149
transform -1 0 29348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__B
timestamp 1644511149
transform -1 0 28244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__C
timestamp 1644511149
transform -1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A1
timestamp 1644511149
transform -1 0 13892 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A2
timestamp 1644511149
transform -1 0 13432 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B1
timestamp 1644511149
transform -1 0 14812 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A
timestamp 1644511149
transform 1 0 15732 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B
timestamp 1644511149
transform -1 0 19412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A2
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B1
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A2
timestamp 1644511149
transform -1 0 29900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A2
timestamp 1644511149
transform 1 0 27140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A
timestamp 1644511149
transform -1 0 14444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B
timestamp 1644511149
transform -1 0 15364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A1
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A2
timestamp 1644511149
transform -1 0 30268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__B1
timestamp 1644511149
transform -1 0 29900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A1
timestamp 1644511149
transform 1 0 27508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A2
timestamp 1644511149
transform 1 0 28612 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A1
timestamp 1644511149
transform -1 0 30820 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A
timestamp 1644511149
transform -1 0 20148 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B
timestamp 1644511149
transform -1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A
timestamp 1644511149
transform -1 0 9936 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A
timestamp 1644511149
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A0
timestamp 1644511149
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A_N
timestamp 1644511149
transform 1 0 5152 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A
timestamp 1644511149
transform -1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A1
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A1
timestamp 1644511149
transform 1 0 4784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A
timestamp 1644511149
transform -1 0 4232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A1
timestamp 1644511149
transform -1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A
timestamp 1644511149
transform -1 0 6900 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A1
timestamp 1644511149
transform 1 0 4600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A_N
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A1
timestamp 1644511149
transform 1 0 5704 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A_N
timestamp 1644511149
transform 1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A1
timestamp 1644511149
transform -1 0 31004 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A_N
timestamp 1644511149
transform -1 0 7360 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A1
timestamp 1644511149
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A_N
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A
timestamp 1644511149
transform -1 0 22540 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A1
timestamp 1644511149
transform -1 0 15916 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__S
timestamp 1644511149
transform 1 0 28060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A_N
timestamp 1644511149
transform -1 0 29900 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A
timestamp 1644511149
transform -1 0 29716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A1
timestamp 1644511149
transform 1 0 2392 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__S
timestamp 1644511149
transform -1 0 3128 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A_N
timestamp 1644511149
transform -1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B
timestamp 1644511149
transform -1 0 21988 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A0
timestamp 1644511149
transform -1 0 29348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A1
timestamp 1644511149
transform -1 0 28244 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__S
timestamp 1644511149
transform -1 0 28796 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A_N
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A1
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__S
timestamp 1644511149
transform 1 0 16836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A_N
timestamp 1644511149
transform -1 0 30268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A0
timestamp 1644511149
transform -1 0 16836 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A1
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__S
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A_N
timestamp 1644511149
transform -1 0 13064 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 1644511149
transform -1 0 23276 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A1
timestamp 1644511149
transform 1 0 2392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__S
timestamp 1644511149
transform 1 0 2944 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A_N
timestamp 1644511149
transform 1 0 28612 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B
timestamp 1644511149
transform -1 0 29716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A
timestamp 1644511149
transform -1 0 8464 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A0
timestamp 1644511149
transform -1 0 17388 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A1
timestamp 1644511149
transform 1 0 18676 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__S
timestamp 1644511149
transform 1 0 19228 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A_N
timestamp 1644511149
transform -1 0 29900 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A
timestamp 1644511149
transform -1 0 11040 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A0
timestamp 1644511149
transform -1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__S
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A_N
timestamp 1644511149
transform 1 0 9200 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A1
timestamp 1644511149
transform -1 0 10488 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__S
timestamp 1644511149
transform -1 0 11592 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A_N
timestamp 1644511149
transform 1 0 12052 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A0
timestamp 1644511149
transform -1 0 21344 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A1
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__S
timestamp 1644511149
transform -1 0 23828 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A_N
timestamp 1644511149
transform 1 0 11960 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A
timestamp 1644511149
transform 1 0 7636 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A0
timestamp 1644511149
transform -1 0 14260 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A1
timestamp 1644511149
transform -1 0 14996 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A_N
timestamp 1644511149
transform -1 0 9752 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A
timestamp 1644511149
transform 1 0 5152 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A0
timestamp 1644511149
transform 1 0 3496 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A1
timestamp 1644511149
transform 1 0 4048 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A0
timestamp 1644511149
transform 1 0 2852 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A0
timestamp 1644511149
transform 1 0 3404 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1644511149
transform -1 0 7728 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A0
timestamp 1644511149
transform 1 0 6072 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A0
timestamp 1644511149
transform 1 0 6992 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A0
timestamp 1644511149
transform 1 0 8004 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A0
timestamp 1644511149
transform 1 0 4324 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A0
timestamp 1644511149
transform 1 0 5520 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__S
timestamp 1644511149
transform -1 0 5888 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A0
timestamp 1644511149
transform 1 0 12512 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__S
timestamp 1644511149
transform -1 0 13616 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A_N
timestamp 1644511149
transform -1 0 30452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__D
timestamp 1644511149
transform -1 0 29716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__D
timestamp 1644511149
transform -1 0 8740 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1644511149
transform -1 0 19964 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1644511149
transform -1 0 23644 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1644511149
transform -1 0 26404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1644511149
transform 1 0 28244 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A
timestamp 1644511149
transform 1 0 29716 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1644511149
transform 1 0 25116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A
timestamp 1644511149
transform 1 0 27692 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A
timestamp 1644511149
transform -1 0 27324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1644511149
transform -1 0 28336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1644511149
transform -1 0 28244 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1644511149
transform 1 0 30084 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A
timestamp 1644511149
transform -1 0 32200 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1644511149
transform -1 0 33672 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1644511149
transform 1 0 34868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A
timestamp 1644511149
transform -1 0 24564 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A
timestamp 1644511149
transform -1 0 29716 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A
timestamp 1644511149
transform -1 0 31556 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1644511149
transform -1 0 24196 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1644511149
transform 1 0 32384 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A
timestamp 1644511149
transform 1 0 35604 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A
timestamp 1644511149
transform -1 0 11040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1644511149
transform -1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1644511149
transform -1 0 30268 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A
timestamp 1644511149
transform -1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A
timestamp 1644511149
transform -1 0 5888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1644511149
transform -1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1644511149
transform -1 0 30820 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1644511149
transform -1 0 30452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1644511149
transform -1 0 11684 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1644511149
transform -1 0 14812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A
timestamp 1644511149
transform -1 0 12236 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1644511149
transform -1 0 9108 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A
timestamp 1644511149
transform -1 0 8464 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A
timestamp 1644511149
transform -1 0 8924 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1644511149
transform -1 0 11040 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A
timestamp 1644511149
transform -1 0 14168 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1644511149
transform -1 0 15548 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A
timestamp 1644511149
transform -1 0 11224 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1644511149
transform -1 0 13248 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_A
timestamp 1644511149
transform -1 0 2852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_A
timestamp 1644511149
transform -1 0 12788 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_A
timestamp 1644511149
transform -1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_A
timestamp 1644511149
transform -1 0 16100 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 23276 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 25116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 2760 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 2116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 2668 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 3312 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 4140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 5060 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 3956 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 1564 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 2116 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 4140 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 2208 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 1564 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 2208 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 2208 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 2208 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 2208 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 2208 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 2208 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 1564 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1644511149
transform -1 0 2760 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1644511149
transform -1 0 22540 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1644511149
transform -1 0 4232 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1644511149
transform -1 0 2116 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1644511149
transform -1 0 23092 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1644511149
transform -1 0 24840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1644511149
transform -1 0 24564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1644511149
transform -1 0 25576 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1644511149
transform -1 0 26128 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1644511149
transform -1 0 25668 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1644511149
transform -1 0 23644 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1644511149
transform -1 0 24196 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1644511149
transform -1 0 25116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1644511149
transform -1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1644511149
transform -1 0 37536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1644511149
transform -1 0 38916 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1644511149
transform -1 0 39836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1644511149
transform -1 0 40756 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1644511149
transform -1 0 41952 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1644511149
transform -1 0 43516 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1644511149
transform -1 0 42780 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1644511149
transform -1 0 41952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1644511149
transform -1 0 43516 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1644511149
transform -1 0 29532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1644511149
transform -1 0 30820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1644511149
transform -1 0 34132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1644511149
transform -1 0 33212 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1644511149
transform -1 0 34684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1644511149
transform -1 0 35420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1644511149
transform -1 0 36156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1644511149
transform -1 0 37444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1644511149
transform -1 0 37996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1644511149
transform -1 0 28796 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1644511149
transform -1 0 38732 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1644511149
transform -1 0 40388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1644511149
transform -1 0 40940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1644511149
transform -1 0 41492 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1644511149
transform -1 0 42780 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1644511149
transform -1 0 42228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1644511149
transform -1 0 43700 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1644511149
transform -1 0 44252 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1644511149
transform -1 0 42964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1644511149
transform -1 0 30084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1644511149
transform -1 0 31372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1644511149
transform -1 0 32476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1644511149
transform -1 0 33764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1644511149
transform -1 0 33948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1644511149
transform -1 0 34868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1644511149
transform -1 0 35420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1644511149
transform -1 0 36708 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1644511149
transform -1 0 37352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1644511149
transform -1 0 25852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1644511149
transform -1 0 23828 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1644511149
transform -1 0 26404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1644511149
transform -1 0 24748 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1644511149
transform -1 0 24564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1644511149
transform -1 0 25668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1644511149
transform -1 0 25300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1644511149
transform -1 0 26220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1644511149
transform -1 0 27324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1644511149
transform -1 0 27876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1644511149
transform -1 0 25852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1644511149
transform -1 0 24196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1644511149
transform -1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1644511149
transform -1 0 26772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1644511149
transform -1 0 24748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1644511149
transform -1 0 26404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1644511149
transform -1 0 25668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1644511149
transform -1 0 25300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1644511149
transform -1 0 26220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1644511149
transform -1 0 25852 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1644511149
transform -1 0 27140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1644511149
transform -1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1644511149
transform -1 0 25208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1644511149
transform -1 0 26772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1644511149
transform -1 0 27692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1644511149
transform -1 0 25760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1644511149
transform -1 0 26404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1644511149
transform -1 0 28152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1644511149
transform -1 0 5428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1644511149
transform -1 0 18400 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1644511149
transform -1 0 20148 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1644511149
transform -1 0 19964 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1644511149
transform -1 0 20700 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1644511149
transform -1 0 20516 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1644511149
transform -1 0 21252 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1644511149
transform -1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1644511149
transform -1 0 21988 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1644511149
transform -1 0 3128 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1644511149
transform -1 0 11040 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1644511149
transform -1 0 13616 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1644511149
transform -1 0 16192 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1644511149
transform -1 0 16836 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1644511149
transform -1 0 17204 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1644511149
transform -1 0 19228 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1644511149
transform -1 0 19780 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1644511149
transform -1 0 20884 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1644511149
transform -1 0 22172 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 1644511149
transform -1 0 23736 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 1644511149
transform -1 0 2852 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 1644511149
transform -1 0 24748 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 1644511149
transform -1 0 26128 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 1644511149
transform -1 0 28152 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 1644511149
transform -1 0 28980 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 1644511149
transform -1 0 31556 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 1644511149
transform -1 0 30636 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 1644511149
transform -1 0 34132 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 1644511149
transform -1 0 33212 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 1644511149
transform -1 0 36708 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 1644511149
transform -1 0 35880 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 1644511149
transform -1 0 3680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 1644511149
transform -1 0 37260 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 1644511149
transform -1 0 38916 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input136_A
timestamp 1644511149
transform -1 0 40204 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input137_A
timestamp 1644511149
transform -1 0 41860 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input138_A
timestamp 1644511149
transform -1 0 41400 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input139_A
timestamp 1644511149
transform -1 0 5152 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input140_A
timestamp 1644511149
transform -1 0 5060 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input141_A
timestamp 1644511149
transform -1 0 8372 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input142_A
timestamp 1644511149
transform -1 0 8004 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input143_A
timestamp 1644511149
transform -1 0 9844 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input144_A
timestamp 1644511149
transform -1 0 10396 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input145_A
timestamp 1644511149
transform -1 0 11500 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input146_A
timestamp 1644511149
transform -1 0 5336 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input147_A
timestamp 1644511149
transform -1 0 4784 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input148_A
timestamp 1644511149
transform -1 0 20700 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input149_A
timestamp 1644511149
transform -1 0 21620 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input150_A
timestamp 1644511149
transform -1 0 22540 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input151_A
timestamp 1644511149
transform -1 0 21252 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input152_A
timestamp 1644511149
transform -1 0 22172 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input153_A
timestamp 1644511149
transform -1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input154_A
timestamp 1644511149
transform -1 0 23092 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input155_A
timestamp 1644511149
transform -1 0 22724 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input156_A
timestamp 1644511149
transform -1 0 25300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input157_A
timestamp 1644511149
transform -1 0 23644 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input158_A
timestamp 1644511149
transform -1 0 21620 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input159_A
timestamp 1644511149
transform -1 0 22540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input160_A
timestamp 1644511149
transform -1 0 23276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input161_A
timestamp 1644511149
transform -1 0 24196 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input162_A
timestamp 1644511149
transform -1 0 22172 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input163_A
timestamp 1644511149
transform -1 0 23092 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input164_A
timestamp 1644511149
transform -1 0 23828 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input165_A
timestamp 1644511149
transform -1 0 24748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input166_A
timestamp 1644511149
transform -1 0 22724 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input167_A
timestamp 1644511149
transform -1 0 25852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input168_A
timestamp 1644511149
transform -1 0 23644 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input169_A
timestamp 1644511149
transform -1 0 24564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input170_A
timestamp 1644511149
transform -1 0 25300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output171_A
timestamp 1644511149
transform -1 0 28980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output172_A
timestamp 1644511149
transform 1 0 37904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output173_A
timestamp 1644511149
transform -1 0 39284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1644511149
transform -1 0 40020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output175_A
timestamp 1644511149
transform 1 0 40756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output176_A
timestamp 1644511149
transform 1 0 41400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output177_A
timestamp 1644511149
transform 1 0 42136 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output178_A
timestamp 1644511149
transform 1 0 42964 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output179_A
timestamp 1644511149
transform 1 0 41584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output180_A
timestamp 1644511149
transform 1 0 43700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output188_A
timestamp 1644511149
transform -1 0 35972 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output189_A
timestamp 1644511149
transform 1 0 36432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output190_A
timestamp 1644511149
transform -1 0 27324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output191_A
timestamp 1644511149
transform -1 0 28244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output207_A
timestamp 1644511149
transform -1 0 27876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output209_A
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output211_A
timestamp 1644511149
transform 1 0 14352 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output217_A
timestamp 1644511149
transform 1 0 22540 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output218_A
timestamp 1644511149
transform 1 0 23092 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output219_A
timestamp 1644511149
transform -1 0 23828 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output221_A
timestamp 1644511149
transform -1 0 25300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output222_A
timestamp 1644511149
transform 1 0 25852 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output223_A
timestamp 1644511149
transform 1 0 27048 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output224_A
timestamp 1644511149
transform 1 0 28428 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output225_A
timestamp 1644511149
transform 1 0 29532 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output226_A
timestamp 1644511149
transform 1 0 31004 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output227_A
timestamp 1644511149
transform 1 0 32016 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output228_A
timestamp 1644511149
transform 1 0 33488 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output229_A
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output230_A
timestamp 1644511149
transform -1 0 36432 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output231_A
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output232_A
timestamp 1644511149
transform 1 0 37812 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output233_A
timestamp 1644511149
transform 1 0 38456 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output234_A
timestamp 1644511149
transform 1 0 39192 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output235_A
timestamp 1644511149
transform -1 0 40756 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output236_A
timestamp 1644511149
transform 1 0 42228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output237_A
timestamp 1644511149
transform 1 0 42964 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output238_A
timestamp 1644511149
transform 1 0 43332 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output239_A
timestamp 1644511149
transform 1 0 43700 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output241_A
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output243_A
timestamp 1644511149
transform 1 0 8280 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output244_A
timestamp 1644511149
transform 1 0 9476 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output245_A
timestamp 1644511149
transform 1 0 11868 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output246_A
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output247_A
timestamp 1644511149
transform 1 0 3128 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output255_A
timestamp 1644511149
transform 1 0 21988 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output256_A
timestamp 1644511149
transform 1 0 23184 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output257_A
timestamp 1644511149
transform -1 0 24564 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output258_A
timestamp 1644511149
transform 1 0 4324 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output259_A
timestamp 1644511149
transform 1 0 25024 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output260_A
timestamp 1644511149
transform 1 0 26312 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output261_A
timestamp 1644511149
transform 1 0 27600 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output262_A
timestamp 1644511149
transform -1 0 30268 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output263_A
timestamp 1644511149
transform 1 0 30268 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output264_A
timestamp 1644511149
transform 1 0 31096 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output265_A
timestamp 1644511149
transform 1 0 32660 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output266_A
timestamp 1644511149
transform 1 0 33580 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output267_A
timestamp 1644511149
transform 1 0 34868 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output268_A
timestamp 1644511149
transform 1 0 36248 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output269_A
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output270_A
timestamp 1644511149
transform 1 0 37812 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output271_A
timestamp 1644511149
transform 1 0 38548 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output272_A
timestamp 1644511149
transform -1 0 40020 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output273_A
timestamp 1644511149
transform 1 0 40756 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output274_A
timestamp 1644511149
transform -1 0 42596 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output275_A
timestamp 1644511149
transform 1 0 42964 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output276_A
timestamp 1644511149
transform 1 0 43700 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output277_A
timestamp 1644511149
transform 1 0 43700 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output281_A
timestamp 1644511149
transform 1 0 10028 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output282_A
timestamp 1644511149
transform 1 0 10764 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output283_A
timestamp 1644511149
transform 1 0 10856 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output284_A
timestamp 1644511149
transform 1 0 13156 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output285_A
timestamp 1644511149
transform 1 0 43332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output286_A
timestamp 1644511149
transform 1 0 43332 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44
timestamp 1644511149
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1644511149
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76
timestamp 1644511149
transform 1 0 8096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1644511149
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1644511149
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129
timestamp 1644511149
transform 1 0 12972 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1644511149
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_190
timestamp 1644511149
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201
timestamp 1644511149
transform 1 0 19596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_206
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1644511149
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_229
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1644511149
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_263
timestamp 1644511149
transform 1 0 25300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_271
timestamp 1644511149
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1644511149
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_319
timestamp 1644511149
transform 1 0 30452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1644511149
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_345
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_353
timestamp 1644511149
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1644511149
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1644511149
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_369
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1644511149
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_404
timestamp 1644511149
transform 1 0 38272 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_410
timestamp 1644511149
transform 1 0 38824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1644511149
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1644511149
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_425
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_435
timestamp 1644511149
transform 1 0 41124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_443
timestamp 1644511149
transform 1 0 41860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1644511149
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1644511149
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_465
timestamp 1644511149
transform 1 0 43884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1644511149
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_47
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1644511149
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1644511149
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_92
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1644511149
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1644511149
transform 1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1644511149
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1644511149
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_138
timestamp 1644511149
transform 1 0 13800 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_147
timestamp 1644511149
transform 1 0 14628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_154
timestamp 1644511149
transform 1 0 15272 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_160
timestamp 1644511149
transform 1 0 15824 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_175
timestamp 1644511149
transform 1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_182
timestamp 1644511149
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1644511149
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_196
timestamp 1644511149
transform 1 0 19136 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_204
timestamp 1644511149
transform 1 0 19872 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_208
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1644511149
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_229
timestamp 1644511149
transform 1 0 22172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_235
timestamp 1644511149
transform 1 0 22724 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_239
timestamp 1644511149
transform 1 0 23092 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_245
timestamp 1644511149
transform 1 0 23644 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1644511149
transform 1 0 24840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_266
timestamp 1644511149
transform 1 0 25576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1644511149
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_283
timestamp 1644511149
transform 1 0 27140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_291
timestamp 1644511149
transform 1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1644511149
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_311
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_319
timestamp 1644511149
transform 1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_327
timestamp 1644511149
transform 1 0 31188 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_345
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_353
timestamp 1644511149
transform 1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_369
timestamp 1644511149
transform 1 0 35052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_377
timestamp 1644511149
transform 1 0 35788 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1644511149
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_397
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_413
timestamp 1644511149
transform 1 0 39100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_421
timestamp 1644511149
transform 1 0 39836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_429
timestamp 1644511149
transform 1 0 40572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_437
timestamp 1644511149
transform 1 0 41308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_441
timestamp 1644511149
transform 1 0 41676 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1644511149
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_457
timestamp 1644511149
transform 1 0 43148 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_469
timestamp 1644511149
transform 1 0 44252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_39
timestamp 1644511149
transform 1 0 4692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_47
timestamp 1644511149
transform 1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_54
timestamp 1644511149
transform 1 0 6072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1644511149
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_92
timestamp 1644511149
transform 1 0 9568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_98
timestamp 1644511149
transform 1 0 10120 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_102
timestamp 1644511149
transform 1 0 10488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1644511149
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_113
timestamp 1644511149
transform 1 0 11500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_120
timestamp 1644511149
transform 1 0 12144 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1644511149
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_150
timestamp 1644511149
transform 1 0 14904 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_156
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_160
timestamp 1644511149
transform 1 0 15824 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_171
timestamp 1644511149
transform 1 0 16836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1644511149
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_208
timestamp 1644511149
transform 1 0 20240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_212
timestamp 1644511149
transform 1 0 20608 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_218
timestamp 1644511149
transform 1 0 21160 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_222
timestamp 1644511149
transform 1 0 21528 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_228
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_232
timestamp 1644511149
transform 1 0 22448 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_243
timestamp 1644511149
transform 1 0 23460 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_256
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_263
timestamp 1644511149
transform 1 0 25300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_269
timestamp 1644511149
transform 1 0 25852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_285
timestamp 1644511149
transform 1 0 27324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1644511149
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1644511149
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_313
timestamp 1644511149
transform 1 0 29900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_329
timestamp 1644511149
transform 1 0 31372 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_339
timestamp 1644511149
transform 1 0 32292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_350
timestamp 1644511149
transform 1 0 33304 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_370
timestamp 1644511149
transform 1 0 35144 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_380
timestamp 1644511149
transform 1 0 36064 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_390
timestamp 1644511149
transform 1 0 36984 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_398
timestamp 1644511149
transform 1 0 37720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_406
timestamp 1644511149
transform 1 0 38456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_414
timestamp 1644511149
transform 1 0 39192 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_425
timestamp 1644511149
transform 1 0 40204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_431
timestamp 1644511149
transform 1 0 40756 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_439
timestamp 1644511149
transform 1 0 41492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_444
timestamp 1644511149
transform 1 0 41952 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_452
timestamp 1644511149
transform 1 0 42688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_456
timestamp 1644511149
transform 1 0 43056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_461
timestamp 1644511149
transform 1 0 43516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_33
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_37
timestamp 1644511149
transform 1 0 4508 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1644511149
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_46
timestamp 1644511149
transform 1 0 5336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1644511149
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_68
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_75
timestamp 1644511149
transform 1 0 8004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_82
timestamp 1644511149
transform 1 0 8648 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_92
timestamp 1644511149
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_98
timestamp 1644511149
transform 1 0 10120 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1644511149
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1644511149
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_121
timestamp 1644511149
transform 1 0 12236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1644511149
transform 1 0 12788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_133
timestamp 1644511149
transform 1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1644511149
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1644511149
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1644511149
transform 1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_157
timestamp 1644511149
transform 1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1644511149
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_171
timestamp 1644511149
transform 1 0 16836 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_179
timestamp 1644511149
transform 1 0 17572 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_187
timestamp 1644511149
transform 1 0 18308 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_191
timestamp 1644511149
transform 1 0 18676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_197
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1644511149
transform 1 0 19596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1644511149
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1644511149
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1644511149
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_227
timestamp 1644511149
transform 1 0 21988 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_233
timestamp 1644511149
transform 1 0 22540 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_239
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_245
timestamp 1644511149
transform 1 0 23644 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_251
timestamp 1644511149
transform 1 0 24196 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_257
timestamp 1644511149
transform 1 0 24748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_263
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_269
timestamp 1644511149
transform 1 0 25852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1644511149
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_288
timestamp 1644511149
transform 1 0 27600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_294
timestamp 1644511149
transform 1 0 28152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_298
timestamp 1644511149
transform 1 0 28520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_301
timestamp 1644511149
transform 1 0 28796 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_309
timestamp 1644511149
transform 1 0 29532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_315
timestamp 1644511149
transform 1 0 30084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_323
timestamp 1644511149
transform 1 0 30820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_341
timestamp 1644511149
transform 1 0 32476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_355
timestamp 1644511149
transform 1 0 33764 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_365
timestamp 1644511149
transform 1 0 34684 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_381
timestamp 1644511149
transform 1 0 36156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1644511149
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_395
timestamp 1644511149
transform 1 0 37444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_401
timestamp 1644511149
transform 1 0 37996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_411
timestamp 1644511149
transform 1 0 38916 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_421
timestamp 1644511149
transform 1 0 39836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_427
timestamp 1644511149
transform 1 0 40388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_433
timestamp 1644511149
transform 1 0 40940 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_444
timestamp 1644511149
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_453
timestamp 1644511149
transform 1 0 42780 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_469
timestamp 1644511149
transform 1 0 44252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_6
timestamp 1644511149
transform 1 0 1656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1644511149
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1644511149
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_31
timestamp 1644511149
transform 1 0 3956 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1644511149
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1644511149
transform 1 0 5244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_57
timestamp 1644511149
transform 1 0 6348 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1644511149
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_69
timestamp 1644511149
transform 1 0 7452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1644511149
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_89
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_95
timestamp 1644511149
transform 1 0 9844 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_103
timestamp 1644511149
transform 1 0 10580 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_111
timestamp 1644511149
transform 1 0 11316 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_117
timestamp 1644511149
transform 1 0 11868 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_127
timestamp 1644511149
transform 1 0 12788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_143
timestamp 1644511149
transform 1 0 14260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1644511149
transform 1 0 14812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_155
timestamp 1644511149
transform 1 0 15364 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_171
timestamp 1644511149
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_183
timestamp 1644511149
transform 1 0 17940 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_199
timestamp 1644511149
transform 1 0 19412 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_205
timestamp 1644511149
transform 1 0 19964 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_211
timestamp 1644511149
transform 1 0 20516 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_217
timestamp 1644511149
transform 1 0 21068 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1644511149
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_229
timestamp 1644511149
transform 1 0 22172 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1644511149
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_241
timestamp 1644511149
transform 1 0 23276 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1644511149
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_255
timestamp 1644511149
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_261
timestamp 1644511149
transform 1 0 25116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_267
timestamp 1644511149
transform 1 0 25668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_273
timestamp 1644511149
transform 1 0 26220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_279
timestamp 1644511149
transform 1 0 26772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_285
timestamp 1644511149
transform 1 0 27324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_291
timestamp 1644511149
transform 1 0 27876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_297
timestamp 1644511149
transform 1 0 28428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_303
timestamp 1644511149
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_353
timestamp 1644511149
transform 1 0 33580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_367
timestamp 1644511149
transform 1 0 34868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_373
timestamp 1644511149
transform 1 0 35420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_379
timestamp 1644511149
transform 1 0 35972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_383
timestamp 1644511149
transform 1 0 36340 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_386
timestamp 1644511149
transform 1 0 36616 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_394
timestamp 1644511149
transform 1 0 37352 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_402
timestamp 1644511149
transform 1 0 38088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1644511149
transform 1 0 38456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_409
timestamp 1644511149
transform 1 0 38732 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_415
timestamp 1644511149
transform 1 0 39284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_423
timestamp 1644511149
transform 1 0 40020 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_439
timestamp 1644511149
transform 1 0 41492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_447
timestamp 1644511149
transform 1 0 42228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_453
timestamp 1644511149
transform 1 0 42780 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_461
timestamp 1644511149
transform 1 0 43516 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1644511149
transform 1 0 1656 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_12
timestamp 1644511149
transform 1 0 2208 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_20
timestamp 1644511149
transform 1 0 2944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_26
timestamp 1644511149
transform 1 0 3496 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_34
timestamp 1644511149
transform 1 0 4232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_40
timestamp 1644511149
transform 1 0 4784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_46
timestamp 1644511149
transform 1 0 5336 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1644511149
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_59
timestamp 1644511149
transform 1 0 6532 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_67
timestamp 1644511149
transform 1 0 7268 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_70
timestamp 1644511149
transform 1 0 7544 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_76
timestamp 1644511149
transform 1 0 8096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_82
timestamp 1644511149
transform 1 0 8648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_88
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_95
timestamp 1644511149
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_101
timestamp 1644511149
transform 1 0 10396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1644511149
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1644511149
transform 1 0 11684 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1644511149
transform 1 0 12236 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_124
timestamp 1644511149
transform 1 0 12512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_130
timestamp 1644511149
transform 1 0 13064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_136
timestamp 1644511149
transform 1 0 13616 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_142
timestamp 1644511149
transform 1 0 14168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_152
timestamp 1644511149
transform 1 0 15088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_158
timestamp 1644511149
transform 1 0 15640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1644511149
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_171
timestamp 1644511149
transform 1 0 16836 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_177
timestamp 1644511149
transform 1 0 17388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_183
timestamp 1644511149
transform 1 0 17940 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_189
timestamp 1644511149
transform 1 0 18492 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1644511149
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_201
timestamp 1644511149
transform 1 0 19596 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_207
timestamp 1644511149
transform 1 0 20148 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_213
timestamp 1644511149
transform 1 0 20700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1644511149
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_227
timestamp 1644511149
transform 1 0 21988 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_233
timestamp 1644511149
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_239
timestamp 1644511149
transform 1 0 23092 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_245
timestamp 1644511149
transform 1 0 23644 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_251
timestamp 1644511149
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_257
timestamp 1644511149
transform 1 0 24748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_263
timestamp 1644511149
transform 1 0 25300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_269
timestamp 1644511149
transform 1 0 25852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1644511149
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_283
timestamp 1644511149
transform 1 0 27140 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_289
timestamp 1644511149
transform 1 0 27692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_295
timestamp 1644511149
transform 1 0 28244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_307
timestamp 1644511149
transform 1 0 29348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_319
timestamp 1644511149
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1644511149
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_437
timestamp 1644511149
transform 1 0 41308 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_440
timestamp 1644511149
transform 1 0 41584 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_453
timestamp 1644511149
transform 1 0 42780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_469
timestamp 1644511149
transform 1 0 44252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_6
timestamp 1644511149
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_12
timestamp 1644511149
transform 1 0 2208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_18
timestamp 1644511149
transform 1 0 2760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_31
timestamp 1644511149
transform 1 0 3956 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_39
timestamp 1644511149
transform 1 0 4692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1644511149
transform 1 0 4968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_48
timestamp 1644511149
transform 1 0 5520 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_54
timestamp 1644511149
transform 1 0 6072 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_62
timestamp 1644511149
transform 1 0 6808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_68
timestamp 1644511149
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_74
timestamp 1644511149
transform 1 0 7912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1644511149
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_89
timestamp 1644511149
transform 1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_96
timestamp 1644511149
transform 1 0 9936 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_100
timestamp 1644511149
transform 1 0 10304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_104
timestamp 1644511149
transform 1 0 10672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_111
timestamp 1644511149
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_117
timestamp 1644511149
transform 1 0 11868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_123
timestamp 1644511149
transform 1 0 12420 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1644511149
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_150
timestamp 1644511149
transform 1 0 14904 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_158
timestamp 1644511149
transform 1 0 15640 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_168
timestamp 1644511149
transform 1 0 16560 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_174
timestamp 1644511149
transform 1 0 17112 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_180
timestamp 1644511149
transform 1 0 17664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1644511149
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1644511149
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_199
timestamp 1644511149
transform 1 0 19412 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_205
timestamp 1644511149
transform 1 0 19964 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_211
timestamp 1644511149
transform 1 0 20516 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_217
timestamp 1644511149
transform 1 0 21068 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1644511149
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_229
timestamp 1644511149
transform 1 0 22172 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_235
timestamp 1644511149
transform 1 0 22724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_241
timestamp 1644511149
transform 1 0 23276 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1644511149
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_255
timestamp 1644511149
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_261
timestamp 1644511149
transform 1 0 25116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_267
timestamp 1644511149
transform 1 0 25668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_273
timestamp 1644511149
transform 1 0 26220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_279
timestamp 1644511149
transform 1 0 26772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_285
timestamp 1644511149
transform 1 0 27324 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_291
timestamp 1644511149
transform 1 0 27876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1644511149
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_439
timestamp 1644511149
transform 1 0 41492 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_442
timestamp 1644511149
transform 1 0 41768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_448
timestamp 1644511149
transform 1 0 42320 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_452
timestamp 1644511149
transform 1 0 42688 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_455
timestamp 1644511149
transform 1 0 42964 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_461
timestamp 1644511149
transform 1 0 43516 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_9
timestamp 1644511149
transform 1 0 1932 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1644511149
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_25
timestamp 1644511149
transform 1 0 3404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp 1644511149
transform 1 0 3956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_37
timestamp 1644511149
transform 1 0 4508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_43
timestamp 1644511149
transform 1 0 5060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_46
timestamp 1644511149
transform 1 0 5336 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1644511149
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1644511149
transform 1 0 6808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_68
timestamp 1644511149
transform 1 0 7360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1644511149
transform 1 0 7912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1644511149
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_95
timestamp 1644511149
transform 1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_99
timestamp 1644511149
transform 1 0 10212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1644511149
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1644511149
transform 1 0 11868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_124
timestamp 1644511149
transform 1 0 12512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_131
timestamp 1644511149
transform 1 0 13156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_138
timestamp 1644511149
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_144
timestamp 1644511149
transform 1 0 14352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_150
timestamp 1644511149
transform 1 0 14904 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1644511149
transform 1 0 15456 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1644511149
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_171
timestamp 1644511149
transform 1 0 16836 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_177
timestamp 1644511149
transform 1 0 17388 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_192
timestamp 1644511149
transform 1 0 18768 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_209
timestamp 1644511149
transform 1 0 20332 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1644511149
transform 1 0 20884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_227
timestamp 1644511149
transform 1 0 21988 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_233
timestamp 1644511149
transform 1 0 22540 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_239
timestamp 1644511149
transform 1 0 23092 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_245
timestamp 1644511149
transform 1 0 23644 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_251
timestamp 1644511149
transform 1 0 24196 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_257
timestamp 1644511149
transform 1 0 24748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_263
timestamp 1644511149
transform 1 0 25300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_269
timestamp 1644511149
transform 1 0 25852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1644511149
transform 1 0 26404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_457
timestamp 1644511149
transform 1 0 43148 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_463
timestamp 1644511149
transform 1 0 43700 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_469
timestamp 1644511149
transform 1 0 44252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_6
timestamp 1644511149
transform 1 0 1656 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_14
timestamp 1644511149
transform 1 0 2392 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_17
timestamp 1644511149
transform 1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1644511149
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_31
timestamp 1644511149
transform 1 0 3956 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_37
timestamp 1644511149
transform 1 0 4508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_45
timestamp 1644511149
transform 1 0 5244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1644511149
transform 1 0 5796 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_57
timestamp 1644511149
transform 1 0 6348 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_63
timestamp 1644511149
transform 1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_70
timestamp 1644511149
transform 1 0 7544 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_76
timestamp 1644511149
transform 1 0 8096 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1644511149
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_93
timestamp 1644511149
transform 1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp 1644511149
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_107
timestamp 1644511149
transform 1 0 10948 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_120
timestamp 1644511149
transform 1 0 12144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1644511149
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1644511149
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_143
timestamp 1644511149
transform 1 0 14260 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1644511149
transform 1 0 14812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_155
timestamp 1644511149
transform 1 0 15364 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_161
timestamp 1644511149
transform 1 0 15916 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_171
timestamp 1644511149
transform 1 0 16836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1644511149
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1644511149
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_206
timestamp 1644511149
transform 1 0 20056 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_213
timestamp 1644511149
transform 1 0 20700 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_225
timestamp 1644511149
transform 1 0 21804 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_239
timestamp 1644511149
transform 1 0 23092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1644511149
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_256
timestamp 1644511149
transform 1 0 24656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_262
timestamp 1644511149
transform 1 0 25208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_268
timestamp 1644511149
transform 1 0 25760 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1644511149
transform 1 0 26864 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_292
timestamp 1644511149
transform 1 0 27968 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1644511149
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_465
timestamp 1644511149
transform 1 0 43884 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_6
timestamp 1644511149
transform 1 0 1656 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1644511149
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_18
timestamp 1644511149
transform 1 0 2760 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_24
timestamp 1644511149
transform 1 0 3312 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_34
timestamp 1644511149
transform 1 0 4232 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_40
timestamp 1644511149
transform 1 0 4784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_43
timestamp 1644511149
transform 1 0 5060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_49
timestamp 1644511149
transform 1 0 5612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1644511149
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_59
timestamp 1644511149
transform 1 0 6532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_66
timestamp 1644511149
transform 1 0 7176 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 1644511149
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_85
timestamp 1644511149
transform 1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1644511149
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1644511149
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_122
timestamp 1644511149
transform 1 0 12328 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_130
timestamp 1644511149
transform 1 0 13064 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp 1644511149
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_180
timestamp 1644511149
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_194
timestamp 1644511149
transform 1 0 18952 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_208
timestamp 1644511149
transform 1 0 20240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1644511149
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_238
timestamp 1644511149
transform 1 0 23000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_252
timestamp 1644511149
transform 1 0 24288 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_258
timestamp 1644511149
transform 1 0 24840 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1644511149
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1644511149
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_6
timestamp 1644511149
transform 1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1644511149
transform 1 0 2208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1644511149
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_31
timestamp 1644511149
transform 1 0 3956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_37
timestamp 1644511149
transform 1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_43
timestamp 1644511149
transform 1 0 5060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_49
timestamp 1644511149
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1644511149
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_63
timestamp 1644511149
transform 1 0 6900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_70
timestamp 1644511149
transform 1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1644511149
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1644511149
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_104
timestamp 1644511149
transform 1 0 10672 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1644511149
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_145
timestamp 1644511149
transform 1 0 14444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_152
timestamp 1644511149
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_159
timestamp 1644511149
transform 1 0 15732 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_166
timestamp 1644511149
transform 1 0 16376 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1644511149
transform 1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1644511149
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_207
timestamp 1644511149
transform 1 0 20148 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1644511149
transform 1 0 20700 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_217
timestamp 1644511149
transform 1 0 21068 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_224
timestamp 1644511149
transform 1 0 21712 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_230
timestamp 1644511149
transform 1 0 22264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_241
timestamp 1644511149
transform 1 0 23276 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1644511149
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_255
timestamp 1644511149
transform 1 0 24564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_261
timestamp 1644511149
transform 1 0 25116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_267
timestamp 1644511149
transform 1 0 25668 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_279
timestamp 1644511149
transform 1 0 26772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_291
timestamp 1644511149
transform 1 0 27876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp 1644511149
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_6
timestamp 1644511149
transform 1 0 1656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_13
timestamp 1644511149
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_20
timestamp 1644511149
transform 1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_26
timestamp 1644511149
transform 1 0 3496 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_34
timestamp 1644511149
transform 1 0 4232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_38
timestamp 1644511149
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_45
timestamp 1644511149
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_63
timestamp 1644511149
transform 1 0 6900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1644511149
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_94
timestamp 1644511149
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_104
timestamp 1644511149
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1644511149
transform 1 0 12420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1644511149
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1644511149
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1644511149
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_175
timestamp 1644511149
transform 1 0 17204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_192
timestamp 1644511149
transform 1 0 18768 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_204
timestamp 1644511149
transform 1 0 19872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_214
timestamp 1644511149
transform 1 0 20792 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1644511149
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_227
timestamp 1644511149
transform 1 0 21988 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_231
timestamp 1644511149
transform 1 0 22356 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_236
timestamp 1644511149
transform 1 0 22816 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_242
timestamp 1644511149
transform 1 0 23368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1644511149
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_254
timestamp 1644511149
transform 1 0 24472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_260
timestamp 1644511149
transform 1 0 25024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_266
timestamp 1644511149
transform 1 0 25576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_272
timestamp 1644511149
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1644511149
transform 1 0 1656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1644511149
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_33
timestamp 1644511149
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_37
timestamp 1644511149
transform 1 0 4508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_45
timestamp 1644511149
transform 1 0 5244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_52
timestamp 1644511149
transform 1 0 5888 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_60
timestamp 1644511149
transform 1 0 6624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_70
timestamp 1644511149
transform 1 0 7544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1644511149
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_107
timestamp 1644511149
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1644511149
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 1644511149
transform 1 0 14352 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_163
timestamp 1644511149
transform 1 0 16100 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_176
timestamp 1644511149
transform 1 0 17296 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_199
timestamp 1644511149
transform 1 0 19412 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1644511149
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1644511149
transform 1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_234
timestamp 1644511149
transform 1 0 22632 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_240
timestamp 1644511149
transform 1 0 23184 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_255
timestamp 1644511149
transform 1 0 24564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_261
timestamp 1644511149
transform 1 0 25116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_269
timestamp 1644511149
transform 1 0 25852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_283
timestamp 1644511149
transform 1 0 27140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_291
timestamp 1644511149
transform 1 0 27876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1644511149
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_10
timestamp 1644511149
transform 1 0 2024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_17
timestamp 1644511149
transform 1 0 2668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_23
timestamp 1644511149
transform 1 0 3220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_34
timestamp 1644511149
transform 1 0 4232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_40
timestamp 1644511149
transform 1 0 4784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_44
timestamp 1644511149
transform 1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1644511149
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_65
timestamp 1644511149
transform 1 0 7084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_75
timestamp 1644511149
transform 1 0 8004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_88
timestamp 1644511149
transform 1 0 9200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_102
timestamp 1644511149
transform 1 0 10488 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1644511149
transform 1 0 12420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_136
timestamp 1644511149
transform 1 0 13616 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1644511149
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_155
timestamp 1644511149
transform 1 0 15364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1644511149
transform 1 0 17112 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_178
timestamp 1644511149
transform 1 0 17480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_188
timestamp 1644511149
transform 1 0 18400 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1644511149
transform 1 0 19596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_211
timestamp 1644511149
transform 1 0 20516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1644511149
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1644511149
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_236
timestamp 1644511149
transform 1 0 22816 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_242
timestamp 1644511149
transform 1 0 23368 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_252
timestamp 1644511149
transform 1 0 24288 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_260
timestamp 1644511149
transform 1 0 25024 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_268
timestamp 1644511149
transform 1 0 25760 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_285
timestamp 1644511149
transform 1 0 27324 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_296
timestamp 1644511149
transform 1 0 28336 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_308
timestamp 1644511149
transform 1 0 29440 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_320
timestamp 1644511149
transform 1 0 30544 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1644511149
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_9
timestamp 1644511149
transform 1 0 1932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_13
timestamp 1644511149
transform 1 0 2300 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_17
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1644511149
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_34
timestamp 1644511149
transform 1 0 4232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_44
timestamp 1644511149
transform 1 0 5152 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1644511149
transform 1 0 6072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_67
timestamp 1644511149
transform 1 0 7268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1644511149
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_91
timestamp 1644511149
transform 1 0 9476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_111
timestamp 1644511149
transform 1 0 11316 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_131
timestamp 1644511149
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_147
timestamp 1644511149
transform 1 0 14628 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_157
timestamp 1644511149
transform 1 0 15548 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_171
timestamp 1644511149
transform 1 0 16836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1644511149
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1644511149
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_203
timestamp 1644511149
transform 1 0 19780 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1644511149
transform 1 0 21160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_224
timestamp 1644511149
transform 1 0 21712 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1644511149
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_236
timestamp 1644511149
transform 1 0 22816 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_242
timestamp 1644511149
transform 1 0 23368 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1644511149
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_256
timestamp 1644511149
transform 1 0 24656 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_262
timestamp 1644511149
transform 1 0 25208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_268
timestamp 1644511149
transform 1 0 25760 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_274
timestamp 1644511149
transform 1 0 26312 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_283
timestamp 1644511149
transform 1 0 27140 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_294
timestamp 1644511149
transform 1 0 28152 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_300
timestamp 1644511149
transform 1 0 28704 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1644511149
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_311
timestamp 1644511149
transform 1 0 29716 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_323
timestamp 1644511149
transform 1 0 30820 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_335
timestamp 1644511149
transform 1 0 31924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_347
timestamp 1644511149
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1644511149
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_461
timestamp 1644511149
transform 1 0 43516 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_10
timestamp 1644511149
transform 1 0 2024 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_14
timestamp 1644511149
transform 1 0 2392 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_20
timestamp 1644511149
transform 1 0 2944 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1644511149
transform 1 0 3312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_32
timestamp 1644511149
transform 1 0 4048 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_42
timestamp 1644511149
transform 1 0 4968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1644511149
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_60
timestamp 1644511149
transform 1 0 6624 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_74
timestamp 1644511149
transform 1 0 7912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1644511149
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1644511149
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_129
timestamp 1644511149
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_142
timestamp 1644511149
transform 1 0 14168 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1644511149
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1644511149
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_171
timestamp 1644511149
transform 1 0 16836 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1644511149
transform 1 0 18400 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1644511149
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_208
timestamp 1644511149
transform 1 0 20240 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_214
timestamp 1644511149
transform 1 0 20792 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_227
timestamp 1644511149
transform 1 0 21988 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_233
timestamp 1644511149
transform 1 0 22540 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_243
timestamp 1644511149
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_247
timestamp 1644511149
transform 1 0 23828 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_250
timestamp 1644511149
transform 1 0 24104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_256
timestamp 1644511149
transform 1 0 24656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_262
timestamp 1644511149
transform 1 0 25208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_268
timestamp 1644511149
transform 1 0 25760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1644511149
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_283
timestamp 1644511149
transform 1 0 27140 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_289
timestamp 1644511149
transform 1 0 27692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_295
timestamp 1644511149
transform 1 0 28244 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_307
timestamp 1644511149
transform 1 0 29348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_319
timestamp 1644511149
transform 1 0 30452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_331
timestamp 1644511149
transform 1 0 31556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_9
timestamp 1644511149
transform 1 0 1932 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_17
timestamp 1644511149
transform 1 0 2668 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1644511149
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_39
timestamp 1644511149
transform 1 0 4692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_52
timestamp 1644511149
transform 1 0 5888 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1644511149
transform 1 0 7176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_106
timestamp 1644511149
transform 1 0 10856 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_126
timestamp 1644511149
transform 1 0 12696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1644511149
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1644511149
transform 1 0 14720 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1644511149
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_168
timestamp 1644511149
transform 1 0 16560 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_183
timestamp 1644511149
transform 1 0 17940 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1644511149
transform 1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1644511149
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1644511149
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_228
timestamp 1644511149
transform 1 0 22080 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_232
timestamp 1644511149
transform 1 0 22448 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_238
timestamp 1644511149
transform 1 0 23000 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_242
timestamp 1644511149
transform 1 0 23368 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_262
timestamp 1644511149
transform 1 0 25208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_268
timestamp 1644511149
transform 1 0 25760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_274
timestamp 1644511149
transform 1 0 26312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_280
timestamp 1644511149
transform 1 0 26864 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_286
timestamp 1644511149
transform 1 0 27416 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_292
timestamp 1644511149
transform 1 0 27968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_298
timestamp 1644511149
transform 1 0 28520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1644511149
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1644511149
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_19
timestamp 1644511149
transform 1 0 2852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_29
timestamp 1644511149
transform 1 0 3772 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1644511149
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1644511149
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1644511149
transform 1 0 8280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_103
timestamp 1644511149
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_129
timestamp 1644511149
transform 1 0 12972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 1644511149
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1644511149
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_185
timestamp 1644511149
transform 1 0 18124 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_194
timestamp 1644511149
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_203
timestamp 1644511149
transform 1 0 19780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1644511149
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1644511149
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_230
timestamp 1644511149
transform 1 0 22264 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1644511149
transform 1 0 23092 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_245
timestamp 1644511149
transform 1 0 23644 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_251
timestamp 1644511149
transform 1 0 24196 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_257
timestamp 1644511149
transform 1 0 24748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_263
timestamp 1644511149
transform 1 0 25300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_269
timestamp 1644511149
transform 1 0 25852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1644511149
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_283
timestamp 1644511149
transform 1 0 27140 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_289
timestamp 1644511149
transform 1 0 27692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1644511149
transform 1 0 28244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_301
timestamp 1644511149
transform 1 0 28796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_307
timestamp 1644511149
transform 1 0 29348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_313
timestamp 1644511149
transform 1 0 29900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_325
timestamp 1644511149
transform 1 0 31004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1644511149
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_10
timestamp 1644511149
transform 1 0 2024 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1644511149
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_55
timestamp 1644511149
transform 1 0 6164 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_106
timestamp 1644511149
transform 1 0 10856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 1644511149
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1644511149
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_168
timestamp 1644511149
transform 1 0 16560 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_178
timestamp 1644511149
transform 1 0 17480 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1644511149
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1644511149
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1644511149
transform 1 0 20424 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_218
timestamp 1644511149
transform 1 0 21160 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_225
timestamp 1644511149
transform 1 0 21804 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_236
timestamp 1644511149
transform 1 0 22816 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1644511149
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_255
timestamp 1644511149
transform 1 0 24564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_261
timestamp 1644511149
transform 1 0 25116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_267
timestamp 1644511149
transform 1 0 25668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_273
timestamp 1644511149
transform 1 0 26220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_279
timestamp 1644511149
transform 1 0 26772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_285
timestamp 1644511149
transform 1 0 27324 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_291
timestamp 1644511149
transform 1 0 27876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_297
timestamp 1644511149
transform 1 0 28428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1644511149
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_311
timestamp 1644511149
transform 1 0 29716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_317
timestamp 1644511149
transform 1 0 30268 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_329
timestamp 1644511149
transform 1 0 31372 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_341
timestamp 1644511149
transform 1 0 32476 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_353
timestamp 1644511149
transform 1 0 33580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_361
timestamp 1644511149
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_9
timestamp 1644511149
transform 1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_32
timestamp 1644511149
transform 1 0 4048 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1644511149
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_74
timestamp 1644511149
transform 1 0 7912 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1644511149
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1644511149
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1644511149
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1644511149
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1644511149
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_195
timestamp 1644511149
transform 1 0 19044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_204
timestamp 1644511149
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_213
timestamp 1644511149
transform 1 0 20700 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_233
timestamp 1644511149
transform 1 0 22540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_239
timestamp 1644511149
transform 1 0 23092 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_248
timestamp 1644511149
transform 1 0 23920 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_254
timestamp 1644511149
transform 1 0 24472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_260
timestamp 1644511149
transform 1 0 25024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_266
timestamp 1644511149
transform 1 0 25576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1644511149
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_283
timestamp 1644511149
transform 1 0 27140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_289
timestamp 1644511149
transform 1 0 27692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1644511149
transform 1 0 28244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_301
timestamp 1644511149
transform 1 0 28796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_307
timestamp 1644511149
transform 1 0 29348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_313
timestamp 1644511149
transform 1 0 29900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_325
timestamp 1644511149
transform 1 0 31004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1644511149
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_9
timestamp 1644511149
transform 1 0 1932 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1644511149
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_35
timestamp 1644511149
transform 1 0 4324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_55
timestamp 1644511149
transform 1 0 6164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1644511149
transform 1 0 10856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_127
timestamp 1644511149
transform 1 0 12788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_157
timestamp 1644511149
transform 1 0 15548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1644511149
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_203
timestamp 1644511149
transform 1 0 19780 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_213
timestamp 1644511149
transform 1 0 20700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1644511149
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1644511149
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_238
timestamp 1644511149
transform 1 0 23000 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_255
timestamp 1644511149
transform 1 0 24564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_261
timestamp 1644511149
transform 1 0 25116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1644511149
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_273
timestamp 1644511149
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_279
timestamp 1644511149
transform 1 0 26772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_285
timestamp 1644511149
transform 1 0 27324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_291
timestamp 1644511149
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_297
timestamp 1644511149
transform 1 0 28428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1644511149
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_311
timestamp 1644511149
transform 1 0 29716 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_317
timestamp 1644511149
transform 1 0 30268 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_323
timestamp 1644511149
transform 1 0 30820 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_335
timestamp 1644511149
transform 1 0 31924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_347
timestamp 1644511149
transform 1 0 33028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_359
timestamp 1644511149
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_6
timestamp 1644511149
transform 1 0 1656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1644511149
transform 1 0 2760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_32
timestamp 1644511149
transform 1 0 4048 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1644511149
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_73
timestamp 1644511149
transform 1 0 7820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1644511149
transform 1 0 10120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1644511149
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_130
timestamp 1644511149
transform 1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1644511149
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1644511149
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_196
timestamp 1644511149
transform 1 0 19136 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_206
timestamp 1644511149
transform 1 0 20056 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_216
timestamp 1644511149
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1644511149
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1644511149
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_246
timestamp 1644511149
transform 1 0 23736 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_253
timestamp 1644511149
transform 1 0 24380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_259
timestamp 1644511149
transform 1 0 24932 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_265
timestamp 1644511149
transform 1 0 25484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_271
timestamp 1644511149
transform 1 0 26036 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_283
timestamp 1644511149
transform 1 0 27140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_289
timestamp 1644511149
transform 1 0 27692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_295
timestamp 1644511149
transform 1 0 28244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_301
timestamp 1644511149
transform 1 0 28796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_307
timestamp 1644511149
transform 1 0 29348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_313
timestamp 1644511149
transform 1 0 29900 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_319
timestamp 1644511149
transform 1 0 30452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_325
timestamp 1644511149
transform 1 0 31004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1644511149
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_10
timestamp 1644511149
transform 1 0 2024 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1644511149
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_40
timestamp 1644511149
transform 1 0 4784 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_60
timestamp 1644511149
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1644511149
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_106
timestamp 1644511149
transform 1 0 10856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_127
timestamp 1644511149
transform 1 0 12788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1644511149
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_158
timestamp 1644511149
transform 1 0 15640 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_178
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_205
timestamp 1644511149
transform 1 0 19964 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1644511149
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_225
timestamp 1644511149
transform 1 0 21804 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1644511149
transform 1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1644511149
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_256
timestamp 1644511149
transform 1 0 24656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_263
timestamp 1644511149
transform 1 0 25300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_269
timestamp 1644511149
transform 1 0 25852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_275
timestamp 1644511149
transform 1 0 26404 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_281
timestamp 1644511149
transform 1 0 26956 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_287
timestamp 1644511149
transform 1 0 27508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_293
timestamp 1644511149
transform 1 0 28060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1644511149
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_311
timestamp 1644511149
transform 1 0 29716 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_317
timestamp 1644511149
transform 1 0 30268 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_323
timestamp 1644511149
transform 1 0 30820 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_335
timestamp 1644511149
transform 1 0 31924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_347
timestamp 1644511149
transform 1 0 33028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_359
timestamp 1644511149
transform 1 0 34132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_18
timestamp 1644511149
transform 1 0 2760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_32
timestamp 1644511149
transform 1 0 4048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_60
timestamp 1644511149
transform 1 0 6624 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_106
timestamp 1644511149
transform 1 0 10856 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_130
timestamp 1644511149
transform 1 0 13064 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_155
timestamp 1644511149
transform 1 0 15364 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_185
timestamp 1644511149
transform 1 0 18124 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_199
timestamp 1644511149
transform 1 0 19412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1644511149
transform 1 0 20424 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_231
timestamp 1644511149
transform 1 0 22356 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_243
timestamp 1644511149
transform 1 0 23460 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_253
timestamp 1644511149
transform 1 0 24380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_263
timestamp 1644511149
transform 1 0 25300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_270
timestamp 1644511149
transform 1 0 25944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_283
timestamp 1644511149
transform 1 0 27140 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_289
timestamp 1644511149
transform 1 0 27692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_295
timestamp 1644511149
transform 1 0 28244 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_301
timestamp 1644511149
transform 1 0 28796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_307
timestamp 1644511149
transform 1 0 29348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_313
timestamp 1644511149
transform 1 0 29900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_319
timestamp 1644511149
transform 1 0 30452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_331
timestamp 1644511149
transform 1 0 31556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_10
timestamp 1644511149
transform 1 0 2024 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1644511149
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_39
timestamp 1644511149
transform 1 0 4692 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_59
timestamp 1644511149
transform 1 0 6532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_158
timestamp 1644511149
transform 1 0 15640 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1644511149
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_203
timestamp 1644511149
transform 1 0 19780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_213
timestamp 1644511149
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_223
timestamp 1644511149
transform 1 0 21620 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_241
timestamp 1644511149
transform 1 0 23276 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_256
timestamp 1644511149
transform 1 0 24656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_263
timestamp 1644511149
transform 1 0 25300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_269
timestamp 1644511149
transform 1 0 25852 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_275
timestamp 1644511149
transform 1 0 26404 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_281
timestamp 1644511149
transform 1 0 26956 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_287
timestamp 1644511149
transform 1 0 27508 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_293
timestamp 1644511149
transform 1 0 28060 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1644511149
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_311
timestamp 1644511149
transform 1 0 29716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_317
timestamp 1644511149
transform 1 0 30268 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_329
timestamp 1644511149
transform 1 0 31372 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_341
timestamp 1644511149
transform 1 0 32476 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_353
timestamp 1644511149
transform 1 0 33580 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_361
timestamp 1644511149
transform 1 0 34316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_12
timestamp 1644511149
transform 1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1644511149
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1644511149
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1644511149
transform 1 0 6808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1644511149
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_130
timestamp 1644511149
transform 1 0 13064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_151
timestamp 1644511149
transform 1 0 14996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1644511149
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_198
timestamp 1644511149
transform 1 0 19320 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1644511149
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1644511149
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_231
timestamp 1644511149
transform 1 0 22356 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_241
timestamp 1644511149
transform 1 0 23276 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_248
timestamp 1644511149
transform 1 0 23920 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_255
timestamp 1644511149
transform 1 0 24564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_267
timestamp 1644511149
transform 1 0 25668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_283
timestamp 1644511149
transform 1 0 27140 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_289
timestamp 1644511149
transform 1 0 27692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_295
timestamp 1644511149
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_301
timestamp 1644511149
transform 1 0 28796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_307
timestamp 1644511149
transform 1 0 29348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_313
timestamp 1644511149
transform 1 0 29900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_319
timestamp 1644511149
transform 1 0 30452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1644511149
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_10
timestamp 1644511149
transform 1 0 2024 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_39
timestamp 1644511149
transform 1 0 4692 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_59
timestamp 1644511149
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1644511149
transform 1 0 9108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1644511149
transform 1 0 11408 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1644511149
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_143
timestamp 1644511149
transform 1 0 14260 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1644511149
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_178
timestamp 1644511149
transform 1 0 17480 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_203
timestamp 1644511149
transform 1 0 19780 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_213
timestamp 1644511149
transform 1 0 20700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_223
timestamp 1644511149
transform 1 0 21620 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_239
timestamp 1644511149
transform 1 0 23092 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_244
timestamp 1644511149
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_255
timestamp 1644511149
transform 1 0 24564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1644511149
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_283
timestamp 1644511149
transform 1 0 27140 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_295
timestamp 1644511149
transform 1 0 28244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_311
timestamp 1644511149
transform 1 0 29716 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_323
timestamp 1644511149
transform 1 0 30820 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_335
timestamp 1644511149
transform 1 0 31924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_347
timestamp 1644511149
transform 1 0 33028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1644511149
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_12
timestamp 1644511149
transform 1 0 2208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_32
timestamp 1644511149
transform 1 0 4048 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_61
timestamp 1644511149
transform 1 0 6716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp 1644511149
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_134
timestamp 1644511149
transform 1 0 13432 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_140
timestamp 1644511149
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_158
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1644511149
transform 1 0 17572 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_189
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_199
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_213
timestamp 1644511149
transform 1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_231
timestamp 1644511149
transform 1 0 22356 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_245
timestamp 1644511149
transform 1 0 23644 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_251
timestamp 1644511149
transform 1 0 24196 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_255
timestamp 1644511149
transform 1 0 24564 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_262
timestamp 1644511149
transform 1 0 25208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_268
timestamp 1644511149
transform 1 0 25760 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1644511149
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_283
timestamp 1644511149
transform 1 0 27140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_289
timestamp 1644511149
transform 1 0 27692 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_295
timestamp 1644511149
transform 1 0 28244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_301
timestamp 1644511149
transform 1 0 28796 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_313
timestamp 1644511149
transform 1 0 29900 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_325
timestamp 1644511149
transform 1 0 31004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1644511149
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_9
timestamp 1644511149
transform 1 0 1932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_13
timestamp 1644511149
transform 1 0 2300 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_35
timestamp 1644511149
transform 1 0 4324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_55
timestamp 1644511149
transform 1 0 6164 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_106
timestamp 1644511149
transform 1 0 10856 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1644511149
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1644511149
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1644511149
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_183
timestamp 1644511149
transform 1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_211
timestamp 1644511149
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1644511149
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_227
timestamp 1644511149
transform 1 0 21988 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1644511149
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_247
timestamp 1644511149
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_255
timestamp 1644511149
transform 1 0 24564 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_261
timestamp 1644511149
transform 1 0 25116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_267
timestamp 1644511149
transform 1 0 25668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_273
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_279
timestamp 1644511149
transform 1 0 26772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_285
timestamp 1644511149
transform 1 0 27324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_291
timestamp 1644511149
transform 1 0 27876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_297
timestamp 1644511149
transform 1 0 28428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_313
timestamp 1644511149
transform 1 0 29900 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_325
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_337
timestamp 1644511149
transform 1 0 32108 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_349
timestamp 1644511149
transform 1 0 33212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1644511149
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_5
timestamp 1644511149
transform 1 0 1564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_18
timestamp 1644511149
transform 1 0 2760 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_32
timestamp 1644511149
transform 1 0 4048 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1644511149
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1644511149
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_134
timestamp 1644511149
transform 1 0 13432 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_140
timestamp 1644511149
transform 1 0 13984 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_157
timestamp 1644511149
transform 1 0 15548 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1644511149
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1644511149
transform 1 0 17480 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_191
timestamp 1644511149
transform 1 0 18676 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_201
timestamp 1644511149
transform 1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_211
timestamp 1644511149
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1644511149
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_233
timestamp 1644511149
transform 1 0 22540 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_240
timestamp 1644511149
transform 1 0 23184 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_246
timestamp 1644511149
transform 1 0 23736 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1644511149
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_258
timestamp 1644511149
transform 1 0 24840 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_264
timestamp 1644511149
transform 1 0 25392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_270
timestamp 1644511149
transform 1 0 25944 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_283
timestamp 1644511149
transform 1 0 27140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_289
timestamp 1644511149
transform 1 0 27692 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_297
timestamp 1644511149
transform 1 0 28428 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_303
timestamp 1644511149
transform 1 0 28980 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_308
timestamp 1644511149
transform 1 0 29440 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_312
timestamp 1644511149
transform 1 0 29808 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_11
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1644511149
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_33
timestamp 1644511149
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_55
timestamp 1644511149
transform 1 0 6164 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1644511149
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_89
timestamp 1644511149
transform 1 0 9292 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_111
timestamp 1644511149
transform 1 0 11316 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_131
timestamp 1644511149
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp 1644511149
transform 1 0 14996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_178
timestamp 1644511149
transform 1 0 17480 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_188
timestamp 1644511149
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_203
timestamp 1644511149
transform 1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_211
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_225
timestamp 1644511149
transform 1 0 21804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_232
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_239
timestamp 1644511149
transform 1 0 23092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_255
timestamp 1644511149
transform 1 0 24564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_267
timestamp 1644511149
transform 1 0 25668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_275
timestamp 1644511149
transform 1 0 26404 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_278
timestamp 1644511149
transform 1 0 26680 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_286
timestamp 1644511149
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1644511149
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1644511149
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_359
timestamp 1644511149
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_6
timestamp 1644511149
transform 1 0 1656 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_19
timestamp 1644511149
transform 1 0 2852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_32
timestamp 1644511149
transform 1 0 4048 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_61
timestamp 1644511149
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_83
timestamp 1644511149
transform 1 0 8740 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_129
timestamp 1644511149
transform 1 0 12972 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_143
timestamp 1644511149
transform 1 0 14260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1644511149
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_186
timestamp 1644511149
transform 1 0 18216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_203
timestamp 1644511149
transform 1 0 19780 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_211
timestamp 1644511149
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1644511149
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_235
timestamp 1644511149
transform 1 0 22724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_241
timestamp 1644511149
transform 1 0 23276 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_247
timestamp 1644511149
transform 1 0 23828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_253
timestamp 1644511149
transform 1 0 24380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_258
timestamp 1644511149
transform 1 0 24840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_266
timestamp 1644511149
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1644511149
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_289
timestamp 1644511149
transform 1 0 27692 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_295
timestamp 1644511149
transform 1 0 28244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_303
timestamp 1644511149
transform 1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_311
timestamp 1644511149
transform 1 0 29716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_342
timestamp 1644511149
transform 1 0 32568 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_350
timestamp 1644511149
transform 1 0 33304 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_358
timestamp 1644511149
transform 1 0 34040 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_363
timestamp 1644511149
transform 1 0 34500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_369
timestamp 1644511149
transform 1 0 35052 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_377
timestamp 1644511149
transform 1 0 35788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1644511149
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1644511149
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_55
timestamp 1644511149
transform 1 0 6164 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1644511149
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1644511149
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_120
timestamp 1644511149
transform 1 0 12144 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_151
timestamp 1644511149
transform 1 0 14996 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_169
timestamp 1644511149
transform 1 0 16652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_176
timestamp 1644511149
transform 1 0 17296 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_186
timestamp 1644511149
transform 1 0 18216 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_205
timestamp 1644511149
transform 1 0 19964 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_211
timestamp 1644511149
transform 1 0 20516 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_222
timestamp 1644511149
transform 1 0 21528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1644511149
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_244
timestamp 1644511149
transform 1 0 23552 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_261
timestamp 1644511149
transform 1 0 25116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_269
timestamp 1644511149
transform 1 0 25852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_275
timestamp 1644511149
transform 1 0 26404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_283
timestamp 1644511149
transform 1 0 27140 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_291
timestamp 1644511149
transform 1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_317
timestamp 1644511149
transform 1 0 30268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_325
timestamp 1644511149
transform 1 0 31004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_331
timestamp 1644511149
transform 1 0 31556 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_335
timestamp 1644511149
transform 1 0 31924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_338
timestamp 1644511149
transform 1 0 32200 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_346
timestamp 1644511149
transform 1 0 32936 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_358
timestamp 1644511149
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_373
timestamp 1644511149
transform 1 0 35420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_381
timestamp 1644511149
transform 1 0 36156 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_393
timestamp 1644511149
transform 1 0 37260 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_405
timestamp 1644511149
transform 1 0 38364 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_417
timestamp 1644511149
transform 1 0 39468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_6
timestamp 1644511149
transform 1 0 1656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_14
timestamp 1644511149
transform 1 0 2392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_24
timestamp 1644511149
transform 1 0 3312 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_38
timestamp 1644511149
transform 1 0 4600 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1644511149
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_62
timestamp 1644511149
transform 1 0 6808 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_87
timestamp 1644511149
transform 1 0 9108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_101
timestamp 1644511149
transform 1 0 10396 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1644511149
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1644511149
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_127
timestamp 1644511149
transform 1 0 12788 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_138
timestamp 1644511149
transform 1 0 13800 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_154
timestamp 1644511149
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1644511149
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1644511149
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_190
timestamp 1644511149
transform 1 0 18584 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_200
timestamp 1644511149
transform 1 0 19504 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_206
timestamp 1644511149
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_212
timestamp 1644511149
transform 1 0 20608 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1644511149
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_227
timestamp 1644511149
transform 1 0 21988 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_243
timestamp 1644511149
transform 1 0 23460 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_253
timestamp 1644511149
transform 1 0 24380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_265
timestamp 1644511149
transform 1 0 25484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_270
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1644511149
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_289
timestamp 1644511149
transform 1 0 27692 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_297
timestamp 1644511149
transform 1 0 28428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_301
timestamp 1644511149
transform 1 0 28796 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_306
timestamp 1644511149
transform 1 0 29256 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_310
timestamp 1644511149
transform 1 0 29624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_313
timestamp 1644511149
transform 1 0 29900 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_325
timestamp 1644511149
transform 1 0 31004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1644511149
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_354
timestamp 1644511149
transform 1 0 33672 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_366
timestamp 1644511149
transform 1 0 34776 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_378
timestamp 1644511149
transform 1 0 35880 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1644511149
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_7
timestamp 1644511149
transform 1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_14
timestamp 1644511149
transform 1 0 2392 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1644511149
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_33
timestamp 1644511149
transform 1 0 4140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_46
timestamp 1644511149
transform 1 0 5336 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_60
timestamp 1644511149
transform 1 0 6624 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_106
timestamp 1644511149
transform 1 0 10856 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_120
timestamp 1644511149
transform 1 0 12144 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_151
timestamp 1644511149
transform 1 0 14996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_161
timestamp 1644511149
transform 1 0 15916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_171
timestamp 1644511149
transform 1 0 16836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1644511149
transform 1 0 17756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_199
timestamp 1644511149
transform 1 0 19412 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_205
timestamp 1644511149
transform 1 0 19964 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_211
timestamp 1644511149
transform 1 0 20516 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_217
timestamp 1644511149
transform 1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1644511149
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_229
timestamp 1644511149
transform 1 0 22172 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1644511149
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_241
timestamp 1644511149
transform 1 0 23276 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1644511149
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_255
timestamp 1644511149
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1644511149
transform 1 0 25300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_275
timestamp 1644511149
transform 1 0 26404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_279
timestamp 1644511149
transform 1 0 26772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_295
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_311
timestamp 1644511149
transform 1 0 29716 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_323
timestamp 1644511149
transform 1 0 30820 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_335
timestamp 1644511149
transform 1 0 31924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_347
timestamp 1644511149
transform 1 0 33028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1644511149
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 1644511149
transform 1 0 2392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1644511149
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_29
timestamp 1644511149
transform 1 0 3772 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1644511149
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1644511149
transform 1 0 6808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_87
timestamp 1644511149
transform 1 0 9108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_101
timestamp 1644511149
transform 1 0 10396 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_122
timestamp 1644511149
transform 1 0 12328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_132
timestamp 1644511149
transform 1 0 13248 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_140
timestamp 1644511149
transform 1 0 13984 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_146
timestamp 1644511149
transform 1 0 14536 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1644511149
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_179
timestamp 1644511149
transform 1 0 17572 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_185
timestamp 1644511149
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_191
timestamp 1644511149
transform 1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_197
timestamp 1644511149
transform 1 0 19228 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1644511149
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_227
timestamp 1644511149
transform 1 0 21988 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_233
timestamp 1644511149
transform 1 0 22540 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_239
timestamp 1644511149
transform 1 0 23092 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_245
timestamp 1644511149
transform 1 0 23644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_251
timestamp 1644511149
transform 1 0 24196 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_263
timestamp 1644511149
transform 1 0 25300 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1644511149
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_291
timestamp 1644511149
transform 1 0 27876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_303
timestamp 1644511149
transform 1 0 28980 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_315
timestamp 1644511149
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1644511149
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_6
timestamp 1644511149
transform 1 0 1656 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1644511149
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1644511149
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_31
timestamp 1644511149
transform 1 0 3956 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_51
timestamp 1644511149
transform 1 0 5796 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_64
timestamp 1644511149
transform 1 0 6992 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1644511149
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_95
timestamp 1644511149
transform 1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_108
timestamp 1644511149
transform 1 0 11040 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1644511149
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1644511149
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_145
timestamp 1644511149
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_159
timestamp 1644511149
transform 1 0 15732 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_175
timestamp 1644511149
transform 1 0 17204 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_181
timestamp 1644511149
transform 1 0 17756 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_185
timestamp 1644511149
transform 1 0 18124 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_190
timestamp 1644511149
transform 1 0 18584 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_201
timestamp 1644511149
transform 1 0 19596 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_215
timestamp 1644511149
transform 1 0 20884 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_229
timestamp 1644511149
transform 1 0 22172 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_241
timestamp 1644511149
transform 1 0 23276 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1644511149
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_6
timestamp 1644511149
transform 1 0 1656 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_12
timestamp 1644511149
transform 1 0 2208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_16
timestamp 1644511149
transform 1 0 2576 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_20
timestamp 1644511149
transform 1 0 2944 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_28
timestamp 1644511149
transform 1 0 3680 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_35
timestamp 1644511149
transform 1 0 4324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_42
timestamp 1644511149
transform 1 0 4968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1644511149
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1644511149
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_71
timestamp 1644511149
transform 1 0 7636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_85
timestamp 1644511149
transform 1 0 8924 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_99
timestamp 1644511149
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1644511149
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1644511149
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_127
timestamp 1644511149
transform 1 0 12788 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_135
timestamp 1644511149
transform 1 0 13524 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_143
timestamp 1644511149
transform 1 0 14260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_150
timestamp 1644511149
transform 1 0 14904 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1644511149
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_162
timestamp 1644511149
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_171
timestamp 1644511149
transform 1 0 16836 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_175
timestamp 1644511149
transform 1 0 17204 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_186
timestamp 1644511149
transform 1 0 18216 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_200
timestamp 1644511149
transform 1 0 19504 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_214
timestamp 1644511149
transform 1 0 20792 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_233
timestamp 1644511149
transform 1 0 22540 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1644511149
transform 1 0 23644 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1644511149
transform 1 0 24748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1644511149
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1644511149
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_313
timestamp 1644511149
transform 1 0 29900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_321
timestamp 1644511149
transform 1 0 30636 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_6
timestamp 1644511149
transform 1 0 1656 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_12
timestamp 1644511149
transform 1 0 2208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_18
timestamp 1644511149
transform 1 0 2760 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1644511149
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_31
timestamp 1644511149
transform 1 0 3956 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_35
timestamp 1644511149
transform 1 0 4324 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_38
timestamp 1644511149
transform 1 0 4600 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_45
timestamp 1644511149
transform 1 0 5244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_52
timestamp 1644511149
transform 1 0 5888 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1644511149
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_75
timestamp 1644511149
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1644511149
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_101
timestamp 1644511149
transform 1 0 10396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_111
timestamp 1644511149
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_119
timestamp 1644511149
transform 1 0 12052 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_127
timestamp 1644511149
transform 1 0 12788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_134
timestamp 1644511149
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_144
timestamp 1644511149
transform 1 0 14352 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_150
timestamp 1644511149
transform 1 0 14904 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_158
timestamp 1644511149
transform 1 0 15640 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_166
timestamp 1644511149
transform 1 0 16376 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_172
timestamp 1644511149
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_176
timestamp 1644511149
transform 1 0 17296 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_180
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_186
timestamp 1644511149
transform 1 0 18216 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_207
timestamp 1644511149
transform 1 0 20148 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_215
timestamp 1644511149
transform 1 0 20884 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_223
timestamp 1644511149
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_231
timestamp 1644511149
transform 1 0 22356 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_243
timestamp 1644511149
transform 1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_293
timestamp 1644511149
transform 1 0 28060 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_317
timestamp 1644511149
transform 1 0 30268 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_325
timestamp 1644511149
transform 1 0 31004 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_341
timestamp 1644511149
transform 1 0 32476 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_353
timestamp 1644511149
transform 1 0 33580 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1644511149
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_6
timestamp 1644511149
transform 1 0 1656 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1644511149
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_20
timestamp 1644511149
transform 1 0 2944 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_26
timestamp 1644511149
transform 1 0 3496 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_32
timestamp 1644511149
transform 1 0 4048 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_41
timestamp 1644511149
transform 1 0 4876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1644511149
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_63
timestamp 1644511149
transform 1 0 6900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_73
timestamp 1644511149
transform 1 0 7820 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_83
timestamp 1644511149
transform 1 0 8740 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_89
timestamp 1644511149
transform 1 0 9292 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_96
timestamp 1644511149
transform 1 0 9936 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_106
timestamp 1644511149
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_117
timestamp 1644511149
transform 1 0 11868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_124
timestamp 1644511149
transform 1 0 12512 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_131
timestamp 1644511149
transform 1 0 13156 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_138
timestamp 1644511149
transform 1 0 13800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_144
timestamp 1644511149
transform 1 0 14352 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_152
timestamp 1644511149
transform 1 0 15088 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_155
timestamp 1644511149
transform 1 0 15364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_175
timestamp 1644511149
transform 1 0 17204 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_187
timestamp 1644511149
transform 1 0 18308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_199
timestamp 1644511149
transform 1 0 19412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_233
timestamp 1644511149
transform 1 0 22540 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1644511149
transform 1 0 24748 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1644511149
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1644511149
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_345
timestamp 1644511149
transform 1 0 32844 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_357
timestamp 1644511149
transform 1 0 33948 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_369
timestamp 1644511149
transform 1 0 35052 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_381
timestamp 1644511149
transform 1 0 36156 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1644511149
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_9
timestamp 1644511149
transform 1 0 1932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1644511149
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_31
timestamp 1644511149
transform 1 0 3956 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_37
timestamp 1644511149
transform 1 0 4508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_43
timestamp 1644511149
transform 1 0 5060 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_49
timestamp 1644511149
transform 1 0 5612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_57
timestamp 1644511149
transform 1 0 6348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_60
timestamp 1644511149
transform 1 0 6624 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_67
timestamp 1644511149
transform 1 0 7268 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_92
timestamp 1644511149
transform 1 0 9568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_100
timestamp 1644511149
transform 1 0 10304 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_107
timestamp 1644511149
transform 1 0 10948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1644511149
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_120
timestamp 1644511149
transform 1 0 12144 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_126
timestamp 1644511149
transform 1 0 12696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1644511149
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_143
timestamp 1644511149
transform 1 0 14260 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1644511149
transform 1 0 14812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_155
timestamp 1644511149
transform 1 0 15364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_161
timestamp 1644511149
transform 1 0 15916 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_167
timestamp 1644511149
transform 1 0 16468 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_173
timestamp 1644511149
transform 1 0 17020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_179
timestamp 1644511149
transform 1 0 17572 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_185
timestamp 1644511149
transform 1 0 18124 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1644511149
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_199
timestamp 1644511149
transform 1 0 19412 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_211
timestamp 1644511149
transform 1 0 20516 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_223
timestamp 1644511149
transform 1 0 21620 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_229
timestamp 1644511149
transform 1 0 22172 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_241
timestamp 1644511149
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1644511149
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_9
timestamp 1644511149
transform 1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_13
timestamp 1644511149
transform 1 0 2300 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_16
timestamp 1644511149
transform 1 0 2576 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_22
timestamp 1644511149
transform 1 0 3128 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_28
timestamp 1644511149
transform 1 0 3680 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_34
timestamp 1644511149
transform 1 0 4232 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_40
timestamp 1644511149
transform 1 0 4784 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_46
timestamp 1644511149
transform 1 0 5336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1644511149
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_61
timestamp 1644511149
transform 1 0 6716 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_68
timestamp 1644511149
transform 1 0 7360 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_75
timestamp 1644511149
transform 1 0 8004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_82
timestamp 1644511149
transform 1 0 8648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_90
timestamp 1644511149
transform 1 0 9384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_97
timestamp 1644511149
transform 1 0 10028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_104
timestamp 1644511149
transform 1 0 10672 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_115
timestamp 1644511149
transform 1 0 11684 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_121
timestamp 1644511149
transform 1 0 12236 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_127
timestamp 1644511149
transform 1 0 12788 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_133
timestamp 1644511149
transform 1 0 13340 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_139
timestamp 1644511149
transform 1 0 13892 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_145
timestamp 1644511149
transform 1 0 14444 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_151
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_157
timestamp 1644511149
transform 1 0 15548 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1644511149
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_171
timestamp 1644511149
transform 1 0 16836 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_177
timestamp 1644511149
transform 1 0 17388 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_189
timestamp 1644511149
transform 1 0 18492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_201
timestamp 1644511149
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_213
timestamp 1644511149
transform 1 0 20700 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1644511149
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_6
timestamp 1644511149
transform 1 0 1656 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_16
timestamp 1644511149
transform 1 0 2576 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_22
timestamp 1644511149
transform 1 0 3128 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_31
timestamp 1644511149
transform 1 0 3956 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_37
timestamp 1644511149
transform 1 0 4508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_43
timestamp 1644511149
transform 1 0 5060 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_47
timestamp 1644511149
transform 1 0 5428 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_50
timestamp 1644511149
transform 1 0 5704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_56
timestamp 1644511149
transform 1 0 6256 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_62
timestamp 1644511149
transform 1 0 6808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_68
timestamp 1644511149
transform 1 0 7360 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1644511149
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_88
timestamp 1644511149
transform 1 0 9200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_95
timestamp 1644511149
transform 1 0 9844 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_101
timestamp 1644511149
transform 1 0 10396 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_107
timestamp 1644511149
transform 1 0 10948 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_110
timestamp 1644511149
transform 1 0 11224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_116
timestamp 1644511149
transform 1 0 11776 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_122
timestamp 1644511149
transform 1 0 12328 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_128
timestamp 1644511149
transform 1 0 12880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1644511149
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_143
timestamp 1644511149
transform 1 0 14260 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_149
timestamp 1644511149
transform 1 0 14812 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_161
timestamp 1644511149
transform 1 0 15916 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_173
timestamp 1644511149
transform 1 0 17020 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_185
timestamp 1644511149
transform 1 0 18124 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1644511149
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_5
timestamp 1644511149
transform 1 0 1564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_11
timestamp 1644511149
transform 1 0 2116 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_21
timestamp 1644511149
transform 1 0 3036 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_33
timestamp 1644511149
transform 1 0 4140 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_45
timestamp 1644511149
transform 1 0 5244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_49
timestamp 1644511149
transform 1 0 5612 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1644511149
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_61
timestamp 1644511149
transform 1 0 6716 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_64
timestamp 1644511149
transform 1 0 6992 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_70
timestamp 1644511149
transform 1 0 7544 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_73
timestamp 1644511149
transform 1 0 7820 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_79
timestamp 1644511149
transform 1 0 8372 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_85
timestamp 1644511149
transform 1 0 8924 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_91
timestamp 1644511149
transform 1 0 9476 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1644511149
transform 1 0 10028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_103
timestamp 1644511149
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_115
timestamp 1644511149
transform 1 0 11684 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_121
timestamp 1644511149
transform 1 0 12236 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_127
timestamp 1644511149
transform 1 0 12788 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_130
timestamp 1644511149
transform 1 0 13064 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_136
timestamp 1644511149
transform 1 0 13616 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_142
timestamp 1644511149
transform 1 0 14168 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_154
timestamp 1644511149
transform 1 0 15272 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1644511149
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_6
timestamp 1644511149
transform 1 0 1656 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_12
timestamp 1644511149
transform 1 0 2208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_18
timestamp 1644511149
transform 1 0 2760 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1644511149
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_31
timestamp 1644511149
transform 1 0 3956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_43
timestamp 1644511149
transform 1 0 5060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_55
timestamp 1644511149
transform 1 0 6164 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_63
timestamp 1644511149
transform 1 0 6900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_66
timestamp 1644511149
transform 1 0 7176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_72
timestamp 1644511149
transform 1 0 7728 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1644511149
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_87
timestamp 1644511149
transform 1 0 9108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_93
timestamp 1644511149
transform 1 0 9660 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_99
timestamp 1644511149
transform 1 0 10212 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_102
timestamp 1644511149
transform 1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_108
timestamp 1644511149
transform 1 0 11040 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_114
timestamp 1644511149
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_120
timestamp 1644511149
transform 1 0 12144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_126
timestamp 1644511149
transform 1 0 12696 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_132
timestamp 1644511149
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_5
timestamp 1644511149
transform 1 0 1564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1644511149
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_17
timestamp 1644511149
transform 1 0 2668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_29
timestamp 1644511149
transform 1 0 3772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_41
timestamp 1644511149
transform 1 0 4876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1644511149
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_77
timestamp 1644511149
transform 1 0 8188 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_83
timestamp 1644511149
transform 1 0 8740 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_87
timestamp 1644511149
transform 1 0 9108 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_90
timestamp 1644511149
transform 1 0 9384 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_96
timestamp 1644511149
transform 1 0 9936 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_102
timestamp 1644511149
transform 1 0 10488 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_115
timestamp 1644511149
transform 1 0 11684 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_121
timestamp 1644511149
transform 1 0 12236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_127
timestamp 1644511149
transform 1 0 12788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_139
timestamp 1644511149
transform 1 0 13892 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_151
timestamp 1644511149
transform 1 0 14996 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1644511149
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_6
timestamp 1644511149
transform 1 0 1656 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 1644511149
transform 1 0 3220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_87
timestamp 1644511149
transform 1 0 9108 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1644511149
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_94
timestamp 1644511149
transform 1 0 9752 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_106
timestamp 1644511149
transform 1 0 10856 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_110
timestamp 1644511149
transform 1 0 11224 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_122
timestamp 1644511149
transform 1 0 12328 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 1644511149
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_9
timestamp 1644511149
transform 1 0 1932 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_21
timestamp 1644511149
transform 1 0 3036 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_33
timestamp 1644511149
transform 1 0 4140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_45
timestamp 1644511149
transform 1 0 5244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1644511149
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_85
timestamp 1644511149
transform 1 0 8924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_97
timestamp 1644511149
transform 1 0 10028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1644511149
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_6
timestamp 1644511149
transform 1 0 1656 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_12
timestamp 1644511149
transform 1 0 2208 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_6
timestamp 1644511149
transform 1 0 1656 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_12
timestamp 1644511149
transform 1 0 2208 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_24
timestamp 1644511149
transform 1 0 3312 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_36
timestamp 1644511149
transform 1 0 4416 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_48
timestamp 1644511149
transform 1 0 5520 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_457
timestamp 1644511149
transform 1 0 43148 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_469
timestamp 1644511149
transform 1 0 44252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_6
timestamp 1644511149
transform 1 0 1656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_12
timestamp 1644511149
transform 1 0 2208 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_24
timestamp 1644511149
transform 1 0 3312 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_36
timestamp 1644511149
transform 1 0 4416 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_48
timestamp 1644511149
transform 1 0 5520 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_9
timestamp 1644511149
transform 1 0 1932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1644511149
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_6
timestamp 1644511149
transform 1 0 1656 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_12
timestamp 1644511149
transform 1 0 2208 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_24
timestamp 1644511149
transform 1 0 3312 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_36
timestamp 1644511149
transform 1 0 4416 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_48
timestamp 1644511149
transform 1 0 5520 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_6
timestamp 1644511149
transform 1 0 1656 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_12
timestamp 1644511149
transform 1 0 2208 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_24
timestamp 1644511149
transform 1 0 3312 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_36
timestamp 1644511149
transform 1 0 4416 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_48
timestamp 1644511149
transform 1 0 5520 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_5
timestamp 1644511149
transform 1 0 1564 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_11
timestamp 1644511149
transform 1 0 2116 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_17
timestamp 1644511149
transform 1 0 2668 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_25
timestamp 1644511149
transform 1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_465
timestamp 1644511149
transform 1 0 43884 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_6
timestamp 1644511149
transform 1 0 1656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_12
timestamp 1644511149
transform 1 0 2208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_18
timestamp 1644511149
transform 1 0 2760 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_24
timestamp 1644511149
transform 1 0 3312 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_36
timestamp 1644511149
transform 1 0 4416 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_48
timestamp 1644511149
transform 1 0 5520 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_465
timestamp 1644511149
transform 1 0 43884 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_6
timestamp 1644511149
transform 1 0 1656 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_13
timestamp 1644511149
transform 1 0 2300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 1644511149
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_31
timestamp 1644511149
transform 1 0 3956 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_37
timestamp 1644511149
transform 1 0 4508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_43
timestamp 1644511149
transform 1 0 5060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_55
timestamp 1644511149
transform 1 0 6164 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_67
timestamp 1644511149
transform 1 0 7268 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_79
timestamp 1644511149
transform 1 0 8372 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_229
timestamp 1644511149
transform 1 0 22172 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_237
timestamp 1644511149
transform 1 0 22908 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_242
timestamp 1644511149
transform 1 0 23368 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1644511149
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_255
timestamp 1644511149
transform 1 0 24564 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_259
timestamp 1644511149
transform 1 0 24932 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_262
timestamp 1644511149
transform 1 0 25208 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_276
timestamp 1644511149
transform 1 0 26496 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_288
timestamp 1644511149
transform 1 0 27600 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_300
timestamp 1644511149
transform 1 0 28704 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_319
timestamp 1644511149
transform 1 0 30452 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_325
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_328
timestamp 1644511149
transform 1 0 31280 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_340
timestamp 1644511149
transform 1 0 32384 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_352
timestamp 1644511149
transform 1 0 33488 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_355
timestamp 1644511149
transform 1 0 33764 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_397
timestamp 1644511149
transform 1 0 37628 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_409
timestamp 1644511149
transform 1 0 38732 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_417
timestamp 1644511149
transform 1 0 39468 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_423
timestamp 1644511149
transform 1 0 40020 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_453
timestamp 1644511149
transform 1 0 42780 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_465
timestamp 1644511149
transform 1 0 43884 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_9
timestamp 1644511149
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_16
timestamp 1644511149
transform 1 0 2576 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_22
timestamp 1644511149
transform 1 0 3128 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_28
timestamp 1644511149
transform 1 0 3680 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_34
timestamp 1644511149
transform 1 0 4232 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_40
timestamp 1644511149
transform 1 0 4784 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_43
timestamp 1644511149
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_59
timestamp 1644511149
transform 1 0 6532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_71
timestamp 1644511149
transform 1 0 7636 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_77
timestamp 1644511149
transform 1 0 8188 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_80
timestamp 1644511149
transform 1 0 8464 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_88
timestamp 1644511149
transform 1 0 9200 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_99
timestamp 1644511149
transform 1 0 10212 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_108
timestamp 1644511149
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_119
timestamp 1644511149
transform 1 0 12052 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_127
timestamp 1644511149
transform 1 0 12788 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_133
timestamp 1644511149
transform 1 0 13340 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_141
timestamp 1644511149
transform 1 0 14076 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_146
timestamp 1644511149
transform 1 0 14536 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_158
timestamp 1644511149
transform 1 0 15640 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1644511149
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_175
timestamp 1644511149
transform 1 0 17204 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_187
timestamp 1644511149
transform 1 0 18308 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_197
timestamp 1644511149
transform 1 0 19228 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_203
timestamp 1644511149
transform 1 0 19780 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_215
timestamp 1644511149
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_229
timestamp 1644511149
transform 1 0 22172 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_235
timestamp 1644511149
transform 1 0 22724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_241
timestamp 1644511149
transform 1 0 23276 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_247
timestamp 1644511149
transform 1 0 23828 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_257
timestamp 1644511149
transform 1 0 24748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_263
timestamp 1644511149
transform 1 0 25300 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_271
timestamp 1644511149
transform 1 0 26036 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_284
timestamp 1644511149
transform 1 0 27232 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_290
timestamp 1644511149
transform 1 0 27784 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_302
timestamp 1644511149
transform 1 0 28888 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_308
timestamp 1644511149
transform 1 0 29440 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_311
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_327
timestamp 1644511149
transform 1 0 31188 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_345
timestamp 1644511149
transform 1 0 32844 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_351
timestamp 1644511149
transform 1 0 33396 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_354
timestamp 1644511149
transform 1 0 33672 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_360
timestamp 1644511149
transform 1 0 34224 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_363
timestamp 1644511149
transform 1 0 34500 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_369
timestamp 1644511149
transform 1 0 35052 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_381
timestamp 1644511149
transform 1 0 36156 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_384
timestamp 1644511149
transform 1 0 36432 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_401
timestamp 1644511149
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_408
timestamp 1644511149
transform 1 0 38640 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_416
timestamp 1644511149
transform 1 0 39376 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_422
timestamp 1644511149
transform 1 0 39928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_425
timestamp 1644511149
transform 1 0 40204 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_431
timestamp 1644511149
transform 1 0 40756 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_435
timestamp 1644511149
transform 1 0 41124 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_438
timestamp 1644511149
transform 1 0 41400 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_446
timestamp 1644511149
transform 1 0 42136 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_451
timestamp 1644511149
transform 1 0 42596 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_469
timestamp 1644511149
transform 1 0 44252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_7
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_11
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_16
timestamp 1644511149
transform 1 0 2576 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_23
timestamp 1644511149
transform 1 0 3220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_33
timestamp 1644511149
transform 1 0 4140 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_43
timestamp 1644511149
transform 1 0 5060 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_51
timestamp 1644511149
transform 1 0 5796 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_56
timestamp 1644511149
transform 1 0 6256 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_64
timestamp 1644511149
transform 1 0 6992 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_69
timestamp 1644511149
transform 1 0 7452 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_75
timestamp 1644511149
transform 1 0 8004 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_89
timestamp 1644511149
transform 1 0 9292 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_95
timestamp 1644511149
transform 1 0 9844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_101
timestamp 1644511149
transform 1 0 10396 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_107
timestamp 1644511149
transform 1 0 10948 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_113
timestamp 1644511149
transform 1 0 11500 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_125
timestamp 1644511149
transform 1 0 12604 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1644511149
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_148
timestamp 1644511149
transform 1 0 14720 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_156
timestamp 1644511149
transform 1 0 15456 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_161
timestamp 1644511149
transform 1 0 15916 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_169
timestamp 1644511149
transform 1 0 16652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_174
timestamp 1644511149
transform 1 0 17112 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_178
timestamp 1644511149
transform 1 0 17480 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_183
timestamp 1644511149
transform 1 0 17940 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_191
timestamp 1644511149
transform 1 0 18676 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_201
timestamp 1644511149
transform 1 0 19596 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_215
timestamp 1644511149
transform 1 0 20884 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_227
timestamp 1644511149
transform 1 0 21988 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_235
timestamp 1644511149
transform 1 0 22724 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_240
timestamp 1644511149
transform 1 0 23184 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_246
timestamp 1644511149
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_257
timestamp 1644511149
transform 1 0 24748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_261
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_266
timestamp 1644511149
transform 1 0 25576 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_272
timestamp 1644511149
transform 1 0 26128 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_280
timestamp 1644511149
transform 1 0 26864 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_288
timestamp 1644511149
transform 1 0 27600 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_293
timestamp 1644511149
transform 1 0 28060 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_299
timestamp 1644511149
transform 1 0 28612 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_313
timestamp 1644511149
transform 1 0 29900 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_327
timestamp 1644511149
transform 1 0 31188 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_332
timestamp 1644511149
transform 1 0 31648 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_338
timestamp 1644511149
transform 1 0 32200 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_346
timestamp 1644511149
transform 1 0 32936 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_349
timestamp 1644511149
transform 1 0 33212 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_359
timestamp 1644511149
transform 1 0 34132 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_372
timestamp 1644511149
transform 1 0 35328 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_378
timestamp 1644511149
transform 1 0 35880 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_384
timestamp 1644511149
transform 1 0 36432 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_390
timestamp 1644511149
transform 1 0 36984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_393
timestamp 1644511149
transform 1 0 37260 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_405
timestamp 1644511149
transform 1 0 38364 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_425
timestamp 1644511149
transform 1 0 40204 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_437
timestamp 1644511149
transform 1 0 41308 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_443
timestamp 1644511149
transform 1 0 41860 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_449
timestamp 1644511149
transform 1 0 42412 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_7
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_25
timestamp 1644511149
transform 1 0 3404 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_33
timestamp 1644511149
transform 1 0 4140 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_38
timestamp 1644511149
transform 1 0 4600 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_44
timestamp 1644511149
transform 1 0 5152 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_65
timestamp 1644511149
transform 1 0 7084 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_73
timestamp 1644511149
transform 1 0 7820 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_78
timestamp 1644511149
transform 1 0 8280 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_86
timestamp 1644511149
transform 1 0 9016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_91
timestamp 1644511149
transform 1 0 9476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_99
timestamp 1644511149
transform 1 0 10212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_103
timestamp 1644511149
transform 1 0 10580 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1644511149
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_117
timestamp 1644511149
transform 1 0 11868 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_135
timestamp 1644511149
transform 1 0 13524 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_139
timestamp 1644511149
transform 1 0 13892 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_144
timestamp 1644511149
transform 1 0 14352 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_158
timestamp 1644511149
transform 1 0 15640 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1644511149
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_171
timestamp 1644511149
transform 1 0 16836 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_185
timestamp 1644511149
transform 1 0 18124 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_191
timestamp 1644511149
transform 1 0 18676 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_196
timestamp 1644511149
transform 1 0 19136 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_200
timestamp 1644511149
transform 1 0 19504 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_211
timestamp 1644511149
transform 1 0 20516 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_219
timestamp 1644511149
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_229
timestamp 1644511149
transform 1 0 22172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_257
timestamp 1644511149
transform 1 0 24748 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_262
timestamp 1644511149
transform 1 0 25208 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_270
timestamp 1644511149
transform 1 0 25944 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 1644511149
transform 1 0 26404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_288
timestamp 1644511149
transform 1 0 27600 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_294
timestamp 1644511149
transform 1 0 28152 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_302
timestamp 1644511149
transform 1 0 28888 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_310
timestamp 1644511149
transform 1 0 29624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_315
timestamp 1644511149
transform 1 0 30084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_323
timestamp 1644511149
transform 1 0 30820 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_331
timestamp 1644511149
transform 1 0 31556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_341
timestamp 1644511149
transform 1 0 32476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_353
timestamp 1644511149
transform 1 0 33580 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_358
timestamp 1644511149
transform 1 0 34040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_362
timestamp 1644511149
transform 1 0 34408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_367
timestamp 1644511149
transform 1 0 34868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_375
timestamp 1644511149
transform 1 0 35604 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_380
timestamp 1644511149
transform 1 0 36064 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1644511149
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_397
timestamp 1644511149
transform 1 0 37628 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_411
timestamp 1644511149
transform 1 0 38916 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_415
timestamp 1644511149
transform 1 0 39284 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_420
timestamp 1644511149
transform 1 0 39744 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_428
timestamp 1644511149
transform 1 0 40480 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_433
timestamp 1644511149
transform 1 0 40940 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_437
timestamp 1644511149
transform 1 0 41308 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_442
timestamp 1644511149
transform 1 0 41768 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_453
timestamp 1644511149
transform 1 0 42780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_469
timestamp 1644511149
transform 1 0 44252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_37
timestamp 1644511149
transform 1 0 4508 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_47
timestamp 1644511149
transform 1 0 5428 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_55
timestamp 1644511149
transform 1 0 6164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_73
timestamp 1644511149
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_79
timestamp 1644511149
transform 1 0 8372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_93
timestamp 1644511149
transform 1 0 9660 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_101
timestamp 1644511149
transform 1 0 10396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_105
timestamp 1644511149
transform 1 0 10764 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_108
timestamp 1644511149
transform 1 0 11040 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_117
timestamp 1644511149
transform 1 0 11868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_126
timestamp 1644511149
transform 1 0 12696 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_134
timestamp 1644511149
transform 1 0 13432 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_151
timestamp 1644511149
transform 1 0 14996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_159
timestamp 1644511149
transform 1 0 15732 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1644511149
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_179
timestamp 1644511149
transform 1 0 17572 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_187
timestamp 1644511149
transform 1 0 18308 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_207
timestamp 1644511149
transform 1 0 20148 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_213
timestamp 1644511149
transform 1 0 20700 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_218
timestamp 1644511149
transform 1 0 21160 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_261
timestamp 1644511149
transform 1 0 25116 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_271
timestamp 1644511149
transform 1 0 26036 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1644511149
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_297
timestamp 1644511149
transform 1 0 28428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_303
timestamp 1644511149
transform 1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_317
timestamp 1644511149
transform 1 0 30268 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_325
timestamp 1644511149
transform 1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_331
timestamp 1644511149
transform 1 0 31556 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1644511149
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_353
timestamp 1644511149
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_359
timestamp 1644511149
transform 1 0 34132 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_373
timestamp 1644511149
transform 1 0 35420 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_381
timestamp 1644511149
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_387
timestamp 1644511149
transform 1 0 36708 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1644511149
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_393
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_397
timestamp 1644511149
transform 1 0 37628 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_404
timestamp 1644511149
transform 1 0 38272 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_412
timestamp 1644511149
transform 1 0 39008 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_431
timestamp 1644511149
transform 1 0 40756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_441
timestamp 1644511149
transform 1 0 41676 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_447
timestamp 1644511149
transform 1 0 42228 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_453
timestamp 1644511149
transform 1 0 42780 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_461
timestamp 1644511149
transform 1 0 43516 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 44896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 44896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 44896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 44896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 44896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 44896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 44896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 44896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 44896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 44896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 44896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 44896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 44896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 44896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 44896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 44896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 44896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 44896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 44896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 44896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 44896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 44896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 44896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 44896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 44896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 44896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 44896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 44896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 44896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 44896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 44896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 44896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 44896 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 44896 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 44896 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 44896 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 44896 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 44896 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 44896 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 44896 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 44896 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 44896 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 44896 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 44896 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 44896 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 44896 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 44896 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 44896 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 44896 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 44896 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 44896 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 44896 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 44896 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 44896 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 44896 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 44896 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 44896 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 44896 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 44896 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 44896 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 44896 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 44896 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 44896 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 42320 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0397_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0398_
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0399_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0400_
timestamp 1644511149
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0401_
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0402_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0403_
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0404_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0405_
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _0406_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2392 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0407_
timestamp 1644511149
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0408_
timestamp 1644511149
transform -1 0 16192 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0409_
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0410_
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0411_
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0412_
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0413_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2392 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0414_
timestamp 1644511149
transform 1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0415_
timestamp 1644511149
transform -1 0 1656 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0416_
timestamp 1644511149
transform -1 0 11040 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0417_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4692 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0418_
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0419_
timestamp 1644511149
transform 1 0 9476 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0420_
timestamp 1644511149
transform 1 0 1472 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0421_
timestamp 1644511149
transform 1 0 2392 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0422_
timestamp 1644511149
transform -1 0 18492 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0423_
timestamp 1644511149
transform -1 0 12144 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0424_
timestamp 1644511149
transform 1 0 1472 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0425_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1644511149
transform 1 0 8372 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0428_
timestamp 1644511149
transform 1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0429_
timestamp 1644511149
transform 1 0 5612 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0430_
timestamp 1644511149
transform -1 0 19412 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0431_
timestamp 1644511149
transform -1 0 4048 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0432_
timestamp 1644511149
transform -1 0 9476 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0433_
timestamp 1644511149
transform -1 0 3312 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0434_
timestamp 1644511149
transform -1 0 2116 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0435_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0436_
timestamp 1644511149
transform -1 0 19780 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0437_
timestamp 1644511149
transform -1 0 9844 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0438_
timestamp 1644511149
transform 1 0 8188 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0439_
timestamp 1644511149
transform 1 0 9476 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0440_
timestamp 1644511149
transform -1 0 10028 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0441_
timestamp 1644511149
transform -1 0 12512 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1644511149
transform -1 0 13432 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1644511149
transform -1 0 14904 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0444_
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0445_
timestamp 1644511149
transform 1 0 16560 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0446_
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0447_
timestamp 1644511149
transform -1 0 10948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0448_
timestamp 1644511149
transform -1 0 20240 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1644511149
transform 1 0 18584 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0450_
timestamp 1644511149
transform -1 0 2024 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1644511149
transform 1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0452_
timestamp 1644511149
transform -1 0 19780 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0453_
timestamp 1644511149
transform -1 0 4692 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0454_
timestamp 1644511149
transform -1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1644511149
transform -1 0 1748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1644511149
transform -1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0458_
timestamp 1644511149
transform -1 0 20700 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0459_
timestamp 1644511149
transform -1 0 12420 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0460_
timestamp 1644511149
transform 1 0 13064 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0461_
timestamp 1644511149
transform 1 0 17848 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0462_
timestamp 1644511149
transform -1 0 20700 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0463_
timestamp 1644511149
transform -1 0 4784 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0464_
timestamp 1644511149
transform 1 0 21068 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1644511149
transform 1 0 23644 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0466_
timestamp 1644511149
transform 1 0 9108 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0467_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1644511149
transform 1 0 3956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1644511149
transform -1 0 7544 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1644511149
transform 1 0 3036 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1644511149
transform 1 0 6624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0472_
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0473_
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0474_
timestamp 1644511149
transform 1 0 4140 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1644511149
transform -1 0 5888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0476_
timestamp 1644511149
transform -1 0 2852 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1644511149
transform 1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0478_
timestamp 1644511149
transform 1 0 9108 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0479_
timestamp 1644511149
transform -1 0 2392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0480_
timestamp 1644511149
transform 1 0 7912 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0481_
timestamp 1644511149
transform 1 0 9568 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1644511149
transform 1 0 4968 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1644511149
transform -1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0484_
timestamp 1644511149
transform -1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0485_
timestamp 1644511149
transform -1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0486_
timestamp 1644511149
transform 1 0 5336 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0487_
timestamp 1644511149
transform 1 0 7544 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0488_
timestamp 1644511149
transform 1 0 10120 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1644511149
transform -1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0490_
timestamp 1644511149
transform 1 0 6532 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0491_
timestamp 1644511149
transform 1 0 8280 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0492_
timestamp 1644511149
transform 1 0 5520 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0493_
timestamp 1644511149
transform -1 0 6164 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0494_
timestamp 1644511149
transform -1 0 4692 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0495_
timestamp 1644511149
transform 1 0 15272 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0496_
timestamp 1644511149
transform 1 0 3220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0497_
timestamp 1644511149
transform -1 0 4048 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0498_
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0499_
timestamp 1644511149
transform 1 0 3128 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0500_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20516 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0501_
timestamp 1644511149
transform -1 0 17204 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0502_
timestamp 1644511149
transform -1 0 22264 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0503_
timestamp 1644511149
transform -1 0 17664 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0504_
timestamp 1644511149
transform -1 0 23092 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0505_
timestamp 1644511149
transform -1 0 19504 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0506_
timestamp 1644511149
transform -1 0 23920 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0507_
timestamp 1644511149
transform -1 0 20884 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0508_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20056 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0509_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0510_
timestamp 1644511149
transform 1 0 21896 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0511_
timestamp 1644511149
transform 1 0 13156 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0512_
timestamp 1644511149
transform 1 0 19872 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0513_
timestamp 1644511149
transform 1 0 16928 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0514_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0515_
timestamp 1644511149
transform -1 0 13616 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0516_
timestamp 1644511149
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0517_
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0518_
timestamp 1644511149
transform 1 0 21988 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0519_
timestamp 1644511149
transform -1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0520_
timestamp 1644511149
transform 1 0 18032 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0521_
timestamp 1644511149
transform 1 0 24472 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0522_
timestamp 1644511149
transform 1 0 18308 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0523_
timestamp 1644511149
transform 1 0 25208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0524_
timestamp 1644511149
transform 1 0 21620 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0525_
timestamp 1644511149
transform 1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0526_
timestamp 1644511149
transform 1 0 20792 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0527_
timestamp 1644511149
transform 1 0 20884 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0528_
timestamp 1644511149
transform 1 0 27508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0529_
timestamp 1644511149
transform -1 0 21252 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0530_
timestamp 1644511149
transform 1 0 28428 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0531_
timestamp 1644511149
transform -1 0 22080 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0532_
timestamp 1644511149
transform 1 0 29900 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0533_
timestamp 1644511149
transform -1 0 23000 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0534_
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0535_
timestamp 1644511149
transform -1 0 23920 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0536_
timestamp 1644511149
transform 1 0 32476 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0537_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20700 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0538_
timestamp 1644511149
transform 1 0 15640 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0539_
timestamp 1644511149
transform -1 0 17296 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0540_
timestamp 1644511149
transform 1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0541_
timestamp 1644511149
transform -1 0 17664 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0542_
timestamp 1644511149
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0543_
timestamp 1644511149
transform -1 0 18584 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0544_
timestamp 1644511149
transform 1 0 15456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0545_
timestamp 1644511149
transform -1 0 19504 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0546_
timestamp 1644511149
transform 1 0 16100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0547_
timestamp 1644511149
transform -1 0 22540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0548_
timestamp 1644511149
transform -1 0 22908 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1644511149
transform 1 0 17204 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0550_
timestamp 1644511149
transform -1 0 23828 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0551_
timestamp 1644511149
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0552_
timestamp 1644511149
transform -1 0 23644 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1644511149
transform 1 0 20424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0554_
timestamp 1644511149
transform 1 0 24656 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1644511149
transform 1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0556_
timestamp 1644511149
transform -1 0 23460 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1644511149
transform -1 0 21804 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0558_
timestamp 1644511149
transform -1 0 24380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 1644511149
transform 1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0560_
timestamp 1644511149
transform -1 0 25300 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0562_
timestamp 1644511149
transform 1 0 27140 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0564_
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0565_
timestamp 1644511149
transform 1 0 11408 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1644511149
transform -1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0567_
timestamp 1644511149
transform 1 0 9844 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0568_
timestamp 1644511149
transform -1 0 18952 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0569_
timestamp 1644511149
transform 1 0 17848 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0570_
timestamp 1644511149
transform 1 0 19320 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0571_
timestamp 1644511149
transform -1 0 19596 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0572_
timestamp 1644511149
transform -1 0 18768 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0573_
timestamp 1644511149
transform 1 0 12696 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0574_
timestamp 1644511149
transform -1 0 20148 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0575_
timestamp 1644511149
transform 1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0576_
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0577_
timestamp 1644511149
transform 1 0 22080 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0578_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0579_
timestamp 1644511149
transform 1 0 22172 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0580_
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0581_
timestamp 1644511149
transform 1 0 22356 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0582_
timestamp 1644511149
transform 1 0 21896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0583_
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0584_
timestamp 1644511149
transform 1 0 23368 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0585_
timestamp 1644511149
transform 1 0 15364 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0586_
timestamp 1644511149
transform 1 0 22448 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0587_
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0588_
timestamp 1644511149
transform 1 0 23552 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0589_
timestamp 1644511149
transform 1 0 17204 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0590_
timestamp 1644511149
transform 1 0 24656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0591_
timestamp 1644511149
transform 1 0 17664 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0592_
timestamp 1644511149
transform 1 0 25852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0593_
timestamp 1644511149
transform 1 0 19228 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0594_
timestamp 1644511149
transform 1 0 27508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0595_
timestamp 1644511149
transform -1 0 17756 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0596_
timestamp 1644511149
transform -1 0 6808 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0597_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11408 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0598_
timestamp 1644511149
transform -1 0 6624 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0599_
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0600_
timestamp 1644511149
transform -1 0 6164 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0601_
timestamp 1644511149
transform 1 0 11316 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0602_
timestamp 1644511149
transform -1 0 5888 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0603_
timestamp 1644511149
transform 1 0 11592 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0604_
timestamp 1644511149
transform -1 0 8280 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 1644511149
transform 1 0 12604 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0606_
timestamp 1644511149
transform -1 0 8924 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0607_
timestamp 1644511149
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0608_
timestamp 1644511149
transform -1 0 13616 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0609_
timestamp 1644511149
transform -1 0 13984 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0610_
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0611_
timestamp 1644511149
transform -1 0 13800 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0612_
timestamp 1644511149
transform -1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0613_
timestamp 1644511149
transform 1 0 17848 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0614_
timestamp 1644511149
transform -1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0615_
timestamp 1644511149
transform -1 0 15272 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0616_
timestamp 1644511149
transform 1 0 14444 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0617_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0618_
timestamp 1644511149
transform 1 0 15364 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0619_
timestamp 1644511149
transform -1 0 15824 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0620_
timestamp 1644511149
transform 1 0 16468 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0621_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1644511149
transform 1 0 17572 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0623_
timestamp 1644511149
transform -1 0 18216 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0624_
timestamp 1644511149
transform -1 0 19596 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0625_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0627_
timestamp 1644511149
transform -1 0 20976 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0628_
timestamp 1644511149
transform 1 0 15548 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0629_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _0630_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 11040 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0631_
timestamp 1644511149
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0632_
timestamp 1644511149
transform -1 0 12144 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0633_
timestamp 1644511149
transform 1 0 18216 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0634_
timestamp 1644511149
transform -1 0 13616 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0635_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0636_
timestamp 1644511149
transform -1 0 13340 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0637_
timestamp 1644511149
transform 1 0 22172 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0638_
timestamp 1644511149
transform -1 0 14168 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0639_
timestamp 1644511149
transform 1 0 22172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0640_
timestamp 1644511149
transform -1 0 15088 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0641_
timestamp 1644511149
transform 1 0 23184 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0642_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0643_
timestamp 1644511149
transform 1 0 25576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0644_
timestamp 1644511149
transform -1 0 16560 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0645_
timestamp 1644511149
transform 1 0 25116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0646_
timestamp 1644511149
transform 1 0 20700 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0647_
timestamp 1644511149
transform 1 0 27324 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0648_
timestamp 1644511149
transform -1 0 17664 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0649_
timestamp 1644511149
transform 1 0 27048 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0650_
timestamp 1644511149
transform -1 0 18768 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0651_
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0652_
timestamp 1644511149
transform -1 0 20056 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0653_
timestamp 1644511149
transform 1 0 29072 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0654_
timestamp 1644511149
transform -1 0 20332 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0655_
timestamp 1644511149
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _0656_
timestamp 1644511149
transform -1 0 21160 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0657_
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0658_
timestamp 1644511149
transform -1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0659_
timestamp 1644511149
transform -1 0 6808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0660_
timestamp 1644511149
transform -1 0 19872 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0661_
timestamp 1644511149
transform -1 0 13616 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0662_
timestamp 1644511149
transform -1 0 20240 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0663_
timestamp 1644511149
transform -1 0 14996 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0664_
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0665_
timestamp 1644511149
transform 1 0 20608 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0666_
timestamp 1644511149
transform -1 0 19320 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0667_
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0668_
timestamp 1644511149
transform 1 0 20240 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0669_
timestamp 1644511149
transform 1 0 26772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0670_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 14720 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0671_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10580 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0672_
timestamp 1644511149
transform -1 0 16560 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0673_
timestamp 1644511149
transform 1 0 15732 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0674_
timestamp 1644511149
transform -1 0 18400 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0675_
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0676_
timestamp 1644511149
transform 1 0 15180 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0677_
timestamp 1644511149
transform -1 0 20424 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0678_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18768 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0679_
timestamp 1644511149
transform 1 0 12788 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0680_
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0681_
timestamp 1644511149
transform -1 0 19872 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0682_
timestamp 1644511149
transform 1 0 6256 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0683_
timestamp 1644511149
transform 1 0 2392 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0684_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0685_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0686_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0687_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19136 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0688_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0689_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16836 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0690_
timestamp 1644511149
transform -1 0 4140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0691_
timestamp 1644511149
transform -1 0 15364 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0692_
timestamp 1644511149
transform -1 0 4876 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0693_
timestamp 1644511149
transform -1 0 16192 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0694_
timestamp 1644511149
transform -1 0 4600 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0695_
timestamp 1644511149
transform -1 0 15180 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0696_
timestamp 1644511149
transform -1 0 12144 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0697_
timestamp 1644511149
transform -1 0 18584 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0698_
timestamp 1644511149
transform -1 0 10212 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0699_
timestamp 1644511149
transform -1 0 18216 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0700_
timestamp 1644511149
transform -1 0 14260 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0701_
timestamp 1644511149
transform -1 0 17388 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0702_
timestamp 1644511149
transform -1 0 15548 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0703_
timestamp 1644511149
transform -1 0 18492 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0704_
timestamp 1644511149
transform -1 0 16284 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0705_
timestamp 1644511149
transform -1 0 22264 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0706_
timestamp 1644511149
transform -1 0 16284 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0707_
timestamp 1644511149
transform -1 0 18952 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0708_
timestamp 1644511149
transform -1 0 15732 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1644511149
transform -1 0 18400 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0710_
timestamp 1644511149
transform -1 0 18768 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0711_
timestamp 1644511149
transform 1 0 14536 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0712_
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0713_
timestamp 1644511149
transform 1 0 20148 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0714_
timestamp 1644511149
transform -1 0 3312 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _0715_
timestamp 1644511149
transform 1 0 20148 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0716_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15088 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0717_
timestamp 1644511149
transform -1 0 22632 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0718_
timestamp 1644511149
transform -1 0 22356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0719_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0720_
timestamp 1644511149
transform 1 0 6992 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0721_
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0722_
timestamp 1644511149
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 1644511149
transform 1 0 24104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0724_
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0725_
timestamp 1644511149
transform 1 0 10304 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0726_
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0727_
timestamp 1644511149
transform 1 0 10580 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0728_
timestamp 1644511149
transform 1 0 10488 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0729_
timestamp 1644511149
transform -1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0730_
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0731_
timestamp 1644511149
transform 1 0 20240 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0732_
timestamp 1644511149
transform 1 0 25024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0733_
timestamp 1644511149
transform 1 0 19504 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0734_
timestamp 1644511149
transform -1 0 10672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0735_
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0736_
timestamp 1644511149
transform 1 0 21068 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0737_
timestamp 1644511149
transform -1 0 11316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0738_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0739_
timestamp 1644511149
transform -1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0740_
timestamp 1644511149
transform 1 0 18492 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0741_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0742_
timestamp 1644511149
transform 1 0 23368 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0743_
timestamp 1644511149
transform -1 0 6624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0744_
timestamp 1644511149
transform 1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0745_
timestamp 1644511149
transform -1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0746_
timestamp 1644511149
transform 1 0 21252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0747_
timestamp 1644511149
transform -1 0 23460 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0748_
timestamp 1644511149
transform -1 0 3312 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0749_
timestamp 1644511149
transform 1 0 10120 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0750_
timestamp 1644511149
transform -1 0 2760 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0751_
timestamp 1644511149
transform -1 0 10948 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0752_
timestamp 1644511149
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0753_
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0754_
timestamp 1644511149
transform 1 0 13616 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0755_
timestamp 1644511149
transform 1 0 21528 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0756_
timestamp 1644511149
transform -1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0757_
timestamp 1644511149
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0758_
timestamp 1644511149
transform 1 0 23184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0759_
timestamp 1644511149
transform -1 0 16560 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0760_
timestamp 1644511149
transform 1 0 11684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0761_
timestamp 1644511149
transform 1 0 17848 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0762_
timestamp 1644511149
transform -1 0 19780 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0763_
timestamp 1644511149
transform -1 0 12788 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0764_
timestamp 1644511149
transform 1 0 13248 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 1644511149
transform -1 0 13800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0766_
timestamp 1644511149
transform -1 0 20976 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0767_
timestamp 1644511149
transform -1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0768_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0769_
timestamp 1644511149
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0770_
timestamp 1644511149
transform -1 0 13524 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0771_
timestamp 1644511149
transform 1 0 22632 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0772_
timestamp 1644511149
transform 1 0 20608 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0773_
timestamp 1644511149
transform 1 0 20148 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _0774_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 14536 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_2  _0775_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2760 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0776_
timestamp 1644511149
transform 1 0 9936 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0777_
timestamp 1644511149
transform 1 0 5520 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1644511149
transform -1 0 8464 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0779_
timestamp 1644511149
transform 1 0 8004 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0780_
timestamp 1644511149
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0781_
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1644511149
transform -1 0 5888 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0783_
timestamp 1644511149
transform -1 0 7544 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0784_
timestamp 1644511149
transform -1 0 7544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1644511149
transform 1 0 8372 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0786_
timestamp 1644511149
transform 1 0 4416 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0787_
timestamp 1644511149
transform 1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1644511149
transform 1 0 4048 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0789_
timestamp 1644511149
transform 1 0 2300 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0790_
timestamp 1644511149
transform -1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1644511149
transform 1 0 8924 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0792_
timestamp 1644511149
transform 1 0 1472 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0793_
timestamp 1644511149
transform -1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0794_
timestamp 1644511149
transform -1 0 4048 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1644511149
transform -1 0 7268 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0796_
timestamp 1644511149
transform -1 0 9844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0797_
timestamp 1644511149
transform -1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0798_
timestamp 1644511149
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0799_
timestamp 1644511149
transform -1 0 4048 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0800_
timestamp 1644511149
transform 1 0 4600 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0801_
timestamp 1644511149
transform -1 0 6256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0802_
timestamp 1644511149
transform 1 0 5060 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0803_
timestamp 1644511149
transform 1 0 2760 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0804_
timestamp 1644511149
transform -1 0 5244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1644511149
transform 1 0 13432 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0806_
timestamp 1644511149
transform -1 0 9660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0807_
timestamp 1644511149
transform -1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1644511149
transform -1 0 3312 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0809_
timestamp 1644511149
transform 1 0 7912 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0810_
timestamp 1644511149
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0811_
timestamp 1644511149
transform 1 0 22172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp 1644511149
transform -1 0 16192 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0813_
timestamp 1644511149
transform 1 0 17572 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0814_
timestamp 1644511149
transform 1 0 23368 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0815_
timestamp 1644511149
transform 1 0 25024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1644511149
transform -1 0 2208 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0817_
timestamp 1644511149
transform 1 0 14996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0818_
timestamp 1644511149
transform 1 0 25668 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0819_
timestamp 1644511149
transform -1 0 19320 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0820_
timestamp 1644511149
transform 1 0 21068 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0821_
timestamp 1644511149
transform 1 0 21528 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0822_
timestamp 1644511149
transform -1 0 16744 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0823_
timestamp 1644511149
transform 1 0 21988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0824_
timestamp 1644511149
transform 1 0 22172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0826_
timestamp 1644511149
transform 1 0 12328 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0827_
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0828_
timestamp 1644511149
transform 1 0 20148 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 1644511149
transform -1 0 2208 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0830_
timestamp 1644511149
transform 1 0 21988 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0831_
timestamp 1644511149
transform 1 0 24288 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0832_
timestamp 1644511149
transform -1 0 9200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0833_
timestamp 1644511149
transform -1 0 17480 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0834_
timestamp 1644511149
transform -1 0 22356 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0835_
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0836_
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0837_
timestamp 1644511149
transform 1 0 9384 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0838_
timestamp 1644511149
transform -1 0 11592 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0839_
timestamp 1644511149
transform -1 0 11040 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0840_
timestamp 1644511149
transform 1 0 10764 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0841_
timestamp 1644511149
transform 1 0 12880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 1644511149
transform 1 0 17848 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0843_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0844_
timestamp 1644511149
transform -1 0 13800 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0845_
timestamp 1644511149
transform -1 0 9384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0847_
timestamp 1644511149
transform 1 0 9016 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0848_
timestamp 1644511149
transform -1 0 14352 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 1644511149
transform -1 0 3312 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0851_
timestamp 1644511149
transform 1 0 2760 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0852_
timestamp 1644511149
transform -1 0 9844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp 1644511149
transform -1 0 4048 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0854_
timestamp 1644511149
transform 1 0 5244 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0855_
timestamp 1644511149
transform 1 0 6992 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 1644511149
transform 1 0 4508 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0857_
timestamp 1644511149
transform -1 0 4692 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0858_
timestamp 1644511149
transform -1 0 3036 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp 1644511149
transform 1 0 2024 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0860_
timestamp 1644511149
transform 1 0 1564 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0861_
timestamp 1644511149
transform -1 0 2392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0862_
timestamp 1644511149
transform 1 0 3404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0863_
timestamp 1644511149
transform -1 0 2760 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0864_
timestamp 1644511149
transform -1 0 7820 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0865_
timestamp 1644511149
transform -1 0 1748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0866_
timestamp 1644511149
transform 1 0 7728 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0867_
timestamp 1644511149
transform -1 0 7636 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0868_
timestamp 1644511149
transform -1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0869_
timestamp 1644511149
transform 1 0 4968 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0870_
timestamp 1644511149
transform -1 0 6992 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0871_
timestamp 1644511149
transform -1 0 6808 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1644511149
transform 1 0 4048 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0873_
timestamp 1644511149
transform 1 0 7176 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0874_
timestamp 1644511149
transform 1 0 5336 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0875_
timestamp 1644511149
transform 1 0 7728 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0876_
timestamp 1644511149
transform -1 0 3312 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0877_
timestamp 1644511149
transform 1 0 4324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0878_
timestamp 1644511149
transform 1 0 7084 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0879_
timestamp 1644511149
transform 1 0 5060 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0880_
timestamp 1644511149
transform 1 0 2760 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1644511149
transform 1 0 5612 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0882_
timestamp 1644511149
transform -1 0 13340 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0883_
timestamp 1644511149
transform -1 0 23276 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0884_
timestamp 1644511149
transform 1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _0885_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13800 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0886_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6992 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0887_
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0889_
timestamp 1644511149
transform 1 0 4416 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1644511149
transform 1 0 5152 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1644511149
transform 1 0 5060 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1644511149
transform 1 0 7084 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1644511149
transform 1 0 16008 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1644511149
transform -1 0 14904 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1644511149
transform 1 0 11224 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1644511149
transform 1 0 6440 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1644511149
transform 1 0 4416 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1644511149
transform -1 0 11040 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1644511149
transform -1 0 11316 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1644511149
transform -1 0 14812 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1644511149
transform 1 0 16008 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0909_
timestamp 1644511149
transform 1 0 14628 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0910_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0911_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0912_
timestamp 1644511149
transform 1 0 14076 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0913_
timestamp 1644511149
transform 1 0 4692 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0914_
timestamp 1644511149
transform 1 0 15916 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0915_
timestamp 1644511149
transform 1 0 6808 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0916_
timestamp 1644511149
transform 1 0 4416 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0917_
timestamp 1644511149
transform 1 0 11684 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0918_
timestamp 1644511149
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0919_
timestamp 1644511149
transform -1 0 13064 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0920_
timestamp 1644511149
transform 1 0 11224 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0921_
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0922_
timestamp 1644511149
transform 1 0 11224 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0923_
timestamp 1644511149
transform -1 0 13064 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0924_
timestamp 1644511149
transform -1 0 13064 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0925_
timestamp 1644511149
transform -1 0 14996 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0926_
timestamp 1644511149
transform -1 0 15640 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0927_
timestamp 1644511149
transform 1 0 6900 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0928_
timestamp 1644511149
transform -1 0 8740 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0929_
timestamp 1644511149
transform 1 0 6900 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0930_
timestamp 1644511149
transform 1 0 14628 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0931_
timestamp 1644511149
transform 1 0 6992 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0932_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0933_
timestamp 1644511149
transform 1 0 14076 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _0934_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11776 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1644511149
transform -1 0 6532 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1644511149
transform 1 0 4416 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1644511149
transform 1 0 4692 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1644511149
transform 1 0 4416 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1644511149
transform 1 0 4416 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1644511149
transform 1 0 2576 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1644511149
transform 1 0 6992 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1644511149
transform 1 0 4416 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1644511149
transform 1 0 2576 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1644511149
transform -1 0 18124 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0945__287 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0946__288
timestamp 1644511149
transform -1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0947__289
timestamp 1644511149
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0948__290
timestamp 1644511149
transform -1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0949__291
timestamp 1644511149
transform -1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0950__292
timestamp 1644511149
transform -1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0951_
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0952_
timestamp 1644511149
transform 1 0 23184 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0953_
timestamp 1644511149
transform 1 0 24748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0954_
timestamp 1644511149
transform 1 0 28428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0955_
timestamp 1644511149
transform 1 0 29900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0956_
timestamp 1644511149
transform -1 0 18492 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0957_
timestamp 1644511149
transform -1 0 25116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0958_
timestamp 1644511149
transform -1 0 27692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 1644511149
transform 1 0 26864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1644511149
transform 1 0 27876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0962_
timestamp 1644511149
transform -1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0963_
timestamp 1644511149
transform -1 0 29716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0964_
timestamp 1644511149
transform 1 0 32568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0965_
timestamp 1644511149
transform 1 0 33672 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0966_
timestamp 1644511149
transform 1 0 35052 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0967_
timestamp 1644511149
transform -1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0968_
timestamp 1644511149
transform -1 0 29256 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0969_
timestamp 1644511149
transform -1 0 31004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0970_
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0971_
timestamp 1644511149
transform 1 0 32936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0972_
timestamp 1644511149
transform 1 0 34132 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0973_
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_8  _0974_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0975_
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0976_
timestamp 1644511149
transform -1 0 10580 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0977_
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0978_
timestamp 1644511149
transform -1 0 10856 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0979_
timestamp 1644511149
transform 1 0 11224 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0980_
timestamp 1644511149
transform 1 0 8188 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0981_
timestamp 1644511149
transform -1 0 8464 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0982_
timestamp 1644511149
transform 1 0 6532 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0983_
timestamp 1644511149
transform -1 0 10856 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0984_
timestamp 1644511149
transform -1 0 10856 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0985_
timestamp 1644511149
transform -1 0 11132 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0986_
timestamp 1644511149
transform -1 0 11040 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0987_
timestamp 1644511149
transform -1 0 11408 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0988_
timestamp 1644511149
transform 1 0 8924 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0989_
timestamp 1644511149
transform -1 0 10856 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0990_
timestamp 1644511149
transform -1 0 10856 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0991_
timestamp 1644511149
transform -1 0 13432 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0992_
timestamp 1644511149
transform -1 0 11316 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0993_
timestamp 1644511149
transform -1 0 13156 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0994_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0995_
timestamp 1644511149
transform -1 0 11040 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0996_
timestamp 1644511149
transform -1 0 8464 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0997_
timestamp 1644511149
transform -1 0 8740 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0998_
timestamp 1644511149
transform -1 0 9108 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _0999_
timestamp 1644511149
transform 1 0 6532 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1000_
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1001_
timestamp 1644511149
transform -1 0 8556 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1002_
timestamp 1644511149
transform -1 0 9108 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1003_
timestamp 1644511149
transform 1 0 6532 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1004_
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1005_
timestamp 1644511149
transform -1 0 6164 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk
timestamp 1644511149
transform -1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 1644511149
transform -1 0 14444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_clk
timestamp 1644511149
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_clk
timestamp 1644511149
transform -1 0 11868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_clk
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_clk
timestamp 1644511149
transform 1 0 13892 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clk
timestamp 1644511149
transform 1 0 3864 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clk
timestamp 1644511149
transform 1 0 6532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clk
timestamp 1644511149
transform 1 0 2024 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clk
timestamp 1644511149
transform -1 0 12788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clk
timestamp 1644511149
transform -1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clk
timestamp 1644511149
transform -1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clk
timestamp 1644511149
transform -1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clk
timestamp 1644511149
transform -1 0 21988 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 2668 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 2668 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform -1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform -1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform -1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform -1 0 1656 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform -1 0 1656 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform -1 0 1656 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform -1 0 1656 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform -1 0 1656 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 2300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 2944 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 2024 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 2668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1644511149
transform -1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1644511149
transform -1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1644511149
transform 1 0 28152 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform -1 0 38272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform -1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1644511149
transform -1 0 41124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1644511149
transform -1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1644511149
transform -1 0 43884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform -1 0 44252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1644511149
transform -1 0 44252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1644511149
transform -1 0 44252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1644511149
transform -1 0 31188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1644511149
transform -1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform -1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1644511149
transform -1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform -1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1644511149
transform -1 0 36524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1644511149
transform -1 0 37628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform -1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1644511149
transform 1 0 28796 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1644511149
transform -1 0 39100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1644511149
transform -1 0 39836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform -1 0 40572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform -1 0 41860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform -1 0 43148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform -1 0 43516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform -1 0 43516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1644511149
transform -1 0 44252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform -1 0 44252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform -1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1644511149
transform -1 0 31188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform -1 0 32844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1644511149
transform -1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform -1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform -1 0 35052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1644511149
transform -1 0 35788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform -1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1644511149
transform -1 0 37720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform -1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1644511149
transform 1 0 20976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1644511149
transform 1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1644511149
transform 1 0 23736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1644511149
transform 1 0 25668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1644511149
transform 1 0 27508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1644511149
transform -1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1644511149
transform -1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1644511149
transform -1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1644511149
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1644511149
transform -1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1644511149
transform -1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1644511149
transform -1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1644511149
transform -1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1644511149
transform -1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1644511149
transform -1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1644511149
transform -1 0 20608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1644511149
transform 1 0 21252 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1644511149
transform 1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1644511149
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1644511149
transform 1 0 25024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input99
timestamp 1644511149
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1644511149
transform 1 0 26956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1644511149
transform 1 0 27876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1644511149
transform 1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1644511149
transform 1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1644511149
transform 1 0 14996 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1644511149
transform 1 0 15548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1644511149
transform -1 0 18676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1644511149
transform 1 0 19320 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input111
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1644511149
transform 1 0 12328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input113
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input114
timestamp 1644511149
transform -1 0 15640 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input115
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input116
timestamp 1644511149
transform 1 0 17204 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input117
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input118
timestamp 1644511149
transform 1 0 19596 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1644511149
transform 1 0 20792 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1644511149
transform 1 0 22172 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1644511149
transform -1 0 23644 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input122
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input123
timestamp 1644511149
transform -1 0 25116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1644511149
transform -1 0 26036 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input125
timestamp 1644511149
transform -1 0 27692 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input126
timestamp 1644511149
transform -1 0 28428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input127
timestamp 1644511149
transform -1 0 30268 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1644511149
transform -1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input129
timestamp 1644511149
transform -1 0 32844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1644511149
transform -1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input131
timestamp 1644511149
transform -1 0 35420 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input132
timestamp 1644511149
transform -1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input133
timestamp 1644511149
transform 1 0 2852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input134
timestamp 1644511149
transform -1 0 37628 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input135 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 38272 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input136
timestamp 1644511149
transform 1 0 40204 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input137
timestamp 1644511149
transform -1 0 41676 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input138
timestamp 1644511149
transform -1 0 41768 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input139
timestamp 1644511149
transform 1 0 4140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input140
timestamp 1644511149
transform 1 0 5060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input141
timestamp 1644511149
transform 1 0 6716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input142
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input143
timestamp 1644511149
transform 1 0 9292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input144
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input145
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1644511149
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input147
timestamp 1644511149
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input148
timestamp 1644511149
transform -1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1644511149
transform -1 0 9568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input150
timestamp 1644511149
transform -1 0 9568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input151
timestamp 1644511149
transform -1 0 10488 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input152
timestamp 1644511149
transform -1 0 10856 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input153
timestamp 1644511149
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input154
timestamp 1644511149
transform -1 0 6072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input155
timestamp 1644511149
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input156
timestamp 1644511149
transform -1 0 7360 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input157
timestamp 1644511149
transform -1 0 7636 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input158
timestamp 1644511149
transform -1 0 8004 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input159
timestamp 1644511149
transform -1 0 8924 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input160
timestamp 1644511149
transform -1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1644511149
transform -1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input162
timestamp 1644511149
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1644511149
transform -1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input164
timestamp 1644511149
transform -1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input165
timestamp 1644511149
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input166
timestamp 1644511149
transform -1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input167
timestamp 1644511149
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input168
timestamp 1644511149
transform -1 0 2300 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input169
timestamp 1644511149
transform -1 0 2300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input170
timestamp 1644511149
transform -1 0 3588 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform -1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform 1 0 38088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform -1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform 1 0 40940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1644511149
transform 1 0 41584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1644511149
transform 1 0 42320 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1644511149
transform 1 0 43884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1644511149
transform 1 0 30268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1644511149
transform 1 0 31004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1644511149
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1644511149
transform 1 0 33856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1644511149
transform 1 0 34776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1644511149
transform 1 0 35696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1644511149
transform 1 0 36616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1644511149
transform -1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1644511149
transform -1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1644511149
transform -1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1644511149
transform -1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1644511149
transform -1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1644511149
transform -1 0 25576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1644511149
transform -1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1644511149
transform -1 0 27600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1644511149
transform -1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1644511149
transform -1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1644511149
transform -1 0 13432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1644511149
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1644511149
transform -1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1644511149
transform -1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1644511149
transform -1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1644511149
transform -1 0 18584 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1644511149
transform -1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1644511149
transform -1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1644511149
transform -1 0 13432 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1644511149
transform -1 0 14352 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1644511149
transform 1 0 15364 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1644511149
transform 1 0 17940 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1644511149
transform 1 0 17572 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1644511149
transform -1 0 19136 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1644511149
transform -1 0 20332 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1644511149
transform -1 0 22172 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1644511149
transform -1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1644511149
transform 1 0 23644 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1644511149
transform -1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1644511149
transform -1 0 25208 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1644511149
transform 1 0 26036 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1644511149
transform 1 0 27232 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1644511149
transform 1 0 28520 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1644511149
transform 1 0 29716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1644511149
transform 1 0 31188 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1644511149
transform 1 0 33672 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1644511149
transform 1 0 34500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1644511149
transform -1 0 36064 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1644511149
transform -1 0 3404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1644511149
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1644511149
transform 1 0 38640 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1644511149
transform 1 0 39376 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1644511149
transform 1 0 42412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1644511149
transform 1 0 43884 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1644511149
transform 1 0 43884 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1644511149
transform 1 0 4232 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1644511149
transform -1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1644511149
transform -1 0 7084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1644511149
transform -1 0 8280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1644511149
transform -1 0 9476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1644511149
transform -1 0 11868 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1644511149
transform -1 0 12604 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1644511149
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1644511149
transform -1 0 13524 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1644511149
transform 1 0 14352 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1644511149
transform 1 0 15548 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1644511149
transform -1 0 17112 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1644511149
transform 1 0 18308 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1644511149
transform -1 0 19596 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1644511149
transform 1 0 20884 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1644511149
transform -1 0 21988 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1644511149
transform -1 0 23184 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1644511149
transform -1 0 2576 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1644511149
transform 1 0 25208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1644511149
transform 1 0 26496 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1644511149
transform -1 0 29900 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1644511149
transform 1 0 30452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1644511149
transform 1 0 31280 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1644511149
transform 1 0 32844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1644511149
transform 1 0 33764 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1644511149
transform 1 0 34960 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1644511149
transform 1 0 36432 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1644511149
transform -1 0 4140 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1644511149
transform 1 0 38732 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1644511149
transform 1 0 43148 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1644511149
transform 1 0 43884 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1644511149
transform 1 0 43884 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1644511149
transform -1 0 5060 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1644511149
transform -1 0 6256 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output280
timestamp 1644511149
transform -1 0 7452 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output281
timestamp 1644511149
transform -1 0 9292 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output282
timestamp 1644511149
transform -1 0 10212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output283
timestamp 1644511149
transform -1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output284
timestamp 1644511149
transform -1 0 12604 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output285
timestamp 1644511149
transform 1 0 43884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output286
timestamp 1644511149
transform 1 0 43884 0 -1 30464
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 280 800 400 6 clk
port 0 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 config_address[0]
port 1 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 config_address[10]
port 2 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 config_address[11]
port 3 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 config_address[12]
port 4 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 config_address[13]
port 5 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 config_address[14]
port 6 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 config_address[15]
port 7 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 config_address[16]
port 8 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 config_address[17]
port 9 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 config_address[18]
port 10 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 config_address[19]
port 11 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 config_address[1]
port 12 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 config_address[20]
port 13 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 config_address[21]
port 14 nsew signal input
rlabel metal3 s 0 28432 800 28552 6 config_address[22]
port 15 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 config_address[23]
port 16 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 config_address[24]
port 17 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 config_address[25]
port 18 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 config_address[26]
port 19 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 config_address[27]
port 20 nsew signal input
rlabel metal3 s 0 35504 800 35624 6 config_address[28]
port 21 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 config_address[29]
port 22 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 config_address[2]
port 23 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 config_address[30]
port 24 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 config_address[31]
port 25 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 config_address[3]
port 26 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 config_address[4]
port 27 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 config_address[5]
port 28 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 config_address[6]
port 29 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 config_address[7]
port 30 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 config_address[8]
port 31 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 config_address[9]
port 32 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 config_data[0]
port 33 nsew signal bidirectional
rlabel metal3 s 0 14968 800 15088 6 config_data[10]
port 34 nsew signal bidirectional
rlabel metal3 s 0 16056 800 16176 6 config_data[11]
port 35 nsew signal bidirectional
rlabel metal3 s 0 17280 800 17400 6 config_data[12]
port 36 nsew signal bidirectional
rlabel metal3 s 0 18504 800 18624 6 config_data[13]
port 37 nsew signal bidirectional
rlabel metal3 s 0 19592 800 19712 6 config_data[14]
port 38 nsew signal bidirectional
rlabel metal3 s 0 20816 800 20936 6 config_data[15]
port 39 nsew signal bidirectional
rlabel metal3 s 0 21904 800 22024 6 config_data[16]
port 40 nsew signal bidirectional
rlabel metal3 s 0 23128 800 23248 6 config_data[17]
port 41 nsew signal bidirectional
rlabel metal3 s 0 24352 800 24472 6 config_data[18]
port 42 nsew signal bidirectional
rlabel metal3 s 0 25440 800 25560 6 config_data[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 4360 800 4480 6 config_data[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 26664 800 26784 6 config_data[20]
port 45 nsew signal bidirectional
rlabel metal3 s 0 27888 800 28008 6 config_data[21]
port 46 nsew signal bidirectional
rlabel metal3 s 0 28976 800 29096 6 config_data[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 30200 800 30320 6 config_data[23]
port 48 nsew signal bidirectional
rlabel metal3 s 0 31424 800 31544 6 config_data[24]
port 49 nsew signal bidirectional
rlabel metal3 s 0 32512 800 32632 6 config_data[25]
port 50 nsew signal bidirectional
rlabel metal3 s 0 33736 800 33856 6 config_data[26]
port 51 nsew signal bidirectional
rlabel metal3 s 0 34960 800 35080 6 config_data[27]
port 52 nsew signal bidirectional
rlabel metal3 s 0 36048 800 36168 6 config_data[28]
port 53 nsew signal bidirectional
rlabel metal3 s 0 37272 800 37392 6 config_data[29]
port 54 nsew signal bidirectional
rlabel metal3 s 0 5448 800 5568 6 config_data[2]
port 55 nsew signal bidirectional
rlabel metal3 s 0 38496 800 38616 6 config_data[30]
port 56 nsew signal bidirectional
rlabel metal3 s 0 39584 800 39704 6 config_data[31]
port 57 nsew signal bidirectional
rlabel metal3 s 0 6672 800 6792 6 config_data[3]
port 58 nsew signal bidirectional
rlabel metal3 s 0 7896 800 8016 6 config_data[4]
port 59 nsew signal bidirectional
rlabel metal3 s 0 8984 800 9104 6 config_data[5]
port 60 nsew signal bidirectional
rlabel metal3 s 0 10208 800 10328 6 config_data[6]
port 61 nsew signal bidirectional
rlabel metal3 s 0 11432 800 11552 6 config_data[7]
port 62 nsew signal bidirectional
rlabel metal3 s 0 12520 800 12640 6 config_data[8]
port 63 nsew signal bidirectional
rlabel metal3 s 0 13744 800 13864 6 config_data[9]
port 64 nsew signal bidirectional
rlabel metal3 s 0 1368 800 1488 6 config_oe
port 65 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 config_we
port 66 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 gpio0_input[0]
port 67 nsew signal tristate
rlabel metal2 s 37554 0 37610 800 6 gpio0_input[10]
port 68 nsew signal tristate
rlabel metal2 s 38474 0 38530 800 6 gpio0_input[11]
port 69 nsew signal tristate
rlabel metal2 s 39486 0 39542 800 6 gpio0_input[12]
port 70 nsew signal tristate
rlabel metal2 s 40406 0 40462 800 6 gpio0_input[13]
port 71 nsew signal tristate
rlabel metal2 s 41326 0 41382 800 6 gpio0_input[14]
port 72 nsew signal tristate
rlabel metal2 s 42246 0 42302 800 6 gpio0_input[15]
port 73 nsew signal tristate
rlabel metal2 s 43258 0 43314 800 6 gpio0_input[16]
port 74 nsew signal tristate
rlabel metal2 s 44178 0 44234 800 6 gpio0_input[17]
port 75 nsew signal tristate
rlabel metal2 s 45098 0 45154 800 6 gpio0_input[18]
port 76 nsew signal tristate
rlabel metal2 s 29090 0 29146 800 6 gpio0_input[1]
port 77 nsew signal tristate
rlabel metal2 s 30010 0 30066 800 6 gpio0_input[2]
port 78 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 gpio0_input[3]
port 79 nsew signal tristate
rlabel metal2 s 31850 0 31906 800 6 gpio0_input[4]
port 80 nsew signal tristate
rlabel metal2 s 32862 0 32918 800 6 gpio0_input[5]
port 81 nsew signal tristate
rlabel metal2 s 33782 0 33838 800 6 gpio0_input[6]
port 82 nsew signal tristate
rlabel metal2 s 34702 0 34758 800 6 gpio0_input[7]
port 83 nsew signal tristate
rlabel metal2 s 35622 0 35678 800 6 gpio0_input[8]
port 84 nsew signal tristate
rlabel metal2 s 36634 0 36690 800 6 gpio0_input[9]
port 85 nsew signal tristate
rlabel metal2 s 28446 0 28502 800 6 gpio0_oe[0]
port 86 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 gpio0_oe[10]
port 87 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 gpio0_oe[11]
port 88 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 gpio0_oe[12]
port 89 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 gpio0_oe[13]
port 90 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 gpio0_oe[14]
port 91 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 gpio0_oe[15]
port 92 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 gpio0_oe[16]
port 93 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 gpio0_oe[17]
port 94 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 gpio0_oe[18]
port 95 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 gpio0_oe[1]
port 96 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 gpio0_oe[2]
port 97 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 gpio0_oe[3]
port 98 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 gpio0_oe[4]
port 99 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 gpio0_oe[5]
port 100 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 gpio0_oe[6]
port 101 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 gpio0_oe[7]
port 102 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 gpio0_oe[8]
port 103 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 gpio0_oe[9]
port 104 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 gpio0_output[0]
port 105 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 gpio0_output[10]
port 106 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 gpio0_output[11]
port 107 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 gpio0_output[12]
port 108 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 gpio0_output[13]
port 109 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 gpio0_output[14]
port 110 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 gpio0_output[15]
port 111 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 gpio0_output[16]
port 112 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 gpio0_output[17]
port 113 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 gpio0_output[18]
port 114 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 gpio0_output[1]
port 115 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 gpio0_output[2]
port 116 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 gpio0_output[3]
port 117 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 gpio0_output[4]
port 118 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 gpio0_output[5]
port 119 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 gpio0_output[6]
port 120 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 gpio0_output[7]
port 121 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 gpio0_output[8]
port 122 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 gpio0_output[9]
port 123 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 gpio1_input[0]
port 124 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 gpio1_input[10]
port 125 nsew signal tristate
rlabel metal2 s 20534 0 20590 800 6 gpio1_input[11]
port 126 nsew signal tristate
rlabel metal2 s 21454 0 21510 800 6 gpio1_input[12]
port 127 nsew signal tristate
rlabel metal2 s 22466 0 22522 800 6 gpio1_input[13]
port 128 nsew signal tristate
rlabel metal2 s 23386 0 23442 800 6 gpio1_input[14]
port 129 nsew signal tristate
rlabel metal2 s 24306 0 24362 800 6 gpio1_input[15]
port 130 nsew signal tristate
rlabel metal2 s 25226 0 25282 800 6 gpio1_input[16]
port 131 nsew signal tristate
rlabel metal2 s 26238 0 26294 800 6 gpio1_input[17]
port 132 nsew signal tristate
rlabel metal2 s 27158 0 27214 800 6 gpio1_input[18]
port 133 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 gpio1_input[1]
port 134 nsew signal tristate
rlabel metal2 s 12070 0 12126 800 6 gpio1_input[2]
port 135 nsew signal tristate
rlabel metal2 s 12990 0 13046 800 6 gpio1_input[3]
port 136 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 gpio1_input[4]
port 137 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 gpio1_input[5]
port 138 nsew signal tristate
rlabel metal2 s 15842 0 15898 800 6 gpio1_input[6]
port 139 nsew signal tristate
rlabel metal2 s 16762 0 16818 800 6 gpio1_input[7]
port 140 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 gpio1_input[8]
port 141 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 gpio1_input[9]
port 142 nsew signal tristate
rlabel metal2 s 10506 0 10562 800 6 gpio1_oe[0]
port 143 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 gpio1_oe[10]
port 144 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 gpio1_oe[11]
port 145 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 gpio1_oe[12]
port 146 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 gpio1_oe[13]
port 147 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 gpio1_oe[14]
port 148 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 gpio1_oe[15]
port 149 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 gpio1_oe[16]
port 150 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 gpio1_oe[17]
port 151 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 gpio1_oe[18]
port 152 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 gpio1_oe[1]
port 153 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 gpio1_oe[2]
port 154 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 gpio1_oe[3]
port 155 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 gpio1_oe[4]
port 156 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 gpio1_oe[5]
port 157 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 gpio1_oe[6]
port 158 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 gpio1_oe[7]
port 159 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 gpio1_oe[8]
port 160 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 gpio1_oe[9]
port 161 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 gpio1_output[0]
port 162 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 gpio1_output[10]
port 163 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 gpio1_output[11]
port 164 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 gpio1_output[12]
port 165 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 gpio1_output[13]
port 166 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 gpio1_output[14]
port 167 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 gpio1_output[15]
port 168 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 gpio1_output[16]
port 169 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 gpio1_output[17]
port 170 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 gpio1_output[18]
port 171 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 gpio1_output[1]
port 172 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 gpio1_output[2]
port 173 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 gpio1_output[3]
port 174 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 gpio1_output[4]
port 175 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 gpio1_output[5]
port 176 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 gpio1_output[6]
port 177 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 gpio1_output[7]
port 178 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 gpio1_output[8]
port 179 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 gpio1_output[9]
port 180 nsew signal input
rlabel metal2 s 202 39200 258 40000 6 io_in[0]
port 181 nsew signal input
rlabel metal2 s 12254 39200 12310 40000 6 io_in[10]
port 182 nsew signal input
rlabel metal2 s 13450 39200 13506 40000 6 io_in[11]
port 183 nsew signal input
rlabel metal2 s 14646 39200 14702 40000 6 io_in[12]
port 184 nsew signal input
rlabel metal2 s 15934 39200 15990 40000 6 io_in[13]
port 185 nsew signal input
rlabel metal2 s 17130 39200 17186 40000 6 io_in[14]
port 186 nsew signal input
rlabel metal2 s 18326 39200 18382 40000 6 io_in[15]
port 187 nsew signal input
rlabel metal2 s 19522 39200 19578 40000 6 io_in[16]
port 188 nsew signal input
rlabel metal2 s 20718 39200 20774 40000 6 io_in[17]
port 189 nsew signal input
rlabel metal2 s 21914 39200 21970 40000 6 io_in[18]
port 190 nsew signal input
rlabel metal2 s 23202 39200 23258 40000 6 io_in[19]
port 191 nsew signal input
rlabel metal2 s 1398 39200 1454 40000 6 io_in[1]
port 192 nsew signal input
rlabel metal2 s 24398 39200 24454 40000 6 io_in[20]
port 193 nsew signal input
rlabel metal2 s 25594 39200 25650 40000 6 io_in[21]
port 194 nsew signal input
rlabel metal2 s 26790 39200 26846 40000 6 io_in[22]
port 195 nsew signal input
rlabel metal2 s 27986 39200 28042 40000 6 io_in[23]
port 196 nsew signal input
rlabel metal2 s 29182 39200 29238 40000 6 io_in[24]
port 197 nsew signal input
rlabel metal2 s 30378 39200 30434 40000 6 io_in[25]
port 198 nsew signal input
rlabel metal2 s 31666 39200 31722 40000 6 io_in[26]
port 199 nsew signal input
rlabel metal2 s 32862 39200 32918 40000 6 io_in[27]
port 200 nsew signal input
rlabel metal2 s 34058 39200 34114 40000 6 io_in[28]
port 201 nsew signal input
rlabel metal2 s 35254 39200 35310 40000 6 io_in[29]
port 202 nsew signal input
rlabel metal2 s 2594 39200 2650 40000 6 io_in[2]
port 203 nsew signal input
rlabel metal2 s 36450 39200 36506 40000 6 io_in[30]
port 204 nsew signal input
rlabel metal2 s 37646 39200 37702 40000 6 io_in[31]
port 205 nsew signal input
rlabel metal2 s 38934 39200 38990 40000 6 io_in[32]
port 206 nsew signal input
rlabel metal2 s 40130 39200 40186 40000 6 io_in[33]
port 207 nsew signal input
rlabel metal2 s 41326 39200 41382 40000 6 io_in[34]
port 208 nsew signal input
rlabel metal2 s 42522 39200 42578 40000 6 io_in[35]
port 209 nsew signal input
rlabel metal2 s 43718 39200 43774 40000 6 io_in[36]
port 210 nsew signal input
rlabel metal2 s 44914 39200 44970 40000 6 io_in[37]
port 211 nsew signal input
rlabel metal2 s 3790 39200 3846 40000 6 io_in[3]
port 212 nsew signal input
rlabel metal2 s 4986 39200 5042 40000 6 io_in[4]
port 213 nsew signal input
rlabel metal2 s 6182 39200 6238 40000 6 io_in[5]
port 214 nsew signal input
rlabel metal2 s 7378 39200 7434 40000 6 io_in[6]
port 215 nsew signal input
rlabel metal2 s 8666 39200 8722 40000 6 io_in[7]
port 216 nsew signal input
rlabel metal2 s 9862 39200 9918 40000 6 io_in[8]
port 217 nsew signal input
rlabel metal2 s 11058 39200 11114 40000 6 io_in[9]
port 218 nsew signal input
rlabel metal2 s 570 39200 626 40000 6 io_oeb[0]
port 219 nsew signal tristate
rlabel metal2 s 12622 39200 12678 40000 6 io_oeb[10]
port 220 nsew signal tristate
rlabel metal2 s 13910 39200 13966 40000 6 io_oeb[11]
port 221 nsew signal tristate
rlabel metal2 s 15106 39200 15162 40000 6 io_oeb[12]
port 222 nsew signal tristate
rlabel metal2 s 16302 39200 16358 40000 6 io_oeb[13]
port 223 nsew signal tristate
rlabel metal2 s 17498 39200 17554 40000 6 io_oeb[14]
port 224 nsew signal tristate
rlabel metal2 s 18694 39200 18750 40000 6 io_oeb[15]
port 225 nsew signal tristate
rlabel metal2 s 19890 39200 19946 40000 6 io_oeb[16]
port 226 nsew signal tristate
rlabel metal2 s 21178 39200 21234 40000 6 io_oeb[17]
port 227 nsew signal tristate
rlabel metal2 s 22374 39200 22430 40000 6 io_oeb[18]
port 228 nsew signal tristate
rlabel metal2 s 23570 39200 23626 40000 6 io_oeb[19]
port 229 nsew signal tristate
rlabel metal2 s 1766 39200 1822 40000 6 io_oeb[1]
port 230 nsew signal tristate
rlabel metal2 s 24766 39200 24822 40000 6 io_oeb[20]
port 231 nsew signal tristate
rlabel metal2 s 25962 39200 26018 40000 6 io_oeb[21]
port 232 nsew signal tristate
rlabel metal2 s 27158 39200 27214 40000 6 io_oeb[22]
port 233 nsew signal tristate
rlabel metal2 s 28446 39200 28502 40000 6 io_oeb[23]
port 234 nsew signal tristate
rlabel metal2 s 29642 39200 29698 40000 6 io_oeb[24]
port 235 nsew signal tristate
rlabel metal2 s 30838 39200 30894 40000 6 io_oeb[25]
port 236 nsew signal tristate
rlabel metal2 s 32034 39200 32090 40000 6 io_oeb[26]
port 237 nsew signal tristate
rlabel metal2 s 33230 39200 33286 40000 6 io_oeb[27]
port 238 nsew signal tristate
rlabel metal2 s 34426 39200 34482 40000 6 io_oeb[28]
port 239 nsew signal tristate
rlabel metal2 s 35622 39200 35678 40000 6 io_oeb[29]
port 240 nsew signal tristate
rlabel metal2 s 2962 39200 3018 40000 6 io_oeb[2]
port 241 nsew signal tristate
rlabel metal2 s 36910 39200 36966 40000 6 io_oeb[30]
port 242 nsew signal tristate
rlabel metal2 s 38106 39200 38162 40000 6 io_oeb[31]
port 243 nsew signal tristate
rlabel metal2 s 39302 39200 39358 40000 6 io_oeb[32]
port 244 nsew signal tristate
rlabel metal2 s 40498 39200 40554 40000 6 io_oeb[33]
port 245 nsew signal tristate
rlabel metal2 s 41694 39200 41750 40000 6 io_oeb[34]
port 246 nsew signal tristate
rlabel metal2 s 42890 39200 42946 40000 6 io_oeb[35]
port 247 nsew signal tristate
rlabel metal2 s 44178 39200 44234 40000 6 io_oeb[36]
port 248 nsew signal tristate
rlabel metal2 s 45374 39200 45430 40000 6 io_oeb[37]
port 249 nsew signal tristate
rlabel metal2 s 4158 39200 4214 40000 6 io_oeb[3]
port 250 nsew signal tristate
rlabel metal2 s 5446 39200 5502 40000 6 io_oeb[4]
port 251 nsew signal tristate
rlabel metal2 s 6642 39200 6698 40000 6 io_oeb[5]
port 252 nsew signal tristate
rlabel metal2 s 7838 39200 7894 40000 6 io_oeb[6]
port 253 nsew signal tristate
rlabel metal2 s 9034 39200 9090 40000 6 io_oeb[7]
port 254 nsew signal tristate
rlabel metal2 s 10230 39200 10286 40000 6 io_oeb[8]
port 255 nsew signal tristate
rlabel metal2 s 11426 39200 11482 40000 6 io_oeb[9]
port 256 nsew signal tristate
rlabel metal2 s 938 39200 994 40000 6 io_out[0]
port 257 nsew signal tristate
rlabel metal2 s 13082 39200 13138 40000 6 io_out[10]
port 258 nsew signal tristate
rlabel metal2 s 14278 39200 14334 40000 6 io_out[11]
port 259 nsew signal tristate
rlabel metal2 s 15474 39200 15530 40000 6 io_out[12]
port 260 nsew signal tristate
rlabel metal2 s 16670 39200 16726 40000 6 io_out[13]
port 261 nsew signal tristate
rlabel metal2 s 17866 39200 17922 40000 6 io_out[14]
port 262 nsew signal tristate
rlabel metal2 s 19154 39200 19210 40000 6 io_out[15]
port 263 nsew signal tristate
rlabel metal2 s 20350 39200 20406 40000 6 io_out[16]
port 264 nsew signal tristate
rlabel metal2 s 21546 39200 21602 40000 6 io_out[17]
port 265 nsew signal tristate
rlabel metal2 s 22742 39200 22798 40000 6 io_out[18]
port 266 nsew signal tristate
rlabel metal2 s 23938 39200 23994 40000 6 io_out[19]
port 267 nsew signal tristate
rlabel metal2 s 2134 39200 2190 40000 6 io_out[1]
port 268 nsew signal tristate
rlabel metal2 s 25134 39200 25190 40000 6 io_out[20]
port 269 nsew signal tristate
rlabel metal2 s 26422 39200 26478 40000 6 io_out[21]
port 270 nsew signal tristate
rlabel metal2 s 27618 39200 27674 40000 6 io_out[22]
port 271 nsew signal tristate
rlabel metal2 s 28814 39200 28870 40000 6 io_out[23]
port 272 nsew signal tristate
rlabel metal2 s 30010 39200 30066 40000 6 io_out[24]
port 273 nsew signal tristate
rlabel metal2 s 31206 39200 31262 40000 6 io_out[25]
port 274 nsew signal tristate
rlabel metal2 s 32402 39200 32458 40000 6 io_out[26]
port 275 nsew signal tristate
rlabel metal2 s 33690 39200 33746 40000 6 io_out[27]
port 276 nsew signal tristate
rlabel metal2 s 34886 39200 34942 40000 6 io_out[28]
port 277 nsew signal tristate
rlabel metal2 s 36082 39200 36138 40000 6 io_out[29]
port 278 nsew signal tristate
rlabel metal2 s 3422 39200 3478 40000 6 io_out[2]
port 279 nsew signal tristate
rlabel metal2 s 37278 39200 37334 40000 6 io_out[30]
port 280 nsew signal tristate
rlabel metal2 s 38474 39200 38530 40000 6 io_out[31]
port 281 nsew signal tristate
rlabel metal2 s 39670 39200 39726 40000 6 io_out[32]
port 282 nsew signal tristate
rlabel metal2 s 40866 39200 40922 40000 6 io_out[33]
port 283 nsew signal tristate
rlabel metal2 s 42154 39200 42210 40000 6 io_out[34]
port 284 nsew signal tristate
rlabel metal2 s 43350 39200 43406 40000 6 io_out[35]
port 285 nsew signal tristate
rlabel metal2 s 44546 39200 44602 40000 6 io_out[36]
port 286 nsew signal tristate
rlabel metal2 s 45742 39200 45798 40000 6 io_out[37]
port 287 nsew signal tristate
rlabel metal2 s 4618 39200 4674 40000 6 io_out[3]
port 288 nsew signal tristate
rlabel metal2 s 5814 39200 5870 40000 6 io_out[4]
port 289 nsew signal tristate
rlabel metal2 s 7010 39200 7066 40000 6 io_out[5]
port 290 nsew signal tristate
rlabel metal2 s 8206 39200 8262 40000 6 io_out[6]
port 291 nsew signal tristate
rlabel metal2 s 9402 39200 9458 40000 6 io_out[7]
port 292 nsew signal tristate
rlabel metal2 s 10690 39200 10746 40000 6 io_out[8]
port 293 nsew signal tristate
rlabel metal2 s 11886 39200 11942 40000 6 io_out[9]
port 294 nsew signal tristate
rlabel metal3 s 45200 9936 46000 10056 6 la_blink[0]
port 295 nsew signal tristate
rlabel metal3 s 45200 29928 46000 30048 6 la_blink[1]
port 296 nsew signal tristate
rlabel metal2 s 5078 0 5134 800 6 pwm_out[0]
port 297 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 pwm_out[10]
port 298 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 pwm_out[11]
port 299 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 pwm_out[12]
port 300 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 pwm_out[13]
port 301 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 pwm_out[14]
port 302 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 pwm_out[15]
port 303 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 pwm_out[1]
port 304 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 pwm_out[2]
port 305 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 pwm_out[3]
port 306 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 pwm_out[4]
port 307 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 pwm_out[5]
port 308 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 pwm_out[6]
port 309 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 pwm_out[7]
port 310 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 pwm_out[8]
port 311 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 pwm_out[9]
port 312 nsew signal input
rlabel metal3 s 0 824 800 944 6 rst
port 313 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 spi_clk[0]
port 314 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 spi_clk[1]
port 315 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 spi_cs[0]
port 316 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 spi_cs[1]
port 317 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 spi_miso[0]
port 318 nsew signal tristate
rlabel metal2 s 4434 0 4490 800 6 spi_miso[1]
port 319 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 spi_mosi[0]
port 320 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 spi_mosi[1]
port 321 nsew signal input
rlabel metal2 s 110 0 166 800 6 uart_rx[0]
port 322 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 uart_rx[1]
port 323 nsew signal tristate
rlabel metal2 s 1306 0 1362 800 6 uart_rx[2]
port 324 nsew signal tristate
rlabel metal2 s 1950 0 2006 800 6 uart_rx[3]
port 325 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 uart_tx[0]
port 326 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 uart_tx[1]
port 327 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 uart_tx[2]
port 328 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 uart_tx[3]
port 329 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 330 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 330 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 331 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 46000 40000
<< end >>
