VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO WishboneInterconnect
  CLASS BLOCK ;
  FOREIGN WishboneInterconnect ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 1100.000 ;
  PIN master0_wb_ack_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END master0_wb_ack_i
  PIN master0_wb_adr_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END master0_wb_adr_o[0]
  PIN master0_wb_adr_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END master0_wb_adr_o[10]
  PIN master0_wb_adr_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END master0_wb_adr_o[11]
  PIN master0_wb_adr_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END master0_wb_adr_o[12]
  PIN master0_wb_adr_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END master0_wb_adr_o[13]
  PIN master0_wb_adr_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END master0_wb_adr_o[14]
  PIN master0_wb_adr_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END master0_wb_adr_o[15]
  PIN master0_wb_adr_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END master0_wb_adr_o[16]
  PIN master0_wb_adr_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END master0_wb_adr_o[17]
  PIN master0_wb_adr_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END master0_wb_adr_o[18]
  PIN master0_wb_adr_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END master0_wb_adr_o[19]
  PIN master0_wb_adr_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END master0_wb_adr_o[1]
  PIN master0_wb_adr_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END master0_wb_adr_o[20]
  PIN master0_wb_adr_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END master0_wb_adr_o[21]
  PIN master0_wb_adr_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END master0_wb_adr_o[22]
  PIN master0_wb_adr_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END master0_wb_adr_o[23]
  PIN master0_wb_adr_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END master0_wb_adr_o[24]
  PIN master0_wb_adr_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END master0_wb_adr_o[25]
  PIN master0_wb_adr_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END master0_wb_adr_o[26]
  PIN master0_wb_adr_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END master0_wb_adr_o[27]
  PIN master0_wb_adr_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END master0_wb_adr_o[2]
  PIN master0_wb_adr_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END master0_wb_adr_o[3]
  PIN master0_wb_adr_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END master0_wb_adr_o[4]
  PIN master0_wb_adr_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END master0_wb_adr_o[5]
  PIN master0_wb_adr_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END master0_wb_adr_o[6]
  PIN master0_wb_adr_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END master0_wb_adr_o[7]
  PIN master0_wb_adr_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END master0_wb_adr_o[8]
  PIN master0_wb_adr_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END master0_wb_adr_o[9]
  PIN master0_wb_cyc_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END master0_wb_cyc_o
  PIN master0_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END master0_wb_data_i[0]
  PIN master0_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END master0_wb_data_i[10]
  PIN master0_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END master0_wb_data_i[11]
  PIN master0_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END master0_wb_data_i[12]
  PIN master0_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END master0_wb_data_i[13]
  PIN master0_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END master0_wb_data_i[14]
  PIN master0_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END master0_wb_data_i[15]
  PIN master0_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END master0_wb_data_i[16]
  PIN master0_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END master0_wb_data_i[17]
  PIN master0_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END master0_wb_data_i[18]
  PIN master0_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END master0_wb_data_i[19]
  PIN master0_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END master0_wb_data_i[1]
  PIN master0_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END master0_wb_data_i[20]
  PIN master0_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END master0_wb_data_i[21]
  PIN master0_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END master0_wb_data_i[22]
  PIN master0_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END master0_wb_data_i[23]
  PIN master0_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END master0_wb_data_i[24]
  PIN master0_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END master0_wb_data_i[25]
  PIN master0_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END master0_wb_data_i[26]
  PIN master0_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END master0_wb_data_i[27]
  PIN master0_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END master0_wb_data_i[28]
  PIN master0_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END master0_wb_data_i[29]
  PIN master0_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END master0_wb_data_i[2]
  PIN master0_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END master0_wb_data_i[30]
  PIN master0_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END master0_wb_data_i[31]
  PIN master0_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END master0_wb_data_i[3]
  PIN master0_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END master0_wb_data_i[4]
  PIN master0_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END master0_wb_data_i[5]
  PIN master0_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END master0_wb_data_i[6]
  PIN master0_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END master0_wb_data_i[7]
  PIN master0_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END master0_wb_data_i[8]
  PIN master0_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END master0_wb_data_i[9]
  PIN master0_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END master0_wb_data_o[0]
  PIN master0_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END master0_wb_data_o[10]
  PIN master0_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END master0_wb_data_o[11]
  PIN master0_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END master0_wb_data_o[12]
  PIN master0_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END master0_wb_data_o[13]
  PIN master0_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END master0_wb_data_o[14]
  PIN master0_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END master0_wb_data_o[15]
  PIN master0_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END master0_wb_data_o[16]
  PIN master0_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END master0_wb_data_o[17]
  PIN master0_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END master0_wb_data_o[18]
  PIN master0_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END master0_wb_data_o[19]
  PIN master0_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END master0_wb_data_o[1]
  PIN master0_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END master0_wb_data_o[20]
  PIN master0_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END master0_wb_data_o[21]
  PIN master0_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END master0_wb_data_o[22]
  PIN master0_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END master0_wb_data_o[23]
  PIN master0_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END master0_wb_data_o[24]
  PIN master0_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END master0_wb_data_o[25]
  PIN master0_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END master0_wb_data_o[26]
  PIN master0_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END master0_wb_data_o[27]
  PIN master0_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END master0_wb_data_o[28]
  PIN master0_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END master0_wb_data_o[29]
  PIN master0_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END master0_wb_data_o[2]
  PIN master0_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END master0_wb_data_o[30]
  PIN master0_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END master0_wb_data_o[31]
  PIN master0_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END master0_wb_data_o[3]
  PIN master0_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END master0_wb_data_o[4]
  PIN master0_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END master0_wb_data_o[5]
  PIN master0_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END master0_wb_data_o[6]
  PIN master0_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END master0_wb_data_o[7]
  PIN master0_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END master0_wb_data_o[8]
  PIN master0_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END master0_wb_data_o[9]
  PIN master0_wb_error_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END master0_wb_error_i
  PIN master0_wb_sel_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END master0_wb_sel_o[0]
  PIN master0_wb_sel_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END master0_wb_sel_o[1]
  PIN master0_wb_sel_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END master0_wb_sel_o[2]
  PIN master0_wb_sel_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END master0_wb_sel_o[3]
  PIN master0_wb_stall_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END master0_wb_stall_i
  PIN master0_wb_stb_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END master0_wb_stb_o
  PIN master0_wb_we_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END master0_wb_we_o
  PIN master1_wb_ack_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END master1_wb_ack_i
  PIN master1_wb_adr_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END master1_wb_adr_o[0]
  PIN master1_wb_adr_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END master1_wb_adr_o[10]
  PIN master1_wb_adr_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END master1_wb_adr_o[11]
  PIN master1_wb_adr_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END master1_wb_adr_o[12]
  PIN master1_wb_adr_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END master1_wb_adr_o[13]
  PIN master1_wb_adr_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.280 4.000 692.880 ;
    END
  END master1_wb_adr_o[14]
  PIN master1_wb_adr_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END master1_wb_adr_o[15]
  PIN master1_wb_adr_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END master1_wb_adr_o[16]
  PIN master1_wb_adr_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END master1_wb_adr_o[17]
  PIN master1_wb_adr_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END master1_wb_adr_o[18]
  PIN master1_wb_adr_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END master1_wb_adr_o[19]
  PIN master1_wb_adr_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END master1_wb_adr_o[1]
  PIN master1_wb_adr_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END master1_wb_adr_o[20]
  PIN master1_wb_adr_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END master1_wb_adr_o[21]
  PIN master1_wb_adr_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END master1_wb_adr_o[22]
  PIN master1_wb_adr_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END master1_wb_adr_o[23]
  PIN master1_wb_adr_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.880 4.000 774.480 ;
    END
  END master1_wb_adr_o[24]
  PIN master1_wb_adr_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END master1_wb_adr_o[25]
  PIN master1_wb_adr_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.200 4.000 790.800 ;
    END
  END master1_wb_adr_o[26]
  PIN master1_wb_adr_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 798.360 4.000 798.960 ;
    END
  END master1_wb_adr_o[27]
  PIN master1_wb_adr_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END master1_wb_adr_o[2]
  PIN master1_wb_adr_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END master1_wb_adr_o[3]
  PIN master1_wb_adr_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END master1_wb_adr_o[4]
  PIN master1_wb_adr_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END master1_wb_adr_o[5]
  PIN master1_wb_adr_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END master1_wb_adr_o[6]
  PIN master1_wb_adr_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END master1_wb_adr_o[7]
  PIN master1_wb_adr_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END master1_wb_adr_o[8]
  PIN master1_wb_adr_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 651.480 4.000 652.080 ;
    END
  END master1_wb_adr_o[9]
  PIN master1_wb_cyc_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END master1_wb_cyc_o
  PIN master1_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END master1_wb_data_i[0]
  PIN master1_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END master1_wb_data_i[10]
  PIN master1_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END master1_wb_data_i[11]
  PIN master1_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END master1_wb_data_i[12]
  PIN master1_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END master1_wb_data_i[13]
  PIN master1_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END master1_wb_data_i[14]
  PIN master1_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END master1_wb_data_i[15]
  PIN master1_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END master1_wb_data_i[16]
  PIN master1_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END master1_wb_data_i[17]
  PIN master1_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END master1_wb_data_i[18]
  PIN master1_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END master1_wb_data_i[19]
  PIN master1_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END master1_wb_data_i[1]
  PIN master1_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END master1_wb_data_i[20]
  PIN master1_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END master1_wb_data_i[21]
  PIN master1_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END master1_wb_data_i[22]
  PIN master1_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END master1_wb_data_i[23]
  PIN master1_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END master1_wb_data_i[24]
  PIN master1_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END master1_wb_data_i[25]
  PIN master1_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END master1_wb_data_i[26]
  PIN master1_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 4.000 801.680 ;
    END
  END master1_wb_data_i[27]
  PIN master1_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 806.520 4.000 807.120 ;
    END
  END master1_wb_data_i[28]
  PIN master1_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.960 4.000 812.560 ;
    END
  END master1_wb_data_i[29]
  PIN master1_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END master1_wb_data_i[2]
  PIN master1_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END master1_wb_data_i[30]
  PIN master1_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END master1_wb_data_i[31]
  PIN master1_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END master1_wb_data_i[3]
  PIN master1_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END master1_wb_data_i[4]
  PIN master1_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END master1_wb_data_i[5]
  PIN master1_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END master1_wb_data_i[6]
  PIN master1_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END master1_wb_data_i[7]
  PIN master1_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END master1_wb_data_i[8]
  PIN master1_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END master1_wb_data_i[9]
  PIN master1_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END master1_wb_data_o[0]
  PIN master1_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END master1_wb_data_o[10]
  PIN master1_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END master1_wb_data_o[11]
  PIN master1_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END master1_wb_data_o[12]
  PIN master1_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END master1_wb_data_o[13]
  PIN master1_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END master1_wb_data_o[14]
  PIN master1_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END master1_wb_data_o[15]
  PIN master1_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END master1_wb_data_o[16]
  PIN master1_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END master1_wb_data_o[17]
  PIN master1_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END master1_wb_data_o[18]
  PIN master1_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END master1_wb_data_o[19]
  PIN master1_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END master1_wb_data_o[1]
  PIN master1_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END master1_wb_data_o[20]
  PIN master1_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END master1_wb_data_o[21]
  PIN master1_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END master1_wb_data_o[22]
  PIN master1_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.160 4.000 771.760 ;
    END
  END master1_wb_data_o[23]
  PIN master1_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END master1_wb_data_o[24]
  PIN master1_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END master1_wb_data_o[25]
  PIN master1_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END master1_wb_data_o[26]
  PIN master1_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.800 4.000 804.400 ;
    END
  END master1_wb_data_o[27]
  PIN master1_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END master1_wb_data_o[28]
  PIN master1_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END master1_wb_data_o[29]
  PIN master1_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END master1_wb_data_o[2]
  PIN master1_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 4.000 820.720 ;
    END
  END master1_wb_data_o[30]
  PIN master1_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END master1_wb_data_o[31]
  PIN master1_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END master1_wb_data_o[3]
  PIN master1_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END master1_wb_data_o[4]
  PIN master1_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END master1_wb_data_o[5]
  PIN master1_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END master1_wb_data_o[6]
  PIN master1_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END master1_wb_data_o[7]
  PIN master1_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END master1_wb_data_o[8]
  PIN master1_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 4.000 657.520 ;
    END
  END master1_wb_data_o[9]
  PIN master1_wb_error_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END master1_wb_error_i
  PIN master1_wb_sel_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END master1_wb_sel_o[0]
  PIN master1_wb_sel_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END master1_wb_sel_o[1]
  PIN master1_wb_sel_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END master1_wb_sel_o[2]
  PIN master1_wb_sel_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END master1_wb_sel_o[3]
  PIN master1_wb_stall_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END master1_wb_stall_i
  PIN master1_wb_stb_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END master1_wb_stb_o
  PIN master1_wb_we_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END master1_wb_we_o
  PIN master2_wb_ack_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END master2_wb_ack_i
  PIN master2_wb_adr_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END master2_wb_adr_o[0]
  PIN master2_wb_adr_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END master2_wb_adr_o[10]
  PIN master2_wb_adr_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END master2_wb_adr_o[11]
  PIN master2_wb_adr_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END master2_wb_adr_o[12]
  PIN master2_wb_adr_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END master2_wb_adr_o[13]
  PIN master2_wb_adr_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END master2_wb_adr_o[14]
  PIN master2_wb_adr_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END master2_wb_adr_o[15]
  PIN master2_wb_adr_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END master2_wb_adr_o[16]
  PIN master2_wb_adr_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END master2_wb_adr_o[17]
  PIN master2_wb_adr_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END master2_wb_adr_o[18]
  PIN master2_wb_adr_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END master2_wb_adr_o[19]
  PIN master2_wb_adr_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END master2_wb_adr_o[1]
  PIN master2_wb_adr_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END master2_wb_adr_o[20]
  PIN master2_wb_adr_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END master2_wb_adr_o[21]
  PIN master2_wb_adr_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END master2_wb_adr_o[22]
  PIN master2_wb_adr_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END master2_wb_adr_o[23]
  PIN master2_wb_adr_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END master2_wb_adr_o[24]
  PIN master2_wb_adr_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END master2_wb_adr_o[25]
  PIN master2_wb_adr_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END master2_wb_adr_o[26]
  PIN master2_wb_adr_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END master2_wb_adr_o[27]
  PIN master2_wb_adr_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END master2_wb_adr_o[2]
  PIN master2_wb_adr_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END master2_wb_adr_o[3]
  PIN master2_wb_adr_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END master2_wb_adr_o[4]
  PIN master2_wb_adr_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END master2_wb_adr_o[5]
  PIN master2_wb_adr_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END master2_wb_adr_o[6]
  PIN master2_wb_adr_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END master2_wb_adr_o[7]
  PIN master2_wb_adr_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END master2_wb_adr_o[8]
  PIN master2_wb_adr_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END master2_wb_adr_o[9]
  PIN master2_wb_cyc_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END master2_wb_cyc_o
  PIN master2_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END master2_wb_data_i[0]
  PIN master2_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END master2_wb_data_i[10]
  PIN master2_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END master2_wb_data_i[11]
  PIN master2_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END master2_wb_data_i[12]
  PIN master2_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END master2_wb_data_i[13]
  PIN master2_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END master2_wb_data_i[14]
  PIN master2_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END master2_wb_data_i[15]
  PIN master2_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END master2_wb_data_i[16]
  PIN master2_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END master2_wb_data_i[17]
  PIN master2_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END master2_wb_data_i[18]
  PIN master2_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END master2_wb_data_i[19]
  PIN master2_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END master2_wb_data_i[1]
  PIN master2_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END master2_wb_data_i[20]
  PIN master2_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END master2_wb_data_i[21]
  PIN master2_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END master2_wb_data_i[22]
  PIN master2_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END master2_wb_data_i[23]
  PIN master2_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END master2_wb_data_i[24]
  PIN master2_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END master2_wb_data_i[25]
  PIN master2_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END master2_wb_data_i[26]
  PIN master2_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END master2_wb_data_i[27]
  PIN master2_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END master2_wb_data_i[28]
  PIN master2_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END master2_wb_data_i[29]
  PIN master2_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END master2_wb_data_i[2]
  PIN master2_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END master2_wb_data_i[30]
  PIN master2_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END master2_wb_data_i[31]
  PIN master2_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END master2_wb_data_i[3]
  PIN master2_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END master2_wb_data_i[4]
  PIN master2_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END master2_wb_data_i[5]
  PIN master2_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END master2_wb_data_i[6]
  PIN master2_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END master2_wb_data_i[7]
  PIN master2_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END master2_wb_data_i[8]
  PIN master2_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END master2_wb_data_i[9]
  PIN master2_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END master2_wb_data_o[0]
  PIN master2_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END master2_wb_data_o[10]
  PIN master2_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END master2_wb_data_o[11]
  PIN master2_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END master2_wb_data_o[12]
  PIN master2_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END master2_wb_data_o[13]
  PIN master2_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END master2_wb_data_o[14]
  PIN master2_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END master2_wb_data_o[15]
  PIN master2_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END master2_wb_data_o[16]
  PIN master2_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END master2_wb_data_o[17]
  PIN master2_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END master2_wb_data_o[18]
  PIN master2_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END master2_wb_data_o[19]
  PIN master2_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END master2_wb_data_o[1]
  PIN master2_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END master2_wb_data_o[20]
  PIN master2_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END master2_wb_data_o[21]
  PIN master2_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END master2_wb_data_o[22]
  PIN master2_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END master2_wb_data_o[23]
  PIN master2_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END master2_wb_data_o[24]
  PIN master2_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END master2_wb_data_o[25]
  PIN master2_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END master2_wb_data_o[26]
  PIN master2_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END master2_wb_data_o[27]
  PIN master2_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END master2_wb_data_o[28]
  PIN master2_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END master2_wb_data_o[29]
  PIN master2_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END master2_wb_data_o[2]
  PIN master2_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END master2_wb_data_o[30]
  PIN master2_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END master2_wb_data_o[31]
  PIN master2_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END master2_wb_data_o[3]
  PIN master2_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END master2_wb_data_o[4]
  PIN master2_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END master2_wb_data_o[5]
  PIN master2_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END master2_wb_data_o[6]
  PIN master2_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END master2_wb_data_o[7]
  PIN master2_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END master2_wb_data_o[8]
  PIN master2_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END master2_wb_data_o[9]
  PIN master2_wb_error_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END master2_wb_error_i
  PIN master2_wb_sel_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END master2_wb_sel_o[0]
  PIN master2_wb_sel_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END master2_wb_sel_o[1]
  PIN master2_wb_sel_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END master2_wb_sel_o[2]
  PIN master2_wb_sel_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END master2_wb_sel_o[3]
  PIN master2_wb_stall_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END master2_wb_stall_i
  PIN master2_wb_stb_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END master2_wb_stb_o
  PIN master2_wb_we_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END master2_wb_we_o
  PIN probe_master0_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END probe_master0_currentSlave[0]
  PIN probe_master0_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END probe_master0_currentSlave[1]
  PIN probe_master1_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END probe_master1_currentSlave[0]
  PIN probe_master1_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END probe_master1_currentSlave[1]
  PIN probe_master2_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END probe_master2_currentSlave[0]
  PIN probe_master2_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END probe_master2_currentSlave[1]
  PIN probe_master3_currentSlave[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END probe_master3_currentSlave[0]
  PIN probe_master3_currentSlave[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END probe_master3_currentSlave[1]
  PIN probe_slave0_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END probe_slave0_currentMaster[0]
  PIN probe_slave0_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END probe_slave0_currentMaster[1]
  PIN probe_slave1_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END probe_slave1_currentMaster[0]
  PIN probe_slave1_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END probe_slave1_currentMaster[1]
  PIN probe_slave2_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END probe_slave2_currentMaster[0]
  PIN probe_slave2_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END probe_slave2_currentMaster[1]
  PIN probe_slave3_currentMaster[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END probe_slave3_currentMaster[0]
  PIN probe_slave3_currentMaster[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END probe_slave3_currentMaster[1]
  PIN slave0_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END slave0_wb_ack_o
  PIN slave0_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 844.600 4.000 845.200 ;
    END
  END slave0_wb_adr_i[0]
  PIN slave0_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.080 4.000 937.680 ;
    END
  END slave0_wb_adr_i[10]
  PIN slave0_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END slave0_wb_adr_i[11]
  PIN slave0_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 953.400 4.000 954.000 ;
    END
  END slave0_wb_adr_i[12]
  PIN slave0_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 961.560 4.000 962.160 ;
    END
  END slave0_wb_adr_i[13]
  PIN slave0_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.720 4.000 970.320 ;
    END
  END slave0_wb_adr_i[14]
  PIN slave0_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.880 4.000 978.480 ;
    END
  END slave0_wb_adr_i[15]
  PIN slave0_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END slave0_wb_adr_i[16]
  PIN slave0_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END slave0_wb_adr_i[17]
  PIN slave0_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1002.360 4.000 1002.960 ;
    END
  END slave0_wb_adr_i[18]
  PIN slave0_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1010.520 4.000 1011.120 ;
    END
  END slave0_wb_adr_i[19]
  PIN slave0_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 855.480 4.000 856.080 ;
    END
  END slave0_wb_adr_i[1]
  PIN slave0_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.680 4.000 1019.280 ;
    END
  END slave0_wb_adr_i[20]
  PIN slave0_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END slave0_wb_adr_i[21]
  PIN slave0_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1035.000 4.000 1035.600 ;
    END
  END slave0_wb_adr_i[22]
  PIN slave0_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.160 4.000 1043.760 ;
    END
  END slave0_wb_adr_i[23]
  PIN slave0_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END slave0_wb_adr_i[2]
  PIN slave0_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END slave0_wb_adr_i[3]
  PIN slave0_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END slave0_wb_adr_i[4]
  PIN slave0_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.280 4.000 896.880 ;
    END
  END slave0_wb_adr_i[5]
  PIN slave0_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END slave0_wb_adr_i[6]
  PIN slave0_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 912.600 4.000 913.200 ;
    END
  END slave0_wb_adr_i[7]
  PIN slave0_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.760 4.000 921.360 ;
    END
  END slave0_wb_adr_i[8]
  PIN slave0_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.920 4.000 929.520 ;
    END
  END slave0_wb_adr_i[9]
  PIN slave0_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.000 4.000 831.600 ;
    END
  END slave0_wb_cyc_i
  PIN slave0_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 847.320 4.000 847.920 ;
    END
  END slave0_wb_data_i[0]
  PIN slave0_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.800 4.000 940.400 ;
    END
  END slave0_wb_data_i[10]
  PIN slave0_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.960 4.000 948.560 ;
    END
  END slave0_wb_data_i[11]
  PIN slave0_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 956.120 4.000 956.720 ;
    END
  END slave0_wb_data_i[12]
  PIN slave0_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.280 4.000 964.880 ;
    END
  END slave0_wb_data_i[13]
  PIN slave0_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END slave0_wb_data_i[14]
  PIN slave0_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END slave0_wb_data_i[15]
  PIN slave0_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 988.760 4.000 989.360 ;
    END
  END slave0_wb_data_i[16]
  PIN slave0_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.920 4.000 997.520 ;
    END
  END slave0_wb_data_i[17]
  PIN slave0_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.080 4.000 1005.680 ;
    END
  END slave0_wb_data_i[18]
  PIN slave0_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END slave0_wb_data_i[19]
  PIN slave0_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.200 4.000 858.800 ;
    END
  END slave0_wb_data_i[1]
  PIN slave0_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1021.400 4.000 1022.000 ;
    END
  END slave0_wb_data_i[20]
  PIN slave0_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END slave0_wb_data_i[21]
  PIN slave0_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.720 4.000 1038.320 ;
    END
  END slave0_wb_data_i[22]
  PIN slave0_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.880 4.000 1046.480 ;
    END
  END slave0_wb_data_i[23]
  PIN slave0_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1051.320 4.000 1051.920 ;
    END
  END slave0_wb_data_i[24]
  PIN slave0_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.760 4.000 1057.360 ;
    END
  END slave0_wb_data_i[25]
  PIN slave0_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.200 4.000 1062.800 ;
    END
  END slave0_wb_data_i[26]
  PIN slave0_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END slave0_wb_data_i[27]
  PIN slave0_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1073.080 4.000 1073.680 ;
    END
  END slave0_wb_data_i[28]
  PIN slave0_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1078.520 4.000 1079.120 ;
    END
  END slave0_wb_data_i[29]
  PIN slave0_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 869.080 4.000 869.680 ;
    END
  END slave0_wb_data_i[2]
  PIN slave0_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1083.960 4.000 1084.560 ;
    END
  END slave0_wb_data_i[30]
  PIN slave0_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1089.400 4.000 1090.000 ;
    END
  END slave0_wb_data_i[31]
  PIN slave0_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.960 4.000 880.560 ;
    END
  END slave0_wb_data_i[3]
  PIN slave0_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END slave0_wb_data_i[4]
  PIN slave0_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END slave0_wb_data_i[5]
  PIN slave0_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.160 4.000 907.760 ;
    END
  END slave0_wb_data_i[6]
  PIN slave0_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 915.320 4.000 915.920 ;
    END
  END slave0_wb_data_i[7]
  PIN slave0_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 923.480 4.000 924.080 ;
    END
  END slave0_wb_data_i[8]
  PIN slave0_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END slave0_wb_data_i[9]
  PIN slave0_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END slave0_wb_data_o[0]
  PIN slave0_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 942.520 4.000 943.120 ;
    END
  END slave0_wb_data_o[10]
  PIN slave0_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.680 4.000 951.280 ;
    END
  END slave0_wb_data_o[11]
  PIN slave0_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END slave0_wb_data_o[12]
  PIN slave0_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 967.000 4.000 967.600 ;
    END
  END slave0_wb_data_o[13]
  PIN slave0_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.160 4.000 975.760 ;
    END
  END slave0_wb_data_o[14]
  PIN slave0_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END slave0_wb_data_o[15]
  PIN slave0_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 991.480 4.000 992.080 ;
    END
  END slave0_wb_data_o[16]
  PIN slave0_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END slave0_wb_data_o[17]
  PIN slave0_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 4.000 1008.400 ;
    END
  END slave0_wb_data_o[18]
  PIN slave0_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1015.960 4.000 1016.560 ;
    END
  END slave0_wb_data_o[19]
  PIN slave0_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.920 4.000 861.520 ;
    END
  END slave0_wb_data_o[1]
  PIN slave0_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.120 4.000 1024.720 ;
    END
  END slave0_wb_data_o[20]
  PIN slave0_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.280 4.000 1032.880 ;
    END
  END slave0_wb_data_o[21]
  PIN slave0_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END slave0_wb_data_o[22]
  PIN slave0_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1048.600 4.000 1049.200 ;
    END
  END slave0_wb_data_o[23]
  PIN slave0_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END slave0_wb_data_o[24]
  PIN slave0_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1059.480 4.000 1060.080 ;
    END
  END slave0_wb_data_o[25]
  PIN slave0_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.920 4.000 1065.520 ;
    END
  END slave0_wb_data_o[26]
  PIN slave0_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1070.360 4.000 1070.960 ;
    END
  END slave0_wb_data_o[27]
  PIN slave0_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.800 4.000 1076.400 ;
    END
  END slave0_wb_data_o[28]
  PIN slave0_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END slave0_wb_data_o[29]
  PIN slave0_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.800 4.000 872.400 ;
    END
  END slave0_wb_data_o[2]
  PIN slave0_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1086.680 4.000 1087.280 ;
    END
  END slave0_wb_data_o[30]
  PIN slave0_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1092.120 4.000 1092.720 ;
    END
  END slave0_wb_data_o[31]
  PIN slave0_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 882.680 4.000 883.280 ;
    END
  END slave0_wb_data_o[3]
  PIN slave0_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END slave0_wb_data_o[4]
  PIN slave0_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.720 4.000 902.320 ;
    END
  END slave0_wb_data_o[5]
  PIN slave0_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END slave0_wb_data_o[6]
  PIN slave0_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END slave0_wb_data_o[7]
  PIN slave0_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.200 4.000 926.800 ;
    END
  END slave0_wb_data_o[8]
  PIN slave0_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 934.360 4.000 934.960 ;
    END
  END slave0_wb_data_o[9]
  PIN slave0_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.720 4.000 834.320 ;
    END
  END slave0_wb_error_o
  PIN slave0_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.760 4.000 853.360 ;
    END
  END slave0_wb_sel_i[0]
  PIN slave0_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END slave0_wb_sel_i[1]
  PIN slave0_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 874.520 4.000 875.120 ;
    END
  END slave0_wb_sel_i[2]
  PIN slave0_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 885.400 4.000 886.000 ;
    END
  END slave0_wb_sel_i[3]
  PIN slave0_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END slave0_wb_stall_o
  PIN slave0_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END slave0_wb_stb_i
  PIN slave0_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 841.880 4.000 842.480 ;
    END
  END slave0_wb_we_i
  PIN slave1_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END slave1_wb_ack_o
  PIN slave1_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END slave1_wb_adr_i[0]
  PIN slave1_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END slave1_wb_adr_i[10]
  PIN slave1_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END slave1_wb_adr_i[11]
  PIN slave1_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END slave1_wb_adr_i[12]
  PIN slave1_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END slave1_wb_adr_i[13]
  PIN slave1_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END slave1_wb_adr_i[14]
  PIN slave1_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END slave1_wb_adr_i[15]
  PIN slave1_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END slave1_wb_adr_i[16]
  PIN slave1_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END slave1_wb_adr_i[17]
  PIN slave1_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END slave1_wb_adr_i[18]
  PIN slave1_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END slave1_wb_adr_i[19]
  PIN slave1_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END slave1_wb_adr_i[1]
  PIN slave1_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END slave1_wb_adr_i[20]
  PIN slave1_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END slave1_wb_adr_i[21]
  PIN slave1_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END slave1_wb_adr_i[22]
  PIN slave1_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END slave1_wb_adr_i[23]
  PIN slave1_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END slave1_wb_adr_i[2]
  PIN slave1_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END slave1_wb_adr_i[3]
  PIN slave1_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END slave1_wb_adr_i[4]
  PIN slave1_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END slave1_wb_adr_i[5]
  PIN slave1_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END slave1_wb_adr_i[6]
  PIN slave1_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END slave1_wb_adr_i[7]
  PIN slave1_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END slave1_wb_adr_i[8]
  PIN slave1_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END slave1_wb_adr_i[9]
  PIN slave1_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END slave1_wb_cyc_i
  PIN slave1_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END slave1_wb_data_i[0]
  PIN slave1_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END slave1_wb_data_i[10]
  PIN slave1_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END slave1_wb_data_i[11]
  PIN slave1_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END slave1_wb_data_i[12]
  PIN slave1_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END slave1_wb_data_i[13]
  PIN slave1_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END slave1_wb_data_i[14]
  PIN slave1_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END slave1_wb_data_i[15]
  PIN slave1_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END slave1_wb_data_i[16]
  PIN slave1_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END slave1_wb_data_i[17]
  PIN slave1_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END slave1_wb_data_i[18]
  PIN slave1_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END slave1_wb_data_i[19]
  PIN slave1_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END slave1_wb_data_i[1]
  PIN slave1_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END slave1_wb_data_i[20]
  PIN slave1_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END slave1_wb_data_i[21]
  PIN slave1_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END slave1_wb_data_i[22]
  PIN slave1_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END slave1_wb_data_i[23]
  PIN slave1_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END slave1_wb_data_i[24]
  PIN slave1_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END slave1_wb_data_i[25]
  PIN slave1_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END slave1_wb_data_i[26]
  PIN slave1_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END slave1_wb_data_i[27]
  PIN slave1_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END slave1_wb_data_i[28]
  PIN slave1_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END slave1_wb_data_i[29]
  PIN slave1_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END slave1_wb_data_i[2]
  PIN slave1_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END slave1_wb_data_i[30]
  PIN slave1_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END slave1_wb_data_i[31]
  PIN slave1_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END slave1_wb_data_i[3]
  PIN slave1_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END slave1_wb_data_i[4]
  PIN slave1_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END slave1_wb_data_i[5]
  PIN slave1_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END slave1_wb_data_i[6]
  PIN slave1_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END slave1_wb_data_i[7]
  PIN slave1_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END slave1_wb_data_i[8]
  PIN slave1_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END slave1_wb_data_i[9]
  PIN slave1_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END slave1_wb_data_o[0]
  PIN slave1_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END slave1_wb_data_o[10]
  PIN slave1_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END slave1_wb_data_o[11]
  PIN slave1_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END slave1_wb_data_o[12]
  PIN slave1_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END slave1_wb_data_o[13]
  PIN slave1_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END slave1_wb_data_o[14]
  PIN slave1_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END slave1_wb_data_o[15]
  PIN slave1_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END slave1_wb_data_o[16]
  PIN slave1_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END slave1_wb_data_o[17]
  PIN slave1_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END slave1_wb_data_o[18]
  PIN slave1_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END slave1_wb_data_o[19]
  PIN slave1_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END slave1_wb_data_o[1]
  PIN slave1_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END slave1_wb_data_o[20]
  PIN slave1_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END slave1_wb_data_o[21]
  PIN slave1_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END slave1_wb_data_o[22]
  PIN slave1_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END slave1_wb_data_o[23]
  PIN slave1_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END slave1_wb_data_o[24]
  PIN slave1_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END slave1_wb_data_o[25]
  PIN slave1_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END slave1_wb_data_o[26]
  PIN slave1_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END slave1_wb_data_o[27]
  PIN slave1_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END slave1_wb_data_o[28]
  PIN slave1_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END slave1_wb_data_o[29]
  PIN slave1_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END slave1_wb_data_o[2]
  PIN slave1_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END slave1_wb_data_o[30]
  PIN slave1_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END slave1_wb_data_o[31]
  PIN slave1_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END slave1_wb_data_o[3]
  PIN slave1_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END slave1_wb_data_o[4]
  PIN slave1_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END slave1_wb_data_o[5]
  PIN slave1_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END slave1_wb_data_o[6]
  PIN slave1_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END slave1_wb_data_o[7]
  PIN slave1_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END slave1_wb_data_o[8]
  PIN slave1_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END slave1_wb_data_o[9]
  PIN slave1_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END slave1_wb_error_o
  PIN slave1_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END slave1_wb_sel_i[0]
  PIN slave1_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END slave1_wb_sel_i[1]
  PIN slave1_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END slave1_wb_sel_i[2]
  PIN slave1_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END slave1_wb_sel_i[3]
  PIN slave1_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END slave1_wb_stall_o
  PIN slave1_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END slave1_wb_stb_i
  PIN slave1_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END slave1_wb_we_i
  PIN slave2_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 1096.000 18.770 1100.000 ;
    END
  END slave2_wb_ack_o
  PIN slave2_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 1096.000 38.090 1100.000 ;
    END
  END slave2_wb_adr_i[0]
  PIN slave2_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 1096.000 147.570 1100.000 ;
    END
  END slave2_wb_adr_i[10]
  PIN slave2_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 1096.000 157.230 1100.000 ;
    END
  END slave2_wb_adr_i[11]
  PIN slave2_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 1096.000 166.890 1100.000 ;
    END
  END slave2_wb_adr_i[12]
  PIN slave2_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 1096.000 176.550 1100.000 ;
    END
  END slave2_wb_adr_i[13]
  PIN slave2_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 1096.000 186.210 1100.000 ;
    END
  END slave2_wb_adr_i[14]
  PIN slave2_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 1096.000 195.870 1100.000 ;
    END
  END slave2_wb_adr_i[15]
  PIN slave2_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 1096.000 205.530 1100.000 ;
    END
  END slave2_wb_adr_i[16]
  PIN slave2_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 1096.000 215.190 1100.000 ;
    END
  END slave2_wb_adr_i[17]
  PIN slave2_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 1096.000 224.850 1100.000 ;
    END
  END slave2_wb_adr_i[18]
  PIN slave2_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 1096.000 234.510 1100.000 ;
    END
  END slave2_wb_adr_i[19]
  PIN slave2_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 1096.000 50.970 1100.000 ;
    END
  END slave2_wb_adr_i[1]
  PIN slave2_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 1096.000 244.170 1100.000 ;
    END
  END slave2_wb_adr_i[20]
  PIN slave2_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 1096.000 253.830 1100.000 ;
    END
  END slave2_wb_adr_i[21]
  PIN slave2_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 1096.000 263.490 1100.000 ;
    END
  END slave2_wb_adr_i[22]
  PIN slave2_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 1096.000 273.150 1100.000 ;
    END
  END slave2_wb_adr_i[23]
  PIN slave2_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 1096.000 63.850 1100.000 ;
    END
  END slave2_wb_adr_i[2]
  PIN slave2_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 1096.000 76.730 1100.000 ;
    END
  END slave2_wb_adr_i[3]
  PIN slave2_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 1096.000 89.610 1100.000 ;
    END
  END slave2_wb_adr_i[4]
  PIN slave2_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 1096.000 99.270 1100.000 ;
    END
  END slave2_wb_adr_i[5]
  PIN slave2_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 1096.000 108.930 1100.000 ;
    END
  END slave2_wb_adr_i[6]
  PIN slave2_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 1096.000 118.590 1100.000 ;
    END
  END slave2_wb_adr_i[7]
  PIN slave2_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 1096.000 128.250 1100.000 ;
    END
  END slave2_wb_adr_i[8]
  PIN slave2_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 1096.000 137.910 1100.000 ;
    END
  END slave2_wb_adr_i[9]
  PIN slave2_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 1096.000 21.990 1100.000 ;
    END
  END slave2_wb_cyc_i
  PIN slave2_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 1096.000 41.310 1100.000 ;
    END
  END slave2_wb_data_i[0]
  PIN slave2_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 1096.000 150.790 1100.000 ;
    END
  END slave2_wb_data_i[10]
  PIN slave2_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 1096.000 160.450 1100.000 ;
    END
  END slave2_wb_data_i[11]
  PIN slave2_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 1096.000 170.110 1100.000 ;
    END
  END slave2_wb_data_i[12]
  PIN slave2_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 1096.000 179.770 1100.000 ;
    END
  END slave2_wb_data_i[13]
  PIN slave2_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 1096.000 189.430 1100.000 ;
    END
  END slave2_wb_data_i[14]
  PIN slave2_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 1096.000 199.090 1100.000 ;
    END
  END slave2_wb_data_i[15]
  PIN slave2_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 1096.000 208.750 1100.000 ;
    END
  END slave2_wb_data_i[16]
  PIN slave2_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 1096.000 218.410 1100.000 ;
    END
  END slave2_wb_data_i[17]
  PIN slave2_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 1096.000 228.070 1100.000 ;
    END
  END slave2_wb_data_i[18]
  PIN slave2_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 1096.000 237.730 1100.000 ;
    END
  END slave2_wb_data_i[19]
  PIN slave2_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 1096.000 54.190 1100.000 ;
    END
  END slave2_wb_data_i[1]
  PIN slave2_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 1096.000 247.390 1100.000 ;
    END
  END slave2_wb_data_i[20]
  PIN slave2_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 1096.000 257.050 1100.000 ;
    END
  END slave2_wb_data_i[21]
  PIN slave2_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 1096.000 266.710 1100.000 ;
    END
  END slave2_wb_data_i[22]
  PIN slave2_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 1096.000 276.370 1100.000 ;
    END
  END slave2_wb_data_i[23]
  PIN slave2_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 1096.000 282.810 1100.000 ;
    END
  END slave2_wb_data_i[24]
  PIN slave2_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 1096.000 289.250 1100.000 ;
    END
  END slave2_wb_data_i[25]
  PIN slave2_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 1096.000 295.690 1100.000 ;
    END
  END slave2_wb_data_i[26]
  PIN slave2_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 1096.000 302.130 1100.000 ;
    END
  END slave2_wb_data_i[27]
  PIN slave2_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 1096.000 308.570 1100.000 ;
    END
  END slave2_wb_data_i[28]
  PIN slave2_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 1096.000 315.010 1100.000 ;
    END
  END slave2_wb_data_i[29]
  PIN slave2_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 1096.000 67.070 1100.000 ;
    END
  END slave2_wb_data_i[2]
  PIN slave2_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 1096.000 321.450 1100.000 ;
    END
  END slave2_wb_data_i[30]
  PIN slave2_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 1096.000 327.890 1100.000 ;
    END
  END slave2_wb_data_i[31]
  PIN slave2_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 1096.000 79.950 1100.000 ;
    END
  END slave2_wb_data_i[3]
  PIN slave2_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 1096.000 92.830 1100.000 ;
    END
  END slave2_wb_data_i[4]
  PIN slave2_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 1096.000 102.490 1100.000 ;
    END
  END slave2_wb_data_i[5]
  PIN slave2_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 1096.000 112.150 1100.000 ;
    END
  END slave2_wb_data_i[6]
  PIN slave2_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 1096.000 121.810 1100.000 ;
    END
  END slave2_wb_data_i[7]
  PIN slave2_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 1096.000 131.470 1100.000 ;
    END
  END slave2_wb_data_i[8]
  PIN slave2_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 1096.000 141.130 1100.000 ;
    END
  END slave2_wb_data_i[9]
  PIN slave2_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 1096.000 44.530 1100.000 ;
    END
  END slave2_wb_data_o[0]
  PIN slave2_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 1096.000 154.010 1100.000 ;
    END
  END slave2_wb_data_o[10]
  PIN slave2_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 1096.000 163.670 1100.000 ;
    END
  END slave2_wb_data_o[11]
  PIN slave2_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 1096.000 173.330 1100.000 ;
    END
  END slave2_wb_data_o[12]
  PIN slave2_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 1096.000 182.990 1100.000 ;
    END
  END slave2_wb_data_o[13]
  PIN slave2_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 1096.000 192.650 1100.000 ;
    END
  END slave2_wb_data_o[14]
  PIN slave2_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 1096.000 202.310 1100.000 ;
    END
  END slave2_wb_data_o[15]
  PIN slave2_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 1096.000 211.970 1100.000 ;
    END
  END slave2_wb_data_o[16]
  PIN slave2_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 1096.000 221.630 1100.000 ;
    END
  END slave2_wb_data_o[17]
  PIN slave2_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 1096.000 231.290 1100.000 ;
    END
  END slave2_wb_data_o[18]
  PIN slave2_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 1096.000 240.950 1100.000 ;
    END
  END slave2_wb_data_o[19]
  PIN slave2_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 1096.000 57.410 1100.000 ;
    END
  END slave2_wb_data_o[1]
  PIN slave2_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 1096.000 250.610 1100.000 ;
    END
  END slave2_wb_data_o[20]
  PIN slave2_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 1096.000 260.270 1100.000 ;
    END
  END slave2_wb_data_o[21]
  PIN slave2_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 1096.000 269.930 1100.000 ;
    END
  END slave2_wb_data_o[22]
  PIN slave2_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 1096.000 279.590 1100.000 ;
    END
  END slave2_wb_data_o[23]
  PIN slave2_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 1096.000 286.030 1100.000 ;
    END
  END slave2_wb_data_o[24]
  PIN slave2_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 1096.000 292.470 1100.000 ;
    END
  END slave2_wb_data_o[25]
  PIN slave2_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 1096.000 298.910 1100.000 ;
    END
  END slave2_wb_data_o[26]
  PIN slave2_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 1096.000 305.350 1100.000 ;
    END
  END slave2_wb_data_o[27]
  PIN slave2_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 1096.000 311.790 1100.000 ;
    END
  END slave2_wb_data_o[28]
  PIN slave2_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 1096.000 318.230 1100.000 ;
    END
  END slave2_wb_data_o[29]
  PIN slave2_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 1096.000 70.290 1100.000 ;
    END
  END slave2_wb_data_o[2]
  PIN slave2_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 1096.000 324.670 1100.000 ;
    END
  END slave2_wb_data_o[30]
  PIN slave2_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 1096.000 331.110 1100.000 ;
    END
  END slave2_wb_data_o[31]
  PIN slave2_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 1096.000 83.170 1100.000 ;
    END
  END slave2_wb_data_o[3]
  PIN slave2_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 1096.000 96.050 1100.000 ;
    END
  END slave2_wb_data_o[4]
  PIN slave2_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 1096.000 105.710 1100.000 ;
    END
  END slave2_wb_data_o[5]
  PIN slave2_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 1096.000 115.370 1100.000 ;
    END
  END slave2_wb_data_o[6]
  PIN slave2_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 1096.000 125.030 1100.000 ;
    END
  END slave2_wb_data_o[7]
  PIN slave2_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 1096.000 134.690 1100.000 ;
    END
  END slave2_wb_data_o[8]
  PIN slave2_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 1096.000 144.350 1100.000 ;
    END
  END slave2_wb_data_o[9]
  PIN slave2_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 1096.000 25.210 1100.000 ;
    END
  END slave2_wb_error_o
  PIN slave2_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 1096.000 47.750 1100.000 ;
    END
  END slave2_wb_sel_i[0]
  PIN slave2_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 1096.000 60.630 1100.000 ;
    END
  END slave2_wb_sel_i[1]
  PIN slave2_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 1096.000 73.510 1100.000 ;
    END
  END slave2_wb_sel_i[2]
  PIN slave2_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 1096.000 86.390 1100.000 ;
    END
  END slave2_wb_sel_i[3]
  PIN slave2_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 1096.000 28.430 1100.000 ;
    END
  END slave2_wb_stall_o
  PIN slave2_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 1096.000 31.650 1100.000 ;
    END
  END slave2_wb_stb_i
  PIN slave2_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 1096.000 34.870 1100.000 ;
    END
  END slave2_wb_we_i
  PIN slave3_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 552.200 350.000 552.800 ;
    END
  END slave3_wb_ack_o
  PIN slave3_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 584.840 350.000 585.440 ;
    END
  END slave3_wb_adr_i[0]
  PIN slave3_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 769.800 350.000 770.400 ;
    END
  END slave3_wb_adr_i[10]
  PIN slave3_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 786.120 350.000 786.720 ;
    END
  END slave3_wb_adr_i[11]
  PIN slave3_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 802.440 350.000 803.040 ;
    END
  END slave3_wb_adr_i[12]
  PIN slave3_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 818.760 350.000 819.360 ;
    END
  END slave3_wb_adr_i[13]
  PIN slave3_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 835.080 350.000 835.680 ;
    END
  END slave3_wb_adr_i[14]
  PIN slave3_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 851.400 350.000 852.000 ;
    END
  END slave3_wb_adr_i[15]
  PIN slave3_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 867.720 350.000 868.320 ;
    END
  END slave3_wb_adr_i[16]
  PIN slave3_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 884.040 350.000 884.640 ;
    END
  END slave3_wb_adr_i[17]
  PIN slave3_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 900.360 350.000 900.960 ;
    END
  END slave3_wb_adr_i[18]
  PIN slave3_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 916.680 350.000 917.280 ;
    END
  END slave3_wb_adr_i[19]
  PIN slave3_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 606.600 350.000 607.200 ;
    END
  END slave3_wb_adr_i[1]
  PIN slave3_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 933.000 350.000 933.600 ;
    END
  END slave3_wb_adr_i[20]
  PIN slave3_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 949.320 350.000 949.920 ;
    END
  END slave3_wb_adr_i[21]
  PIN slave3_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 965.640 350.000 966.240 ;
    END
  END slave3_wb_adr_i[22]
  PIN slave3_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 981.960 350.000 982.560 ;
    END
  END slave3_wb_adr_i[23]
  PIN slave3_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 628.360 350.000 628.960 ;
    END
  END slave3_wb_adr_i[2]
  PIN slave3_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 650.120 350.000 650.720 ;
    END
  END slave3_wb_adr_i[3]
  PIN slave3_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 671.880 350.000 672.480 ;
    END
  END slave3_wb_adr_i[4]
  PIN slave3_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 688.200 350.000 688.800 ;
    END
  END slave3_wb_adr_i[5]
  PIN slave3_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 704.520 350.000 705.120 ;
    END
  END slave3_wb_adr_i[6]
  PIN slave3_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 720.840 350.000 721.440 ;
    END
  END slave3_wb_adr_i[7]
  PIN slave3_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 737.160 350.000 737.760 ;
    END
  END slave3_wb_adr_i[8]
  PIN slave3_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 753.480 350.000 754.080 ;
    END
  END slave3_wb_adr_i[9]
  PIN slave3_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 557.640 350.000 558.240 ;
    END
  END slave3_wb_cyc_i
  PIN slave3_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 590.280 350.000 590.880 ;
    END
  END slave3_wb_data_i[0]
  PIN slave3_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 775.240 350.000 775.840 ;
    END
  END slave3_wb_data_i[10]
  PIN slave3_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 791.560 350.000 792.160 ;
    END
  END slave3_wb_data_i[11]
  PIN slave3_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 807.880 350.000 808.480 ;
    END
  END slave3_wb_data_i[12]
  PIN slave3_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 824.200 350.000 824.800 ;
    END
  END slave3_wb_data_i[13]
  PIN slave3_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 840.520 350.000 841.120 ;
    END
  END slave3_wb_data_i[14]
  PIN slave3_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 856.840 350.000 857.440 ;
    END
  END slave3_wb_data_i[15]
  PIN slave3_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 873.160 350.000 873.760 ;
    END
  END slave3_wb_data_i[16]
  PIN slave3_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 889.480 350.000 890.080 ;
    END
  END slave3_wb_data_i[17]
  PIN slave3_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 905.800 350.000 906.400 ;
    END
  END slave3_wb_data_i[18]
  PIN slave3_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 922.120 350.000 922.720 ;
    END
  END slave3_wb_data_i[19]
  PIN slave3_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 612.040 350.000 612.640 ;
    END
  END slave3_wb_data_i[1]
  PIN slave3_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 938.440 350.000 939.040 ;
    END
  END slave3_wb_data_i[20]
  PIN slave3_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 954.760 350.000 955.360 ;
    END
  END slave3_wb_data_i[21]
  PIN slave3_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 971.080 350.000 971.680 ;
    END
  END slave3_wb_data_i[22]
  PIN slave3_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 987.400 350.000 988.000 ;
    END
  END slave3_wb_data_i[23]
  PIN slave3_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 998.280 350.000 998.880 ;
    END
  END slave3_wb_data_i[24]
  PIN slave3_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1009.160 350.000 1009.760 ;
    END
  END slave3_wb_data_i[25]
  PIN slave3_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1020.040 350.000 1020.640 ;
    END
  END slave3_wb_data_i[26]
  PIN slave3_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1030.920 350.000 1031.520 ;
    END
  END slave3_wb_data_i[27]
  PIN slave3_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1041.800 350.000 1042.400 ;
    END
  END slave3_wb_data_i[28]
  PIN slave3_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1052.680 350.000 1053.280 ;
    END
  END slave3_wb_data_i[29]
  PIN slave3_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 633.800 350.000 634.400 ;
    END
  END slave3_wb_data_i[2]
  PIN slave3_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1063.560 350.000 1064.160 ;
    END
  END slave3_wb_data_i[30]
  PIN slave3_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1074.440 350.000 1075.040 ;
    END
  END slave3_wb_data_i[31]
  PIN slave3_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 655.560 350.000 656.160 ;
    END
  END slave3_wb_data_i[3]
  PIN slave3_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 677.320 350.000 677.920 ;
    END
  END slave3_wb_data_i[4]
  PIN slave3_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 693.640 350.000 694.240 ;
    END
  END slave3_wb_data_i[5]
  PIN slave3_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 709.960 350.000 710.560 ;
    END
  END slave3_wb_data_i[6]
  PIN slave3_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 726.280 350.000 726.880 ;
    END
  END slave3_wb_data_i[7]
  PIN slave3_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 742.600 350.000 743.200 ;
    END
  END slave3_wb_data_i[8]
  PIN slave3_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 758.920 350.000 759.520 ;
    END
  END slave3_wb_data_i[9]
  PIN slave3_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 595.720 350.000 596.320 ;
    END
  END slave3_wb_data_o[0]
  PIN slave3_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 780.680 350.000 781.280 ;
    END
  END slave3_wb_data_o[10]
  PIN slave3_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 797.000 350.000 797.600 ;
    END
  END slave3_wb_data_o[11]
  PIN slave3_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 813.320 350.000 813.920 ;
    END
  END slave3_wb_data_o[12]
  PIN slave3_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 829.640 350.000 830.240 ;
    END
  END slave3_wb_data_o[13]
  PIN slave3_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 845.960 350.000 846.560 ;
    END
  END slave3_wb_data_o[14]
  PIN slave3_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 862.280 350.000 862.880 ;
    END
  END slave3_wb_data_o[15]
  PIN slave3_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 878.600 350.000 879.200 ;
    END
  END slave3_wb_data_o[16]
  PIN slave3_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 894.920 350.000 895.520 ;
    END
  END slave3_wb_data_o[17]
  PIN slave3_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 911.240 350.000 911.840 ;
    END
  END slave3_wb_data_o[18]
  PIN slave3_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 927.560 350.000 928.160 ;
    END
  END slave3_wb_data_o[19]
  PIN slave3_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 617.480 350.000 618.080 ;
    END
  END slave3_wb_data_o[1]
  PIN slave3_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 943.880 350.000 944.480 ;
    END
  END slave3_wb_data_o[20]
  PIN slave3_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 960.200 350.000 960.800 ;
    END
  END slave3_wb_data_o[21]
  PIN slave3_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 976.520 350.000 977.120 ;
    END
  END slave3_wb_data_o[22]
  PIN slave3_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 992.840 350.000 993.440 ;
    END
  END slave3_wb_data_o[23]
  PIN slave3_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1003.720 350.000 1004.320 ;
    END
  END slave3_wb_data_o[24]
  PIN slave3_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1014.600 350.000 1015.200 ;
    END
  END slave3_wb_data_o[25]
  PIN slave3_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1025.480 350.000 1026.080 ;
    END
  END slave3_wb_data_o[26]
  PIN slave3_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1036.360 350.000 1036.960 ;
    END
  END slave3_wb_data_o[27]
  PIN slave3_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1047.240 350.000 1047.840 ;
    END
  END slave3_wb_data_o[28]
  PIN slave3_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1058.120 350.000 1058.720 ;
    END
  END slave3_wb_data_o[29]
  PIN slave3_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 639.240 350.000 639.840 ;
    END
  END slave3_wb_data_o[2]
  PIN slave3_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1069.000 350.000 1069.600 ;
    END
  END slave3_wb_data_o[30]
  PIN slave3_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1079.880 350.000 1080.480 ;
    END
  END slave3_wb_data_o[31]
  PIN slave3_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 661.000 350.000 661.600 ;
    END
  END slave3_wb_data_o[3]
  PIN slave3_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 682.760 350.000 683.360 ;
    END
  END slave3_wb_data_o[4]
  PIN slave3_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 699.080 350.000 699.680 ;
    END
  END slave3_wb_data_o[5]
  PIN slave3_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 715.400 350.000 716.000 ;
    END
  END slave3_wb_data_o[6]
  PIN slave3_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 731.720 350.000 732.320 ;
    END
  END slave3_wb_data_o[7]
  PIN slave3_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 748.040 350.000 748.640 ;
    END
  END slave3_wb_data_o[8]
  PIN slave3_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 764.360 350.000 764.960 ;
    END
  END slave3_wb_data_o[9]
  PIN slave3_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 563.080 350.000 563.680 ;
    END
  END slave3_wb_error_o
  PIN slave3_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 601.160 350.000 601.760 ;
    END
  END slave3_wb_sel_i[0]
  PIN slave3_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 622.920 350.000 623.520 ;
    END
  END slave3_wb_sel_i[1]
  PIN slave3_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 644.680 350.000 645.280 ;
    END
  END slave3_wb_sel_i[2]
  PIN slave3_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 666.440 350.000 667.040 ;
    END
  END slave3_wb_sel_i[3]
  PIN slave3_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 568.520 350.000 569.120 ;
    END
  END slave3_wb_stall_o
  PIN slave3_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 573.960 350.000 574.560 ;
    END
  END slave3_wb_stb_i
  PIN slave3_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 579.400 350.000 580.000 ;
    END
  END slave3_wb_we_i
  PIN slave4_wb_ack_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 19.080 350.000 19.680 ;
    END
  END slave4_wb_ack_o
  PIN slave4_wb_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 51.720 350.000 52.320 ;
    END
  END slave4_wb_adr_i[0]
  PIN slave4_wb_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 236.680 350.000 237.280 ;
    END
  END slave4_wb_adr_i[10]
  PIN slave4_wb_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 253.000 350.000 253.600 ;
    END
  END slave4_wb_adr_i[11]
  PIN slave4_wb_adr_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 269.320 350.000 269.920 ;
    END
  END slave4_wb_adr_i[12]
  PIN slave4_wb_adr_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 285.640 350.000 286.240 ;
    END
  END slave4_wb_adr_i[13]
  PIN slave4_wb_adr_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 301.960 350.000 302.560 ;
    END
  END slave4_wb_adr_i[14]
  PIN slave4_wb_adr_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 318.280 350.000 318.880 ;
    END
  END slave4_wb_adr_i[15]
  PIN slave4_wb_adr_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 334.600 350.000 335.200 ;
    END
  END slave4_wb_adr_i[16]
  PIN slave4_wb_adr_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 350.920 350.000 351.520 ;
    END
  END slave4_wb_adr_i[17]
  PIN slave4_wb_adr_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 367.240 350.000 367.840 ;
    END
  END slave4_wb_adr_i[18]
  PIN slave4_wb_adr_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 383.560 350.000 384.160 ;
    END
  END slave4_wb_adr_i[19]
  PIN slave4_wb_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 73.480 350.000 74.080 ;
    END
  END slave4_wb_adr_i[1]
  PIN slave4_wb_adr_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 399.880 350.000 400.480 ;
    END
  END slave4_wb_adr_i[20]
  PIN slave4_wb_adr_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 416.200 350.000 416.800 ;
    END
  END slave4_wb_adr_i[21]
  PIN slave4_wb_adr_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 432.520 350.000 433.120 ;
    END
  END slave4_wb_adr_i[22]
  PIN slave4_wb_adr_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 448.840 350.000 449.440 ;
    END
  END slave4_wb_adr_i[23]
  PIN slave4_wb_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 95.240 350.000 95.840 ;
    END
  END slave4_wb_adr_i[2]
  PIN slave4_wb_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 117.000 350.000 117.600 ;
    END
  END slave4_wb_adr_i[3]
  PIN slave4_wb_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 138.760 350.000 139.360 ;
    END
  END slave4_wb_adr_i[4]
  PIN slave4_wb_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 155.080 350.000 155.680 ;
    END
  END slave4_wb_adr_i[5]
  PIN slave4_wb_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 171.400 350.000 172.000 ;
    END
  END slave4_wb_adr_i[6]
  PIN slave4_wb_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 187.720 350.000 188.320 ;
    END
  END slave4_wb_adr_i[7]
  PIN slave4_wb_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 204.040 350.000 204.640 ;
    END
  END slave4_wb_adr_i[8]
  PIN slave4_wb_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 220.360 350.000 220.960 ;
    END
  END slave4_wb_adr_i[9]
  PIN slave4_wb_cyc_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 24.520 350.000 25.120 ;
    END
  END slave4_wb_cyc_i
  PIN slave4_wb_data_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 57.160 350.000 57.760 ;
    END
  END slave4_wb_data_i[0]
  PIN slave4_wb_data_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 242.120 350.000 242.720 ;
    END
  END slave4_wb_data_i[10]
  PIN slave4_wb_data_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 258.440 350.000 259.040 ;
    END
  END slave4_wb_data_i[11]
  PIN slave4_wb_data_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 274.760 350.000 275.360 ;
    END
  END slave4_wb_data_i[12]
  PIN slave4_wb_data_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 291.080 350.000 291.680 ;
    END
  END slave4_wb_data_i[13]
  PIN slave4_wb_data_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 307.400 350.000 308.000 ;
    END
  END slave4_wb_data_i[14]
  PIN slave4_wb_data_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 323.720 350.000 324.320 ;
    END
  END slave4_wb_data_i[15]
  PIN slave4_wb_data_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 340.040 350.000 340.640 ;
    END
  END slave4_wb_data_i[16]
  PIN slave4_wb_data_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 356.360 350.000 356.960 ;
    END
  END slave4_wb_data_i[17]
  PIN slave4_wb_data_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 372.680 350.000 373.280 ;
    END
  END slave4_wb_data_i[18]
  PIN slave4_wb_data_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 389.000 350.000 389.600 ;
    END
  END slave4_wb_data_i[19]
  PIN slave4_wb_data_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 78.920 350.000 79.520 ;
    END
  END slave4_wb_data_i[1]
  PIN slave4_wb_data_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 405.320 350.000 405.920 ;
    END
  END slave4_wb_data_i[20]
  PIN slave4_wb_data_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 421.640 350.000 422.240 ;
    END
  END slave4_wb_data_i[21]
  PIN slave4_wb_data_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 437.960 350.000 438.560 ;
    END
  END slave4_wb_data_i[22]
  PIN slave4_wb_data_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 454.280 350.000 454.880 ;
    END
  END slave4_wb_data_i[23]
  PIN slave4_wb_data_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 465.160 350.000 465.760 ;
    END
  END slave4_wb_data_i[24]
  PIN slave4_wb_data_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 476.040 350.000 476.640 ;
    END
  END slave4_wb_data_i[25]
  PIN slave4_wb_data_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 486.920 350.000 487.520 ;
    END
  END slave4_wb_data_i[26]
  PIN slave4_wb_data_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 497.800 350.000 498.400 ;
    END
  END slave4_wb_data_i[27]
  PIN slave4_wb_data_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 508.680 350.000 509.280 ;
    END
  END slave4_wb_data_i[28]
  PIN slave4_wb_data_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 519.560 350.000 520.160 ;
    END
  END slave4_wb_data_i[29]
  PIN slave4_wb_data_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 100.680 350.000 101.280 ;
    END
  END slave4_wb_data_i[2]
  PIN slave4_wb_data_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 530.440 350.000 531.040 ;
    END
  END slave4_wb_data_i[30]
  PIN slave4_wb_data_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 541.320 350.000 541.920 ;
    END
  END slave4_wb_data_i[31]
  PIN slave4_wb_data_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 122.440 350.000 123.040 ;
    END
  END slave4_wb_data_i[3]
  PIN slave4_wb_data_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 144.200 350.000 144.800 ;
    END
  END slave4_wb_data_i[4]
  PIN slave4_wb_data_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 160.520 350.000 161.120 ;
    END
  END slave4_wb_data_i[5]
  PIN slave4_wb_data_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 176.840 350.000 177.440 ;
    END
  END slave4_wb_data_i[6]
  PIN slave4_wb_data_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 193.160 350.000 193.760 ;
    END
  END slave4_wb_data_i[7]
  PIN slave4_wb_data_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 209.480 350.000 210.080 ;
    END
  END slave4_wb_data_i[8]
  PIN slave4_wb_data_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 225.800 350.000 226.400 ;
    END
  END slave4_wb_data_i[9]
  PIN slave4_wb_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 62.600 350.000 63.200 ;
    END
  END slave4_wb_data_o[0]
  PIN slave4_wb_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 247.560 350.000 248.160 ;
    END
  END slave4_wb_data_o[10]
  PIN slave4_wb_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 263.880 350.000 264.480 ;
    END
  END slave4_wb_data_o[11]
  PIN slave4_wb_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 280.200 350.000 280.800 ;
    END
  END slave4_wb_data_o[12]
  PIN slave4_wb_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 296.520 350.000 297.120 ;
    END
  END slave4_wb_data_o[13]
  PIN slave4_wb_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 312.840 350.000 313.440 ;
    END
  END slave4_wb_data_o[14]
  PIN slave4_wb_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 329.160 350.000 329.760 ;
    END
  END slave4_wb_data_o[15]
  PIN slave4_wb_data_o[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 345.480 350.000 346.080 ;
    END
  END slave4_wb_data_o[16]
  PIN slave4_wb_data_o[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 361.800 350.000 362.400 ;
    END
  END slave4_wb_data_o[17]
  PIN slave4_wb_data_o[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 378.120 350.000 378.720 ;
    END
  END slave4_wb_data_o[18]
  PIN slave4_wb_data_o[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 394.440 350.000 395.040 ;
    END
  END slave4_wb_data_o[19]
  PIN slave4_wb_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 84.360 350.000 84.960 ;
    END
  END slave4_wb_data_o[1]
  PIN slave4_wb_data_o[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 410.760 350.000 411.360 ;
    END
  END slave4_wb_data_o[20]
  PIN slave4_wb_data_o[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 427.080 350.000 427.680 ;
    END
  END slave4_wb_data_o[21]
  PIN slave4_wb_data_o[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 443.400 350.000 444.000 ;
    END
  END slave4_wb_data_o[22]
  PIN slave4_wb_data_o[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 459.720 350.000 460.320 ;
    END
  END slave4_wb_data_o[23]
  PIN slave4_wb_data_o[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 470.600 350.000 471.200 ;
    END
  END slave4_wb_data_o[24]
  PIN slave4_wb_data_o[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 481.480 350.000 482.080 ;
    END
  END slave4_wb_data_o[25]
  PIN slave4_wb_data_o[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 492.360 350.000 492.960 ;
    END
  END slave4_wb_data_o[26]
  PIN slave4_wb_data_o[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 503.240 350.000 503.840 ;
    END
  END slave4_wb_data_o[27]
  PIN slave4_wb_data_o[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 514.120 350.000 514.720 ;
    END
  END slave4_wb_data_o[28]
  PIN slave4_wb_data_o[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 525.000 350.000 525.600 ;
    END
  END slave4_wb_data_o[29]
  PIN slave4_wb_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 106.120 350.000 106.720 ;
    END
  END slave4_wb_data_o[2]
  PIN slave4_wb_data_o[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 535.880 350.000 536.480 ;
    END
  END slave4_wb_data_o[30]
  PIN slave4_wb_data_o[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 546.760 350.000 547.360 ;
    END
  END slave4_wb_data_o[31]
  PIN slave4_wb_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 127.880 350.000 128.480 ;
    END
  END slave4_wb_data_o[3]
  PIN slave4_wb_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 149.640 350.000 150.240 ;
    END
  END slave4_wb_data_o[4]
  PIN slave4_wb_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 165.960 350.000 166.560 ;
    END
  END slave4_wb_data_o[5]
  PIN slave4_wb_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 182.280 350.000 182.880 ;
    END
  END slave4_wb_data_o[6]
  PIN slave4_wb_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 198.600 350.000 199.200 ;
    END
  END slave4_wb_data_o[7]
  PIN slave4_wb_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 214.920 350.000 215.520 ;
    END
  END slave4_wb_data_o[8]
  PIN slave4_wb_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 231.240 350.000 231.840 ;
    END
  END slave4_wb_data_o[9]
  PIN slave4_wb_error_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 29.960 350.000 30.560 ;
    END
  END slave4_wb_error_o
  PIN slave4_wb_sel_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 68.040 350.000 68.640 ;
    END
  END slave4_wb_sel_i[0]
  PIN slave4_wb_sel_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 89.800 350.000 90.400 ;
    END
  END slave4_wb_sel_i[1]
  PIN slave4_wb_sel_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 111.560 350.000 112.160 ;
    END
  END slave4_wb_sel_i[2]
  PIN slave4_wb_sel_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 133.320 350.000 133.920 ;
    END
  END slave4_wb_sel_i[3]
  PIN slave4_wb_stall_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 35.400 350.000 36.000 ;
    END
  END slave4_wb_stall_o
  PIN slave4_wb_stb_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 40.840 350.000 41.440 ;
    END
  END slave4_wb_stb_i
  PIN slave4_wb_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 46.280 350.000 46.880 ;
    END
  END slave4_wb_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1088.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1088.240 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 1088.085 ;
      LAYER met1 ;
        RECT 0.070 4.460 345.390 1096.460 ;
      LAYER met2 ;
        RECT 0.100 1095.720 18.210 1097.250 ;
        RECT 19.050 1095.720 21.430 1097.250 ;
        RECT 22.270 1095.720 24.650 1097.250 ;
        RECT 25.490 1095.720 27.870 1097.250 ;
        RECT 28.710 1095.720 31.090 1097.250 ;
        RECT 31.930 1095.720 34.310 1097.250 ;
        RECT 35.150 1095.720 37.530 1097.250 ;
        RECT 38.370 1095.720 40.750 1097.250 ;
        RECT 41.590 1095.720 43.970 1097.250 ;
        RECT 44.810 1095.720 47.190 1097.250 ;
        RECT 48.030 1095.720 50.410 1097.250 ;
        RECT 51.250 1095.720 53.630 1097.250 ;
        RECT 54.470 1095.720 56.850 1097.250 ;
        RECT 57.690 1095.720 60.070 1097.250 ;
        RECT 60.910 1095.720 63.290 1097.250 ;
        RECT 64.130 1095.720 66.510 1097.250 ;
        RECT 67.350 1095.720 69.730 1097.250 ;
        RECT 70.570 1095.720 72.950 1097.250 ;
        RECT 73.790 1095.720 76.170 1097.250 ;
        RECT 77.010 1095.720 79.390 1097.250 ;
        RECT 80.230 1095.720 82.610 1097.250 ;
        RECT 83.450 1095.720 85.830 1097.250 ;
        RECT 86.670 1095.720 89.050 1097.250 ;
        RECT 89.890 1095.720 92.270 1097.250 ;
        RECT 93.110 1095.720 95.490 1097.250 ;
        RECT 96.330 1095.720 98.710 1097.250 ;
        RECT 99.550 1095.720 101.930 1097.250 ;
        RECT 102.770 1095.720 105.150 1097.250 ;
        RECT 105.990 1095.720 108.370 1097.250 ;
        RECT 109.210 1095.720 111.590 1097.250 ;
        RECT 112.430 1095.720 114.810 1097.250 ;
        RECT 115.650 1095.720 118.030 1097.250 ;
        RECT 118.870 1095.720 121.250 1097.250 ;
        RECT 122.090 1095.720 124.470 1097.250 ;
        RECT 125.310 1095.720 127.690 1097.250 ;
        RECT 128.530 1095.720 130.910 1097.250 ;
        RECT 131.750 1095.720 134.130 1097.250 ;
        RECT 134.970 1095.720 137.350 1097.250 ;
        RECT 138.190 1095.720 140.570 1097.250 ;
        RECT 141.410 1095.720 143.790 1097.250 ;
        RECT 144.630 1095.720 147.010 1097.250 ;
        RECT 147.850 1095.720 150.230 1097.250 ;
        RECT 151.070 1095.720 153.450 1097.250 ;
        RECT 154.290 1095.720 156.670 1097.250 ;
        RECT 157.510 1095.720 159.890 1097.250 ;
        RECT 160.730 1095.720 163.110 1097.250 ;
        RECT 163.950 1095.720 166.330 1097.250 ;
        RECT 167.170 1095.720 169.550 1097.250 ;
        RECT 170.390 1095.720 172.770 1097.250 ;
        RECT 173.610 1095.720 175.990 1097.250 ;
        RECT 176.830 1095.720 179.210 1097.250 ;
        RECT 180.050 1095.720 182.430 1097.250 ;
        RECT 183.270 1095.720 185.650 1097.250 ;
        RECT 186.490 1095.720 188.870 1097.250 ;
        RECT 189.710 1095.720 192.090 1097.250 ;
        RECT 192.930 1095.720 195.310 1097.250 ;
        RECT 196.150 1095.720 198.530 1097.250 ;
        RECT 199.370 1095.720 201.750 1097.250 ;
        RECT 202.590 1095.720 204.970 1097.250 ;
        RECT 205.810 1095.720 208.190 1097.250 ;
        RECT 209.030 1095.720 211.410 1097.250 ;
        RECT 212.250 1095.720 214.630 1097.250 ;
        RECT 215.470 1095.720 217.850 1097.250 ;
        RECT 218.690 1095.720 221.070 1097.250 ;
        RECT 221.910 1095.720 224.290 1097.250 ;
        RECT 225.130 1095.720 227.510 1097.250 ;
        RECT 228.350 1095.720 230.730 1097.250 ;
        RECT 231.570 1095.720 233.950 1097.250 ;
        RECT 234.790 1095.720 237.170 1097.250 ;
        RECT 238.010 1095.720 240.390 1097.250 ;
        RECT 241.230 1095.720 243.610 1097.250 ;
        RECT 244.450 1095.720 246.830 1097.250 ;
        RECT 247.670 1095.720 250.050 1097.250 ;
        RECT 250.890 1095.720 253.270 1097.250 ;
        RECT 254.110 1095.720 256.490 1097.250 ;
        RECT 257.330 1095.720 259.710 1097.250 ;
        RECT 260.550 1095.720 262.930 1097.250 ;
        RECT 263.770 1095.720 266.150 1097.250 ;
        RECT 266.990 1095.720 269.370 1097.250 ;
        RECT 270.210 1095.720 272.590 1097.250 ;
        RECT 273.430 1095.720 275.810 1097.250 ;
        RECT 276.650 1095.720 279.030 1097.250 ;
        RECT 279.870 1095.720 282.250 1097.250 ;
        RECT 283.090 1095.720 285.470 1097.250 ;
        RECT 286.310 1095.720 288.690 1097.250 ;
        RECT 289.530 1095.720 291.910 1097.250 ;
        RECT 292.750 1095.720 295.130 1097.250 ;
        RECT 295.970 1095.720 298.350 1097.250 ;
        RECT 299.190 1095.720 301.570 1097.250 ;
        RECT 302.410 1095.720 304.790 1097.250 ;
        RECT 305.630 1095.720 308.010 1097.250 ;
        RECT 308.850 1095.720 311.230 1097.250 ;
        RECT 312.070 1095.720 314.450 1097.250 ;
        RECT 315.290 1095.720 317.670 1097.250 ;
        RECT 318.510 1095.720 320.890 1097.250 ;
        RECT 321.730 1095.720 324.110 1097.250 ;
        RECT 324.950 1095.720 327.330 1097.250 ;
        RECT 328.170 1095.720 330.550 1097.250 ;
        RECT 331.390 1095.720 345.370 1097.250 ;
        RECT 0.100 4.280 345.370 1095.720 ;
        RECT 0.100 3.670 10.390 4.280 ;
        RECT 11.230 3.670 13.150 4.280 ;
        RECT 13.990 3.670 15.910 4.280 ;
        RECT 16.750 3.670 18.670 4.280 ;
        RECT 19.510 3.670 21.430 4.280 ;
        RECT 22.270 3.670 24.190 4.280 ;
        RECT 25.030 3.670 26.950 4.280 ;
        RECT 27.790 3.670 29.710 4.280 ;
        RECT 30.550 3.670 32.470 4.280 ;
        RECT 33.310 3.670 35.230 4.280 ;
        RECT 36.070 3.670 37.990 4.280 ;
        RECT 38.830 3.670 40.750 4.280 ;
        RECT 41.590 3.670 43.510 4.280 ;
        RECT 44.350 3.670 46.270 4.280 ;
        RECT 47.110 3.670 49.030 4.280 ;
        RECT 49.870 3.670 51.790 4.280 ;
        RECT 52.630 3.670 54.550 4.280 ;
        RECT 55.390 3.670 57.310 4.280 ;
        RECT 58.150 3.670 60.070 4.280 ;
        RECT 60.910 3.670 62.830 4.280 ;
        RECT 63.670 3.670 65.590 4.280 ;
        RECT 66.430 3.670 68.350 4.280 ;
        RECT 69.190 3.670 71.110 4.280 ;
        RECT 71.950 3.670 73.870 4.280 ;
        RECT 74.710 3.670 76.630 4.280 ;
        RECT 77.470 3.670 79.390 4.280 ;
        RECT 80.230 3.670 82.150 4.280 ;
        RECT 82.990 3.670 84.910 4.280 ;
        RECT 85.750 3.670 87.670 4.280 ;
        RECT 88.510 3.670 90.430 4.280 ;
        RECT 91.270 3.670 93.190 4.280 ;
        RECT 94.030 3.670 95.950 4.280 ;
        RECT 96.790 3.670 98.710 4.280 ;
        RECT 99.550 3.670 101.470 4.280 ;
        RECT 102.310 3.670 104.230 4.280 ;
        RECT 105.070 3.670 106.990 4.280 ;
        RECT 107.830 3.670 109.750 4.280 ;
        RECT 110.590 3.670 112.510 4.280 ;
        RECT 113.350 3.670 115.270 4.280 ;
        RECT 116.110 3.670 118.030 4.280 ;
        RECT 118.870 3.670 120.790 4.280 ;
        RECT 121.630 3.670 123.550 4.280 ;
        RECT 124.390 3.670 126.310 4.280 ;
        RECT 127.150 3.670 129.070 4.280 ;
        RECT 129.910 3.670 131.830 4.280 ;
        RECT 132.670 3.670 134.590 4.280 ;
        RECT 135.430 3.670 137.350 4.280 ;
        RECT 138.190 3.670 140.110 4.280 ;
        RECT 140.950 3.670 142.870 4.280 ;
        RECT 143.710 3.670 145.630 4.280 ;
        RECT 146.470 3.670 148.390 4.280 ;
        RECT 149.230 3.670 151.150 4.280 ;
        RECT 151.990 3.670 153.910 4.280 ;
        RECT 154.750 3.670 156.670 4.280 ;
        RECT 157.510 3.670 159.430 4.280 ;
        RECT 160.270 3.670 162.190 4.280 ;
        RECT 163.030 3.670 164.950 4.280 ;
        RECT 165.790 3.670 167.710 4.280 ;
        RECT 168.550 3.670 170.470 4.280 ;
        RECT 171.310 3.670 173.230 4.280 ;
        RECT 174.070 3.670 175.990 4.280 ;
        RECT 176.830 3.670 178.750 4.280 ;
        RECT 179.590 3.670 181.510 4.280 ;
        RECT 182.350 3.670 184.270 4.280 ;
        RECT 185.110 3.670 187.030 4.280 ;
        RECT 187.870 3.670 189.790 4.280 ;
        RECT 190.630 3.670 192.550 4.280 ;
        RECT 193.390 3.670 195.310 4.280 ;
        RECT 196.150 3.670 198.070 4.280 ;
        RECT 198.910 3.670 200.830 4.280 ;
        RECT 201.670 3.670 203.590 4.280 ;
        RECT 204.430 3.670 206.350 4.280 ;
        RECT 207.190 3.670 209.110 4.280 ;
        RECT 209.950 3.670 211.870 4.280 ;
        RECT 212.710 3.670 214.630 4.280 ;
        RECT 215.470 3.670 217.390 4.280 ;
        RECT 218.230 3.670 220.150 4.280 ;
        RECT 220.990 3.670 222.910 4.280 ;
        RECT 223.750 3.670 225.670 4.280 ;
        RECT 226.510 3.670 228.430 4.280 ;
        RECT 229.270 3.670 231.190 4.280 ;
        RECT 232.030 3.670 233.950 4.280 ;
        RECT 234.790 3.670 236.710 4.280 ;
        RECT 237.550 3.670 239.470 4.280 ;
        RECT 240.310 3.670 242.230 4.280 ;
        RECT 243.070 3.670 244.990 4.280 ;
        RECT 245.830 3.670 247.750 4.280 ;
        RECT 248.590 3.670 250.510 4.280 ;
        RECT 251.350 3.670 253.270 4.280 ;
        RECT 254.110 3.670 256.030 4.280 ;
        RECT 256.870 3.670 258.790 4.280 ;
        RECT 259.630 3.670 261.550 4.280 ;
        RECT 262.390 3.670 264.310 4.280 ;
        RECT 265.150 3.670 267.070 4.280 ;
        RECT 267.910 3.670 269.830 4.280 ;
        RECT 270.670 3.670 272.590 4.280 ;
        RECT 273.430 3.670 275.350 4.280 ;
        RECT 276.190 3.670 278.110 4.280 ;
        RECT 278.950 3.670 280.870 4.280 ;
        RECT 281.710 3.670 283.630 4.280 ;
        RECT 284.470 3.670 286.390 4.280 ;
        RECT 287.230 3.670 289.150 4.280 ;
        RECT 289.990 3.670 291.910 4.280 ;
        RECT 292.750 3.670 294.670 4.280 ;
        RECT 295.510 3.670 297.430 4.280 ;
        RECT 298.270 3.670 300.190 4.280 ;
        RECT 301.030 3.670 302.950 4.280 ;
        RECT 303.790 3.670 305.710 4.280 ;
        RECT 306.550 3.670 308.470 4.280 ;
        RECT 309.310 3.670 311.230 4.280 ;
        RECT 312.070 3.670 313.990 4.280 ;
        RECT 314.830 3.670 316.750 4.280 ;
        RECT 317.590 3.670 319.510 4.280 ;
        RECT 320.350 3.670 322.270 4.280 ;
        RECT 323.110 3.670 325.030 4.280 ;
        RECT 325.870 3.670 327.790 4.280 ;
        RECT 328.630 3.670 330.550 4.280 ;
        RECT 331.390 3.670 333.310 4.280 ;
        RECT 334.150 3.670 336.070 4.280 ;
        RECT 336.910 3.670 338.830 4.280 ;
        RECT 339.670 3.670 345.370 4.280 ;
      LAYER met3 ;
        RECT 4.400 1091.720 346.000 1092.585 ;
        RECT 3.950 1090.400 346.000 1091.720 ;
        RECT 4.400 1089.000 346.000 1090.400 ;
        RECT 3.950 1087.680 346.000 1089.000 ;
        RECT 4.400 1086.280 346.000 1087.680 ;
        RECT 3.950 1084.960 346.000 1086.280 ;
        RECT 4.400 1083.560 346.000 1084.960 ;
        RECT 3.950 1082.240 346.000 1083.560 ;
        RECT 4.400 1080.880 346.000 1082.240 ;
        RECT 4.400 1080.840 345.600 1080.880 ;
        RECT 3.950 1079.520 345.600 1080.840 ;
        RECT 4.400 1079.480 345.600 1079.520 ;
        RECT 4.400 1078.120 346.000 1079.480 ;
        RECT 3.950 1076.800 346.000 1078.120 ;
        RECT 4.400 1075.440 346.000 1076.800 ;
        RECT 4.400 1075.400 345.600 1075.440 ;
        RECT 3.950 1074.080 345.600 1075.400 ;
        RECT 4.400 1074.040 345.600 1074.080 ;
        RECT 4.400 1072.680 346.000 1074.040 ;
        RECT 3.950 1071.360 346.000 1072.680 ;
        RECT 4.400 1070.000 346.000 1071.360 ;
        RECT 4.400 1069.960 345.600 1070.000 ;
        RECT 3.950 1068.640 345.600 1069.960 ;
        RECT 4.400 1068.600 345.600 1068.640 ;
        RECT 4.400 1067.240 346.000 1068.600 ;
        RECT 3.950 1065.920 346.000 1067.240 ;
        RECT 4.400 1064.560 346.000 1065.920 ;
        RECT 4.400 1064.520 345.600 1064.560 ;
        RECT 3.950 1063.200 345.600 1064.520 ;
        RECT 4.400 1063.160 345.600 1063.200 ;
        RECT 4.400 1061.800 346.000 1063.160 ;
        RECT 3.950 1060.480 346.000 1061.800 ;
        RECT 4.400 1059.120 346.000 1060.480 ;
        RECT 4.400 1059.080 345.600 1059.120 ;
        RECT 3.950 1057.760 345.600 1059.080 ;
        RECT 4.400 1057.720 345.600 1057.760 ;
        RECT 4.400 1056.360 346.000 1057.720 ;
        RECT 3.950 1055.040 346.000 1056.360 ;
        RECT 4.400 1053.680 346.000 1055.040 ;
        RECT 4.400 1053.640 345.600 1053.680 ;
        RECT 3.950 1052.320 345.600 1053.640 ;
        RECT 4.400 1052.280 345.600 1052.320 ;
        RECT 4.400 1050.920 346.000 1052.280 ;
        RECT 3.950 1049.600 346.000 1050.920 ;
        RECT 4.400 1048.240 346.000 1049.600 ;
        RECT 4.400 1048.200 345.600 1048.240 ;
        RECT 3.950 1046.880 345.600 1048.200 ;
        RECT 4.400 1046.840 345.600 1046.880 ;
        RECT 4.400 1045.480 346.000 1046.840 ;
        RECT 3.950 1044.160 346.000 1045.480 ;
        RECT 4.400 1042.800 346.000 1044.160 ;
        RECT 4.400 1042.760 345.600 1042.800 ;
        RECT 3.950 1041.440 345.600 1042.760 ;
        RECT 4.400 1041.400 345.600 1041.440 ;
        RECT 4.400 1040.040 346.000 1041.400 ;
        RECT 3.950 1038.720 346.000 1040.040 ;
        RECT 4.400 1037.360 346.000 1038.720 ;
        RECT 4.400 1037.320 345.600 1037.360 ;
        RECT 3.950 1036.000 345.600 1037.320 ;
        RECT 4.400 1035.960 345.600 1036.000 ;
        RECT 4.400 1034.600 346.000 1035.960 ;
        RECT 3.950 1033.280 346.000 1034.600 ;
        RECT 4.400 1031.920 346.000 1033.280 ;
        RECT 4.400 1031.880 345.600 1031.920 ;
        RECT 3.950 1030.560 345.600 1031.880 ;
        RECT 4.400 1030.520 345.600 1030.560 ;
        RECT 4.400 1029.160 346.000 1030.520 ;
        RECT 3.950 1027.840 346.000 1029.160 ;
        RECT 4.400 1026.480 346.000 1027.840 ;
        RECT 4.400 1026.440 345.600 1026.480 ;
        RECT 3.950 1025.120 345.600 1026.440 ;
        RECT 4.400 1025.080 345.600 1025.120 ;
        RECT 4.400 1023.720 346.000 1025.080 ;
        RECT 3.950 1022.400 346.000 1023.720 ;
        RECT 4.400 1021.040 346.000 1022.400 ;
        RECT 4.400 1021.000 345.600 1021.040 ;
        RECT 3.950 1019.680 345.600 1021.000 ;
        RECT 4.400 1019.640 345.600 1019.680 ;
        RECT 4.400 1018.280 346.000 1019.640 ;
        RECT 3.950 1016.960 346.000 1018.280 ;
        RECT 4.400 1015.600 346.000 1016.960 ;
        RECT 4.400 1015.560 345.600 1015.600 ;
        RECT 3.950 1014.240 345.600 1015.560 ;
        RECT 4.400 1014.200 345.600 1014.240 ;
        RECT 4.400 1012.840 346.000 1014.200 ;
        RECT 3.950 1011.520 346.000 1012.840 ;
        RECT 4.400 1010.160 346.000 1011.520 ;
        RECT 4.400 1010.120 345.600 1010.160 ;
        RECT 3.950 1008.800 345.600 1010.120 ;
        RECT 4.400 1008.760 345.600 1008.800 ;
        RECT 4.400 1007.400 346.000 1008.760 ;
        RECT 3.950 1006.080 346.000 1007.400 ;
        RECT 4.400 1004.720 346.000 1006.080 ;
        RECT 4.400 1004.680 345.600 1004.720 ;
        RECT 3.950 1003.360 345.600 1004.680 ;
        RECT 4.400 1003.320 345.600 1003.360 ;
        RECT 4.400 1001.960 346.000 1003.320 ;
        RECT 3.950 1000.640 346.000 1001.960 ;
        RECT 4.400 999.280 346.000 1000.640 ;
        RECT 4.400 999.240 345.600 999.280 ;
        RECT 3.950 997.920 345.600 999.240 ;
        RECT 4.400 997.880 345.600 997.920 ;
        RECT 4.400 996.520 346.000 997.880 ;
        RECT 3.950 995.200 346.000 996.520 ;
        RECT 4.400 993.840 346.000 995.200 ;
        RECT 4.400 993.800 345.600 993.840 ;
        RECT 3.950 992.480 345.600 993.800 ;
        RECT 4.400 992.440 345.600 992.480 ;
        RECT 4.400 991.080 346.000 992.440 ;
        RECT 3.950 989.760 346.000 991.080 ;
        RECT 4.400 988.400 346.000 989.760 ;
        RECT 4.400 988.360 345.600 988.400 ;
        RECT 3.950 987.040 345.600 988.360 ;
        RECT 4.400 987.000 345.600 987.040 ;
        RECT 4.400 985.640 346.000 987.000 ;
        RECT 3.950 984.320 346.000 985.640 ;
        RECT 4.400 982.960 346.000 984.320 ;
        RECT 4.400 982.920 345.600 982.960 ;
        RECT 3.950 981.600 345.600 982.920 ;
        RECT 4.400 981.560 345.600 981.600 ;
        RECT 4.400 980.200 346.000 981.560 ;
        RECT 3.950 978.880 346.000 980.200 ;
        RECT 4.400 977.520 346.000 978.880 ;
        RECT 4.400 977.480 345.600 977.520 ;
        RECT 3.950 976.160 345.600 977.480 ;
        RECT 4.400 976.120 345.600 976.160 ;
        RECT 4.400 974.760 346.000 976.120 ;
        RECT 3.950 973.440 346.000 974.760 ;
        RECT 4.400 972.080 346.000 973.440 ;
        RECT 4.400 972.040 345.600 972.080 ;
        RECT 3.950 970.720 345.600 972.040 ;
        RECT 4.400 970.680 345.600 970.720 ;
        RECT 4.400 969.320 346.000 970.680 ;
        RECT 3.950 968.000 346.000 969.320 ;
        RECT 4.400 966.640 346.000 968.000 ;
        RECT 4.400 966.600 345.600 966.640 ;
        RECT 3.950 965.280 345.600 966.600 ;
        RECT 4.400 965.240 345.600 965.280 ;
        RECT 4.400 963.880 346.000 965.240 ;
        RECT 3.950 962.560 346.000 963.880 ;
        RECT 4.400 961.200 346.000 962.560 ;
        RECT 4.400 961.160 345.600 961.200 ;
        RECT 3.950 959.840 345.600 961.160 ;
        RECT 4.400 959.800 345.600 959.840 ;
        RECT 4.400 958.440 346.000 959.800 ;
        RECT 3.950 957.120 346.000 958.440 ;
        RECT 4.400 955.760 346.000 957.120 ;
        RECT 4.400 955.720 345.600 955.760 ;
        RECT 3.950 954.400 345.600 955.720 ;
        RECT 4.400 954.360 345.600 954.400 ;
        RECT 4.400 953.000 346.000 954.360 ;
        RECT 3.950 951.680 346.000 953.000 ;
        RECT 4.400 950.320 346.000 951.680 ;
        RECT 4.400 950.280 345.600 950.320 ;
        RECT 3.950 948.960 345.600 950.280 ;
        RECT 4.400 948.920 345.600 948.960 ;
        RECT 4.400 947.560 346.000 948.920 ;
        RECT 3.950 946.240 346.000 947.560 ;
        RECT 4.400 944.880 346.000 946.240 ;
        RECT 4.400 944.840 345.600 944.880 ;
        RECT 3.950 943.520 345.600 944.840 ;
        RECT 4.400 943.480 345.600 943.520 ;
        RECT 4.400 942.120 346.000 943.480 ;
        RECT 3.950 940.800 346.000 942.120 ;
        RECT 4.400 939.440 346.000 940.800 ;
        RECT 4.400 939.400 345.600 939.440 ;
        RECT 3.950 938.080 345.600 939.400 ;
        RECT 4.400 938.040 345.600 938.080 ;
        RECT 4.400 936.680 346.000 938.040 ;
        RECT 3.950 935.360 346.000 936.680 ;
        RECT 4.400 934.000 346.000 935.360 ;
        RECT 4.400 933.960 345.600 934.000 ;
        RECT 3.950 932.640 345.600 933.960 ;
        RECT 4.400 932.600 345.600 932.640 ;
        RECT 4.400 931.240 346.000 932.600 ;
        RECT 3.950 929.920 346.000 931.240 ;
        RECT 4.400 928.560 346.000 929.920 ;
        RECT 4.400 928.520 345.600 928.560 ;
        RECT 3.950 927.200 345.600 928.520 ;
        RECT 4.400 927.160 345.600 927.200 ;
        RECT 4.400 925.800 346.000 927.160 ;
        RECT 3.950 924.480 346.000 925.800 ;
        RECT 4.400 923.120 346.000 924.480 ;
        RECT 4.400 923.080 345.600 923.120 ;
        RECT 3.950 921.760 345.600 923.080 ;
        RECT 4.400 921.720 345.600 921.760 ;
        RECT 4.400 920.360 346.000 921.720 ;
        RECT 3.950 919.040 346.000 920.360 ;
        RECT 4.400 917.680 346.000 919.040 ;
        RECT 4.400 917.640 345.600 917.680 ;
        RECT 3.950 916.320 345.600 917.640 ;
        RECT 4.400 916.280 345.600 916.320 ;
        RECT 4.400 914.920 346.000 916.280 ;
        RECT 3.950 913.600 346.000 914.920 ;
        RECT 4.400 912.240 346.000 913.600 ;
        RECT 4.400 912.200 345.600 912.240 ;
        RECT 3.950 910.880 345.600 912.200 ;
        RECT 4.400 910.840 345.600 910.880 ;
        RECT 4.400 909.480 346.000 910.840 ;
        RECT 3.950 908.160 346.000 909.480 ;
        RECT 4.400 906.800 346.000 908.160 ;
        RECT 4.400 906.760 345.600 906.800 ;
        RECT 3.950 905.440 345.600 906.760 ;
        RECT 4.400 905.400 345.600 905.440 ;
        RECT 4.400 904.040 346.000 905.400 ;
        RECT 3.950 902.720 346.000 904.040 ;
        RECT 4.400 901.360 346.000 902.720 ;
        RECT 4.400 901.320 345.600 901.360 ;
        RECT 3.950 900.000 345.600 901.320 ;
        RECT 4.400 899.960 345.600 900.000 ;
        RECT 4.400 898.600 346.000 899.960 ;
        RECT 3.950 897.280 346.000 898.600 ;
        RECT 4.400 895.920 346.000 897.280 ;
        RECT 4.400 895.880 345.600 895.920 ;
        RECT 3.950 894.560 345.600 895.880 ;
        RECT 4.400 894.520 345.600 894.560 ;
        RECT 4.400 893.160 346.000 894.520 ;
        RECT 3.950 891.840 346.000 893.160 ;
        RECT 4.400 890.480 346.000 891.840 ;
        RECT 4.400 890.440 345.600 890.480 ;
        RECT 3.950 889.120 345.600 890.440 ;
        RECT 4.400 889.080 345.600 889.120 ;
        RECT 4.400 887.720 346.000 889.080 ;
        RECT 3.950 886.400 346.000 887.720 ;
        RECT 4.400 885.040 346.000 886.400 ;
        RECT 4.400 885.000 345.600 885.040 ;
        RECT 3.950 883.680 345.600 885.000 ;
        RECT 4.400 883.640 345.600 883.680 ;
        RECT 4.400 882.280 346.000 883.640 ;
        RECT 3.950 880.960 346.000 882.280 ;
        RECT 4.400 879.600 346.000 880.960 ;
        RECT 4.400 879.560 345.600 879.600 ;
        RECT 3.950 878.240 345.600 879.560 ;
        RECT 4.400 878.200 345.600 878.240 ;
        RECT 4.400 876.840 346.000 878.200 ;
        RECT 3.950 875.520 346.000 876.840 ;
        RECT 4.400 874.160 346.000 875.520 ;
        RECT 4.400 874.120 345.600 874.160 ;
        RECT 3.950 872.800 345.600 874.120 ;
        RECT 4.400 872.760 345.600 872.800 ;
        RECT 4.400 871.400 346.000 872.760 ;
        RECT 3.950 870.080 346.000 871.400 ;
        RECT 4.400 868.720 346.000 870.080 ;
        RECT 4.400 868.680 345.600 868.720 ;
        RECT 3.950 867.360 345.600 868.680 ;
        RECT 4.400 867.320 345.600 867.360 ;
        RECT 4.400 865.960 346.000 867.320 ;
        RECT 3.950 864.640 346.000 865.960 ;
        RECT 4.400 863.280 346.000 864.640 ;
        RECT 4.400 863.240 345.600 863.280 ;
        RECT 3.950 861.920 345.600 863.240 ;
        RECT 4.400 861.880 345.600 861.920 ;
        RECT 4.400 860.520 346.000 861.880 ;
        RECT 3.950 859.200 346.000 860.520 ;
        RECT 4.400 857.840 346.000 859.200 ;
        RECT 4.400 857.800 345.600 857.840 ;
        RECT 3.950 856.480 345.600 857.800 ;
        RECT 4.400 856.440 345.600 856.480 ;
        RECT 4.400 855.080 346.000 856.440 ;
        RECT 3.950 853.760 346.000 855.080 ;
        RECT 4.400 852.400 346.000 853.760 ;
        RECT 4.400 852.360 345.600 852.400 ;
        RECT 3.950 851.040 345.600 852.360 ;
        RECT 4.400 851.000 345.600 851.040 ;
        RECT 4.400 849.640 346.000 851.000 ;
        RECT 3.950 848.320 346.000 849.640 ;
        RECT 4.400 846.960 346.000 848.320 ;
        RECT 4.400 846.920 345.600 846.960 ;
        RECT 3.950 845.600 345.600 846.920 ;
        RECT 4.400 845.560 345.600 845.600 ;
        RECT 4.400 844.200 346.000 845.560 ;
        RECT 3.950 842.880 346.000 844.200 ;
        RECT 4.400 841.520 346.000 842.880 ;
        RECT 4.400 841.480 345.600 841.520 ;
        RECT 3.950 840.160 345.600 841.480 ;
        RECT 4.400 840.120 345.600 840.160 ;
        RECT 4.400 838.760 346.000 840.120 ;
        RECT 3.950 837.440 346.000 838.760 ;
        RECT 4.400 836.080 346.000 837.440 ;
        RECT 4.400 836.040 345.600 836.080 ;
        RECT 3.950 834.720 345.600 836.040 ;
        RECT 4.400 834.680 345.600 834.720 ;
        RECT 4.400 833.320 346.000 834.680 ;
        RECT 3.950 832.000 346.000 833.320 ;
        RECT 4.400 830.640 346.000 832.000 ;
        RECT 4.400 830.600 345.600 830.640 ;
        RECT 3.950 829.280 345.600 830.600 ;
        RECT 4.400 829.240 345.600 829.280 ;
        RECT 4.400 827.880 346.000 829.240 ;
        RECT 3.950 826.560 346.000 827.880 ;
        RECT 4.400 825.200 346.000 826.560 ;
        RECT 4.400 825.160 345.600 825.200 ;
        RECT 3.950 823.840 345.600 825.160 ;
        RECT 4.400 823.800 345.600 823.840 ;
        RECT 4.400 822.440 346.000 823.800 ;
        RECT 3.950 821.120 346.000 822.440 ;
        RECT 4.400 819.760 346.000 821.120 ;
        RECT 4.400 819.720 345.600 819.760 ;
        RECT 3.950 818.400 345.600 819.720 ;
        RECT 4.400 818.360 345.600 818.400 ;
        RECT 4.400 817.000 346.000 818.360 ;
        RECT 3.950 815.680 346.000 817.000 ;
        RECT 4.400 814.320 346.000 815.680 ;
        RECT 4.400 814.280 345.600 814.320 ;
        RECT 3.950 812.960 345.600 814.280 ;
        RECT 4.400 812.920 345.600 812.960 ;
        RECT 4.400 811.560 346.000 812.920 ;
        RECT 3.950 810.240 346.000 811.560 ;
        RECT 4.400 808.880 346.000 810.240 ;
        RECT 4.400 808.840 345.600 808.880 ;
        RECT 3.950 807.520 345.600 808.840 ;
        RECT 4.400 807.480 345.600 807.520 ;
        RECT 4.400 806.120 346.000 807.480 ;
        RECT 3.950 804.800 346.000 806.120 ;
        RECT 4.400 803.440 346.000 804.800 ;
        RECT 4.400 803.400 345.600 803.440 ;
        RECT 3.950 802.080 345.600 803.400 ;
        RECT 4.400 802.040 345.600 802.080 ;
        RECT 4.400 800.680 346.000 802.040 ;
        RECT 3.950 799.360 346.000 800.680 ;
        RECT 4.400 798.000 346.000 799.360 ;
        RECT 4.400 797.960 345.600 798.000 ;
        RECT 3.950 796.640 345.600 797.960 ;
        RECT 4.400 796.600 345.600 796.640 ;
        RECT 4.400 795.240 346.000 796.600 ;
        RECT 3.950 793.920 346.000 795.240 ;
        RECT 4.400 792.560 346.000 793.920 ;
        RECT 4.400 792.520 345.600 792.560 ;
        RECT 3.950 791.200 345.600 792.520 ;
        RECT 4.400 791.160 345.600 791.200 ;
        RECT 4.400 789.800 346.000 791.160 ;
        RECT 3.950 788.480 346.000 789.800 ;
        RECT 4.400 787.120 346.000 788.480 ;
        RECT 4.400 787.080 345.600 787.120 ;
        RECT 3.950 785.760 345.600 787.080 ;
        RECT 4.400 785.720 345.600 785.760 ;
        RECT 4.400 784.360 346.000 785.720 ;
        RECT 3.950 783.040 346.000 784.360 ;
        RECT 4.400 781.680 346.000 783.040 ;
        RECT 4.400 781.640 345.600 781.680 ;
        RECT 3.950 780.320 345.600 781.640 ;
        RECT 4.400 780.280 345.600 780.320 ;
        RECT 4.400 778.920 346.000 780.280 ;
        RECT 3.950 777.600 346.000 778.920 ;
        RECT 4.400 776.240 346.000 777.600 ;
        RECT 4.400 776.200 345.600 776.240 ;
        RECT 3.950 774.880 345.600 776.200 ;
        RECT 4.400 774.840 345.600 774.880 ;
        RECT 4.400 773.480 346.000 774.840 ;
        RECT 3.950 772.160 346.000 773.480 ;
        RECT 4.400 770.800 346.000 772.160 ;
        RECT 4.400 770.760 345.600 770.800 ;
        RECT 3.950 769.440 345.600 770.760 ;
        RECT 4.400 769.400 345.600 769.440 ;
        RECT 4.400 768.040 346.000 769.400 ;
        RECT 3.950 766.720 346.000 768.040 ;
        RECT 4.400 765.360 346.000 766.720 ;
        RECT 4.400 765.320 345.600 765.360 ;
        RECT 3.950 764.000 345.600 765.320 ;
        RECT 4.400 763.960 345.600 764.000 ;
        RECT 4.400 762.600 346.000 763.960 ;
        RECT 3.950 761.280 346.000 762.600 ;
        RECT 4.400 759.920 346.000 761.280 ;
        RECT 4.400 759.880 345.600 759.920 ;
        RECT 3.950 758.560 345.600 759.880 ;
        RECT 4.400 758.520 345.600 758.560 ;
        RECT 4.400 757.160 346.000 758.520 ;
        RECT 3.950 755.840 346.000 757.160 ;
        RECT 4.400 754.480 346.000 755.840 ;
        RECT 4.400 754.440 345.600 754.480 ;
        RECT 3.950 753.120 345.600 754.440 ;
        RECT 4.400 753.080 345.600 753.120 ;
        RECT 4.400 751.720 346.000 753.080 ;
        RECT 3.950 750.400 346.000 751.720 ;
        RECT 4.400 749.040 346.000 750.400 ;
        RECT 4.400 749.000 345.600 749.040 ;
        RECT 3.950 747.680 345.600 749.000 ;
        RECT 4.400 747.640 345.600 747.680 ;
        RECT 4.400 746.280 346.000 747.640 ;
        RECT 3.950 744.960 346.000 746.280 ;
        RECT 4.400 743.600 346.000 744.960 ;
        RECT 4.400 743.560 345.600 743.600 ;
        RECT 3.950 742.240 345.600 743.560 ;
        RECT 4.400 742.200 345.600 742.240 ;
        RECT 4.400 740.840 346.000 742.200 ;
        RECT 3.950 739.520 346.000 740.840 ;
        RECT 4.400 738.160 346.000 739.520 ;
        RECT 4.400 738.120 345.600 738.160 ;
        RECT 3.950 736.800 345.600 738.120 ;
        RECT 4.400 736.760 345.600 736.800 ;
        RECT 4.400 735.400 346.000 736.760 ;
        RECT 3.950 734.080 346.000 735.400 ;
        RECT 4.400 732.720 346.000 734.080 ;
        RECT 4.400 732.680 345.600 732.720 ;
        RECT 3.950 731.360 345.600 732.680 ;
        RECT 4.400 731.320 345.600 731.360 ;
        RECT 4.400 729.960 346.000 731.320 ;
        RECT 3.950 728.640 346.000 729.960 ;
        RECT 4.400 727.280 346.000 728.640 ;
        RECT 4.400 727.240 345.600 727.280 ;
        RECT 3.950 725.920 345.600 727.240 ;
        RECT 4.400 725.880 345.600 725.920 ;
        RECT 4.400 724.520 346.000 725.880 ;
        RECT 3.950 723.200 346.000 724.520 ;
        RECT 4.400 721.840 346.000 723.200 ;
        RECT 4.400 721.800 345.600 721.840 ;
        RECT 3.950 720.480 345.600 721.800 ;
        RECT 4.400 720.440 345.600 720.480 ;
        RECT 4.400 719.080 346.000 720.440 ;
        RECT 3.950 717.760 346.000 719.080 ;
        RECT 4.400 716.400 346.000 717.760 ;
        RECT 4.400 716.360 345.600 716.400 ;
        RECT 3.950 715.040 345.600 716.360 ;
        RECT 4.400 715.000 345.600 715.040 ;
        RECT 4.400 713.640 346.000 715.000 ;
        RECT 3.950 712.320 346.000 713.640 ;
        RECT 4.400 710.960 346.000 712.320 ;
        RECT 4.400 710.920 345.600 710.960 ;
        RECT 3.950 709.600 345.600 710.920 ;
        RECT 4.400 709.560 345.600 709.600 ;
        RECT 4.400 708.200 346.000 709.560 ;
        RECT 3.950 706.880 346.000 708.200 ;
        RECT 4.400 705.520 346.000 706.880 ;
        RECT 4.400 705.480 345.600 705.520 ;
        RECT 3.950 704.160 345.600 705.480 ;
        RECT 4.400 704.120 345.600 704.160 ;
        RECT 4.400 702.760 346.000 704.120 ;
        RECT 3.950 701.440 346.000 702.760 ;
        RECT 4.400 700.080 346.000 701.440 ;
        RECT 4.400 700.040 345.600 700.080 ;
        RECT 3.950 698.720 345.600 700.040 ;
        RECT 4.400 698.680 345.600 698.720 ;
        RECT 4.400 697.320 346.000 698.680 ;
        RECT 3.950 696.000 346.000 697.320 ;
        RECT 4.400 694.640 346.000 696.000 ;
        RECT 4.400 694.600 345.600 694.640 ;
        RECT 3.950 693.280 345.600 694.600 ;
        RECT 4.400 693.240 345.600 693.280 ;
        RECT 4.400 691.880 346.000 693.240 ;
        RECT 3.950 690.560 346.000 691.880 ;
        RECT 4.400 689.200 346.000 690.560 ;
        RECT 4.400 689.160 345.600 689.200 ;
        RECT 3.950 687.840 345.600 689.160 ;
        RECT 4.400 687.800 345.600 687.840 ;
        RECT 4.400 686.440 346.000 687.800 ;
        RECT 3.950 685.120 346.000 686.440 ;
        RECT 4.400 683.760 346.000 685.120 ;
        RECT 4.400 683.720 345.600 683.760 ;
        RECT 3.950 682.400 345.600 683.720 ;
        RECT 4.400 682.360 345.600 682.400 ;
        RECT 4.400 681.000 346.000 682.360 ;
        RECT 3.950 679.680 346.000 681.000 ;
        RECT 4.400 678.320 346.000 679.680 ;
        RECT 4.400 678.280 345.600 678.320 ;
        RECT 3.950 676.960 345.600 678.280 ;
        RECT 4.400 676.920 345.600 676.960 ;
        RECT 4.400 675.560 346.000 676.920 ;
        RECT 3.950 674.240 346.000 675.560 ;
        RECT 4.400 672.880 346.000 674.240 ;
        RECT 4.400 672.840 345.600 672.880 ;
        RECT 3.950 671.520 345.600 672.840 ;
        RECT 4.400 671.480 345.600 671.520 ;
        RECT 4.400 670.120 346.000 671.480 ;
        RECT 3.950 668.800 346.000 670.120 ;
        RECT 4.400 667.440 346.000 668.800 ;
        RECT 4.400 667.400 345.600 667.440 ;
        RECT 3.950 666.080 345.600 667.400 ;
        RECT 4.400 666.040 345.600 666.080 ;
        RECT 4.400 664.680 346.000 666.040 ;
        RECT 3.950 663.360 346.000 664.680 ;
        RECT 4.400 662.000 346.000 663.360 ;
        RECT 4.400 661.960 345.600 662.000 ;
        RECT 3.950 660.640 345.600 661.960 ;
        RECT 4.400 660.600 345.600 660.640 ;
        RECT 4.400 659.240 346.000 660.600 ;
        RECT 3.950 657.920 346.000 659.240 ;
        RECT 4.400 656.560 346.000 657.920 ;
        RECT 4.400 656.520 345.600 656.560 ;
        RECT 3.950 655.200 345.600 656.520 ;
        RECT 4.400 655.160 345.600 655.200 ;
        RECT 4.400 653.800 346.000 655.160 ;
        RECT 3.950 652.480 346.000 653.800 ;
        RECT 4.400 651.120 346.000 652.480 ;
        RECT 4.400 651.080 345.600 651.120 ;
        RECT 3.950 649.760 345.600 651.080 ;
        RECT 4.400 649.720 345.600 649.760 ;
        RECT 4.400 648.360 346.000 649.720 ;
        RECT 3.950 647.040 346.000 648.360 ;
        RECT 4.400 645.680 346.000 647.040 ;
        RECT 4.400 645.640 345.600 645.680 ;
        RECT 3.950 644.320 345.600 645.640 ;
        RECT 4.400 644.280 345.600 644.320 ;
        RECT 4.400 642.920 346.000 644.280 ;
        RECT 3.950 641.600 346.000 642.920 ;
        RECT 4.400 640.240 346.000 641.600 ;
        RECT 4.400 640.200 345.600 640.240 ;
        RECT 3.950 638.880 345.600 640.200 ;
        RECT 4.400 638.840 345.600 638.880 ;
        RECT 4.400 637.480 346.000 638.840 ;
        RECT 3.950 636.160 346.000 637.480 ;
        RECT 4.400 634.800 346.000 636.160 ;
        RECT 4.400 634.760 345.600 634.800 ;
        RECT 3.950 633.440 345.600 634.760 ;
        RECT 4.400 633.400 345.600 633.440 ;
        RECT 4.400 632.040 346.000 633.400 ;
        RECT 3.950 630.720 346.000 632.040 ;
        RECT 4.400 629.360 346.000 630.720 ;
        RECT 4.400 629.320 345.600 629.360 ;
        RECT 3.950 628.000 345.600 629.320 ;
        RECT 4.400 627.960 345.600 628.000 ;
        RECT 4.400 626.600 346.000 627.960 ;
        RECT 3.950 625.280 346.000 626.600 ;
        RECT 4.400 623.920 346.000 625.280 ;
        RECT 4.400 623.880 345.600 623.920 ;
        RECT 3.950 622.560 345.600 623.880 ;
        RECT 4.400 622.520 345.600 622.560 ;
        RECT 4.400 621.160 346.000 622.520 ;
        RECT 3.950 619.840 346.000 621.160 ;
        RECT 4.400 618.480 346.000 619.840 ;
        RECT 4.400 618.440 345.600 618.480 ;
        RECT 3.950 617.120 345.600 618.440 ;
        RECT 4.400 617.080 345.600 617.120 ;
        RECT 4.400 615.720 346.000 617.080 ;
        RECT 3.950 614.400 346.000 615.720 ;
        RECT 4.400 613.040 346.000 614.400 ;
        RECT 4.400 613.000 345.600 613.040 ;
        RECT 3.950 611.680 345.600 613.000 ;
        RECT 4.400 611.640 345.600 611.680 ;
        RECT 4.400 610.280 346.000 611.640 ;
        RECT 3.950 608.960 346.000 610.280 ;
        RECT 4.400 607.600 346.000 608.960 ;
        RECT 4.400 607.560 345.600 607.600 ;
        RECT 3.950 606.240 345.600 607.560 ;
        RECT 4.400 606.200 345.600 606.240 ;
        RECT 4.400 604.840 346.000 606.200 ;
        RECT 3.950 603.520 346.000 604.840 ;
        RECT 4.400 602.160 346.000 603.520 ;
        RECT 4.400 602.120 345.600 602.160 ;
        RECT 3.950 600.800 345.600 602.120 ;
        RECT 4.400 600.760 345.600 600.800 ;
        RECT 4.400 599.400 346.000 600.760 ;
        RECT 3.950 598.080 346.000 599.400 ;
        RECT 4.400 596.720 346.000 598.080 ;
        RECT 4.400 596.680 345.600 596.720 ;
        RECT 3.950 595.360 345.600 596.680 ;
        RECT 4.400 595.320 345.600 595.360 ;
        RECT 4.400 593.960 346.000 595.320 ;
        RECT 3.950 592.640 346.000 593.960 ;
        RECT 4.400 591.280 346.000 592.640 ;
        RECT 4.400 591.240 345.600 591.280 ;
        RECT 3.950 589.920 345.600 591.240 ;
        RECT 4.400 589.880 345.600 589.920 ;
        RECT 4.400 588.520 346.000 589.880 ;
        RECT 3.950 587.200 346.000 588.520 ;
        RECT 4.400 585.840 346.000 587.200 ;
        RECT 4.400 585.800 345.600 585.840 ;
        RECT 3.950 584.480 345.600 585.800 ;
        RECT 4.400 584.440 345.600 584.480 ;
        RECT 4.400 583.080 346.000 584.440 ;
        RECT 3.950 581.760 346.000 583.080 ;
        RECT 4.400 580.400 346.000 581.760 ;
        RECT 4.400 580.360 345.600 580.400 ;
        RECT 3.950 579.040 345.600 580.360 ;
        RECT 4.400 579.000 345.600 579.040 ;
        RECT 4.400 577.640 346.000 579.000 ;
        RECT 3.950 576.320 346.000 577.640 ;
        RECT 4.400 574.960 346.000 576.320 ;
        RECT 4.400 574.920 345.600 574.960 ;
        RECT 3.950 573.600 345.600 574.920 ;
        RECT 4.400 573.560 345.600 573.600 ;
        RECT 4.400 572.200 346.000 573.560 ;
        RECT 3.950 570.880 346.000 572.200 ;
        RECT 4.400 569.520 346.000 570.880 ;
        RECT 4.400 569.480 345.600 569.520 ;
        RECT 3.950 568.160 345.600 569.480 ;
        RECT 4.400 568.120 345.600 568.160 ;
        RECT 4.400 566.760 346.000 568.120 ;
        RECT 3.950 565.440 346.000 566.760 ;
        RECT 4.400 564.080 346.000 565.440 ;
        RECT 4.400 564.040 345.600 564.080 ;
        RECT 3.950 562.720 345.600 564.040 ;
        RECT 4.400 562.680 345.600 562.720 ;
        RECT 4.400 561.320 346.000 562.680 ;
        RECT 3.950 560.000 346.000 561.320 ;
        RECT 4.400 558.640 346.000 560.000 ;
        RECT 4.400 558.600 345.600 558.640 ;
        RECT 3.950 557.280 345.600 558.600 ;
        RECT 4.400 557.240 345.600 557.280 ;
        RECT 4.400 555.880 346.000 557.240 ;
        RECT 3.950 554.560 346.000 555.880 ;
        RECT 4.400 553.200 346.000 554.560 ;
        RECT 4.400 553.160 345.600 553.200 ;
        RECT 3.950 551.840 345.600 553.160 ;
        RECT 4.400 551.800 345.600 551.840 ;
        RECT 4.400 550.440 346.000 551.800 ;
        RECT 3.950 549.120 346.000 550.440 ;
        RECT 4.400 547.760 346.000 549.120 ;
        RECT 4.400 547.720 345.600 547.760 ;
        RECT 3.950 546.400 345.600 547.720 ;
        RECT 4.400 546.360 345.600 546.400 ;
        RECT 4.400 545.000 346.000 546.360 ;
        RECT 3.950 543.680 346.000 545.000 ;
        RECT 4.400 542.320 346.000 543.680 ;
        RECT 4.400 542.280 345.600 542.320 ;
        RECT 3.950 540.960 345.600 542.280 ;
        RECT 4.400 540.920 345.600 540.960 ;
        RECT 4.400 539.560 346.000 540.920 ;
        RECT 3.950 538.240 346.000 539.560 ;
        RECT 4.400 536.880 346.000 538.240 ;
        RECT 4.400 536.840 345.600 536.880 ;
        RECT 3.950 535.520 345.600 536.840 ;
        RECT 4.400 535.480 345.600 535.520 ;
        RECT 4.400 534.120 346.000 535.480 ;
        RECT 3.950 532.800 346.000 534.120 ;
        RECT 4.400 531.440 346.000 532.800 ;
        RECT 4.400 531.400 345.600 531.440 ;
        RECT 3.950 530.080 345.600 531.400 ;
        RECT 4.400 530.040 345.600 530.080 ;
        RECT 4.400 528.680 346.000 530.040 ;
        RECT 3.950 527.360 346.000 528.680 ;
        RECT 4.400 526.000 346.000 527.360 ;
        RECT 4.400 525.960 345.600 526.000 ;
        RECT 3.950 524.640 345.600 525.960 ;
        RECT 4.400 524.600 345.600 524.640 ;
        RECT 4.400 523.240 346.000 524.600 ;
        RECT 3.950 521.920 346.000 523.240 ;
        RECT 4.400 520.560 346.000 521.920 ;
        RECT 4.400 520.520 345.600 520.560 ;
        RECT 3.950 519.200 345.600 520.520 ;
        RECT 4.400 519.160 345.600 519.200 ;
        RECT 4.400 517.800 346.000 519.160 ;
        RECT 3.950 516.480 346.000 517.800 ;
        RECT 4.400 515.120 346.000 516.480 ;
        RECT 4.400 515.080 345.600 515.120 ;
        RECT 3.950 513.760 345.600 515.080 ;
        RECT 4.400 513.720 345.600 513.760 ;
        RECT 4.400 512.360 346.000 513.720 ;
        RECT 3.950 511.040 346.000 512.360 ;
        RECT 4.400 509.680 346.000 511.040 ;
        RECT 4.400 509.640 345.600 509.680 ;
        RECT 3.950 508.320 345.600 509.640 ;
        RECT 4.400 508.280 345.600 508.320 ;
        RECT 4.400 506.920 346.000 508.280 ;
        RECT 3.950 505.600 346.000 506.920 ;
        RECT 4.400 504.240 346.000 505.600 ;
        RECT 4.400 504.200 345.600 504.240 ;
        RECT 3.950 502.880 345.600 504.200 ;
        RECT 4.400 502.840 345.600 502.880 ;
        RECT 4.400 501.480 346.000 502.840 ;
        RECT 3.950 500.160 346.000 501.480 ;
        RECT 4.400 498.800 346.000 500.160 ;
        RECT 4.400 498.760 345.600 498.800 ;
        RECT 3.950 497.440 345.600 498.760 ;
        RECT 4.400 497.400 345.600 497.440 ;
        RECT 4.400 496.040 346.000 497.400 ;
        RECT 3.950 494.720 346.000 496.040 ;
        RECT 4.400 493.360 346.000 494.720 ;
        RECT 4.400 493.320 345.600 493.360 ;
        RECT 3.950 492.000 345.600 493.320 ;
        RECT 4.400 491.960 345.600 492.000 ;
        RECT 4.400 490.600 346.000 491.960 ;
        RECT 3.950 489.280 346.000 490.600 ;
        RECT 4.400 487.920 346.000 489.280 ;
        RECT 4.400 487.880 345.600 487.920 ;
        RECT 3.950 486.560 345.600 487.880 ;
        RECT 4.400 486.520 345.600 486.560 ;
        RECT 4.400 485.160 346.000 486.520 ;
        RECT 3.950 483.840 346.000 485.160 ;
        RECT 4.400 482.480 346.000 483.840 ;
        RECT 4.400 482.440 345.600 482.480 ;
        RECT 3.950 481.120 345.600 482.440 ;
        RECT 4.400 481.080 345.600 481.120 ;
        RECT 4.400 479.720 346.000 481.080 ;
        RECT 3.950 478.400 346.000 479.720 ;
        RECT 4.400 477.040 346.000 478.400 ;
        RECT 4.400 477.000 345.600 477.040 ;
        RECT 3.950 475.680 345.600 477.000 ;
        RECT 4.400 475.640 345.600 475.680 ;
        RECT 4.400 474.280 346.000 475.640 ;
        RECT 3.950 472.960 346.000 474.280 ;
        RECT 4.400 471.600 346.000 472.960 ;
        RECT 4.400 471.560 345.600 471.600 ;
        RECT 3.950 470.240 345.600 471.560 ;
        RECT 4.400 470.200 345.600 470.240 ;
        RECT 4.400 468.840 346.000 470.200 ;
        RECT 3.950 467.520 346.000 468.840 ;
        RECT 4.400 466.160 346.000 467.520 ;
        RECT 4.400 466.120 345.600 466.160 ;
        RECT 3.950 464.800 345.600 466.120 ;
        RECT 4.400 464.760 345.600 464.800 ;
        RECT 4.400 463.400 346.000 464.760 ;
        RECT 3.950 462.080 346.000 463.400 ;
        RECT 4.400 460.720 346.000 462.080 ;
        RECT 4.400 460.680 345.600 460.720 ;
        RECT 3.950 459.360 345.600 460.680 ;
        RECT 4.400 459.320 345.600 459.360 ;
        RECT 4.400 457.960 346.000 459.320 ;
        RECT 3.950 456.640 346.000 457.960 ;
        RECT 4.400 455.280 346.000 456.640 ;
        RECT 4.400 455.240 345.600 455.280 ;
        RECT 3.950 453.920 345.600 455.240 ;
        RECT 4.400 453.880 345.600 453.920 ;
        RECT 4.400 452.520 346.000 453.880 ;
        RECT 3.950 451.200 346.000 452.520 ;
        RECT 4.400 449.840 346.000 451.200 ;
        RECT 4.400 449.800 345.600 449.840 ;
        RECT 3.950 448.480 345.600 449.800 ;
        RECT 4.400 448.440 345.600 448.480 ;
        RECT 4.400 447.080 346.000 448.440 ;
        RECT 3.950 445.760 346.000 447.080 ;
        RECT 4.400 444.400 346.000 445.760 ;
        RECT 4.400 444.360 345.600 444.400 ;
        RECT 3.950 443.040 345.600 444.360 ;
        RECT 4.400 443.000 345.600 443.040 ;
        RECT 4.400 441.640 346.000 443.000 ;
        RECT 3.950 440.320 346.000 441.640 ;
        RECT 4.400 438.960 346.000 440.320 ;
        RECT 4.400 438.920 345.600 438.960 ;
        RECT 3.950 437.600 345.600 438.920 ;
        RECT 4.400 437.560 345.600 437.600 ;
        RECT 4.400 436.200 346.000 437.560 ;
        RECT 3.950 434.880 346.000 436.200 ;
        RECT 4.400 433.520 346.000 434.880 ;
        RECT 4.400 433.480 345.600 433.520 ;
        RECT 3.950 432.160 345.600 433.480 ;
        RECT 4.400 432.120 345.600 432.160 ;
        RECT 4.400 430.760 346.000 432.120 ;
        RECT 3.950 429.440 346.000 430.760 ;
        RECT 4.400 428.080 346.000 429.440 ;
        RECT 4.400 428.040 345.600 428.080 ;
        RECT 3.950 426.720 345.600 428.040 ;
        RECT 4.400 426.680 345.600 426.720 ;
        RECT 4.400 425.320 346.000 426.680 ;
        RECT 3.950 424.000 346.000 425.320 ;
        RECT 4.400 422.640 346.000 424.000 ;
        RECT 4.400 422.600 345.600 422.640 ;
        RECT 3.950 421.280 345.600 422.600 ;
        RECT 4.400 421.240 345.600 421.280 ;
        RECT 4.400 419.880 346.000 421.240 ;
        RECT 3.950 418.560 346.000 419.880 ;
        RECT 4.400 417.200 346.000 418.560 ;
        RECT 4.400 417.160 345.600 417.200 ;
        RECT 3.950 415.840 345.600 417.160 ;
        RECT 4.400 415.800 345.600 415.840 ;
        RECT 4.400 414.440 346.000 415.800 ;
        RECT 3.950 413.120 346.000 414.440 ;
        RECT 4.400 411.760 346.000 413.120 ;
        RECT 4.400 411.720 345.600 411.760 ;
        RECT 3.950 410.400 345.600 411.720 ;
        RECT 4.400 410.360 345.600 410.400 ;
        RECT 4.400 409.000 346.000 410.360 ;
        RECT 3.950 407.680 346.000 409.000 ;
        RECT 4.400 406.320 346.000 407.680 ;
        RECT 4.400 406.280 345.600 406.320 ;
        RECT 3.950 404.960 345.600 406.280 ;
        RECT 4.400 404.920 345.600 404.960 ;
        RECT 4.400 403.560 346.000 404.920 ;
        RECT 3.950 402.240 346.000 403.560 ;
        RECT 4.400 400.880 346.000 402.240 ;
        RECT 4.400 400.840 345.600 400.880 ;
        RECT 3.950 399.520 345.600 400.840 ;
        RECT 4.400 399.480 345.600 399.520 ;
        RECT 4.400 398.120 346.000 399.480 ;
        RECT 3.950 396.800 346.000 398.120 ;
        RECT 4.400 395.440 346.000 396.800 ;
        RECT 4.400 395.400 345.600 395.440 ;
        RECT 3.950 394.080 345.600 395.400 ;
        RECT 4.400 394.040 345.600 394.080 ;
        RECT 4.400 392.680 346.000 394.040 ;
        RECT 3.950 391.360 346.000 392.680 ;
        RECT 4.400 390.000 346.000 391.360 ;
        RECT 4.400 389.960 345.600 390.000 ;
        RECT 3.950 388.640 345.600 389.960 ;
        RECT 4.400 388.600 345.600 388.640 ;
        RECT 4.400 387.240 346.000 388.600 ;
        RECT 3.950 385.920 346.000 387.240 ;
        RECT 4.400 384.560 346.000 385.920 ;
        RECT 4.400 384.520 345.600 384.560 ;
        RECT 3.950 383.200 345.600 384.520 ;
        RECT 4.400 383.160 345.600 383.200 ;
        RECT 4.400 381.800 346.000 383.160 ;
        RECT 3.950 380.480 346.000 381.800 ;
        RECT 4.400 379.120 346.000 380.480 ;
        RECT 4.400 379.080 345.600 379.120 ;
        RECT 3.950 377.760 345.600 379.080 ;
        RECT 4.400 377.720 345.600 377.760 ;
        RECT 4.400 376.360 346.000 377.720 ;
        RECT 3.950 375.040 346.000 376.360 ;
        RECT 4.400 373.680 346.000 375.040 ;
        RECT 4.400 373.640 345.600 373.680 ;
        RECT 3.950 372.320 345.600 373.640 ;
        RECT 4.400 372.280 345.600 372.320 ;
        RECT 4.400 370.920 346.000 372.280 ;
        RECT 3.950 369.600 346.000 370.920 ;
        RECT 4.400 368.240 346.000 369.600 ;
        RECT 4.400 368.200 345.600 368.240 ;
        RECT 3.950 366.880 345.600 368.200 ;
        RECT 4.400 366.840 345.600 366.880 ;
        RECT 4.400 365.480 346.000 366.840 ;
        RECT 3.950 364.160 346.000 365.480 ;
        RECT 4.400 362.800 346.000 364.160 ;
        RECT 4.400 362.760 345.600 362.800 ;
        RECT 3.950 361.440 345.600 362.760 ;
        RECT 4.400 361.400 345.600 361.440 ;
        RECT 4.400 360.040 346.000 361.400 ;
        RECT 3.950 358.720 346.000 360.040 ;
        RECT 4.400 357.360 346.000 358.720 ;
        RECT 4.400 357.320 345.600 357.360 ;
        RECT 3.950 356.000 345.600 357.320 ;
        RECT 4.400 355.960 345.600 356.000 ;
        RECT 4.400 354.600 346.000 355.960 ;
        RECT 3.950 353.280 346.000 354.600 ;
        RECT 4.400 351.920 346.000 353.280 ;
        RECT 4.400 351.880 345.600 351.920 ;
        RECT 3.950 350.560 345.600 351.880 ;
        RECT 4.400 350.520 345.600 350.560 ;
        RECT 4.400 349.160 346.000 350.520 ;
        RECT 3.950 347.840 346.000 349.160 ;
        RECT 4.400 346.480 346.000 347.840 ;
        RECT 4.400 346.440 345.600 346.480 ;
        RECT 3.950 345.120 345.600 346.440 ;
        RECT 4.400 345.080 345.600 345.120 ;
        RECT 4.400 343.720 346.000 345.080 ;
        RECT 3.950 342.400 346.000 343.720 ;
        RECT 4.400 341.040 346.000 342.400 ;
        RECT 4.400 341.000 345.600 341.040 ;
        RECT 3.950 339.680 345.600 341.000 ;
        RECT 4.400 339.640 345.600 339.680 ;
        RECT 4.400 338.280 346.000 339.640 ;
        RECT 3.950 336.960 346.000 338.280 ;
        RECT 4.400 335.600 346.000 336.960 ;
        RECT 4.400 335.560 345.600 335.600 ;
        RECT 3.950 334.240 345.600 335.560 ;
        RECT 4.400 334.200 345.600 334.240 ;
        RECT 4.400 332.840 346.000 334.200 ;
        RECT 3.950 331.520 346.000 332.840 ;
        RECT 4.400 330.160 346.000 331.520 ;
        RECT 4.400 330.120 345.600 330.160 ;
        RECT 3.950 328.800 345.600 330.120 ;
        RECT 4.400 328.760 345.600 328.800 ;
        RECT 4.400 327.400 346.000 328.760 ;
        RECT 3.950 326.080 346.000 327.400 ;
        RECT 4.400 324.720 346.000 326.080 ;
        RECT 4.400 324.680 345.600 324.720 ;
        RECT 3.950 323.360 345.600 324.680 ;
        RECT 4.400 323.320 345.600 323.360 ;
        RECT 4.400 321.960 346.000 323.320 ;
        RECT 3.950 320.640 346.000 321.960 ;
        RECT 4.400 319.280 346.000 320.640 ;
        RECT 4.400 319.240 345.600 319.280 ;
        RECT 3.950 317.920 345.600 319.240 ;
        RECT 4.400 317.880 345.600 317.920 ;
        RECT 4.400 316.520 346.000 317.880 ;
        RECT 3.950 315.200 346.000 316.520 ;
        RECT 4.400 313.840 346.000 315.200 ;
        RECT 4.400 313.800 345.600 313.840 ;
        RECT 3.950 312.480 345.600 313.800 ;
        RECT 4.400 312.440 345.600 312.480 ;
        RECT 4.400 311.080 346.000 312.440 ;
        RECT 3.950 309.760 346.000 311.080 ;
        RECT 4.400 308.400 346.000 309.760 ;
        RECT 4.400 308.360 345.600 308.400 ;
        RECT 3.950 307.040 345.600 308.360 ;
        RECT 4.400 307.000 345.600 307.040 ;
        RECT 4.400 305.640 346.000 307.000 ;
        RECT 3.950 304.320 346.000 305.640 ;
        RECT 4.400 302.960 346.000 304.320 ;
        RECT 4.400 302.920 345.600 302.960 ;
        RECT 3.950 301.600 345.600 302.920 ;
        RECT 4.400 301.560 345.600 301.600 ;
        RECT 4.400 300.200 346.000 301.560 ;
        RECT 3.950 298.880 346.000 300.200 ;
        RECT 4.400 297.520 346.000 298.880 ;
        RECT 4.400 297.480 345.600 297.520 ;
        RECT 3.950 296.160 345.600 297.480 ;
        RECT 4.400 296.120 345.600 296.160 ;
        RECT 4.400 294.760 346.000 296.120 ;
        RECT 3.950 293.440 346.000 294.760 ;
        RECT 4.400 292.080 346.000 293.440 ;
        RECT 4.400 292.040 345.600 292.080 ;
        RECT 3.950 290.720 345.600 292.040 ;
        RECT 4.400 290.680 345.600 290.720 ;
        RECT 4.400 289.320 346.000 290.680 ;
        RECT 3.950 288.000 346.000 289.320 ;
        RECT 4.400 286.640 346.000 288.000 ;
        RECT 4.400 286.600 345.600 286.640 ;
        RECT 3.950 285.280 345.600 286.600 ;
        RECT 4.400 285.240 345.600 285.280 ;
        RECT 4.400 283.880 346.000 285.240 ;
        RECT 3.950 282.560 346.000 283.880 ;
        RECT 4.400 281.200 346.000 282.560 ;
        RECT 4.400 281.160 345.600 281.200 ;
        RECT 3.950 279.840 345.600 281.160 ;
        RECT 4.400 279.800 345.600 279.840 ;
        RECT 4.400 278.440 346.000 279.800 ;
        RECT 3.950 277.120 346.000 278.440 ;
        RECT 4.400 275.760 346.000 277.120 ;
        RECT 4.400 275.720 345.600 275.760 ;
        RECT 3.950 274.400 345.600 275.720 ;
        RECT 4.400 274.360 345.600 274.400 ;
        RECT 4.400 273.000 346.000 274.360 ;
        RECT 3.950 271.680 346.000 273.000 ;
        RECT 4.400 270.320 346.000 271.680 ;
        RECT 4.400 270.280 345.600 270.320 ;
        RECT 3.950 268.960 345.600 270.280 ;
        RECT 4.400 268.920 345.600 268.960 ;
        RECT 4.400 267.560 346.000 268.920 ;
        RECT 3.950 266.240 346.000 267.560 ;
        RECT 4.400 264.880 346.000 266.240 ;
        RECT 4.400 264.840 345.600 264.880 ;
        RECT 3.950 263.520 345.600 264.840 ;
        RECT 4.400 263.480 345.600 263.520 ;
        RECT 4.400 262.120 346.000 263.480 ;
        RECT 3.950 260.800 346.000 262.120 ;
        RECT 4.400 259.440 346.000 260.800 ;
        RECT 4.400 259.400 345.600 259.440 ;
        RECT 3.950 258.080 345.600 259.400 ;
        RECT 4.400 258.040 345.600 258.080 ;
        RECT 4.400 256.680 346.000 258.040 ;
        RECT 3.950 255.360 346.000 256.680 ;
        RECT 4.400 254.000 346.000 255.360 ;
        RECT 4.400 253.960 345.600 254.000 ;
        RECT 3.950 252.640 345.600 253.960 ;
        RECT 4.400 252.600 345.600 252.640 ;
        RECT 4.400 251.240 346.000 252.600 ;
        RECT 3.950 249.920 346.000 251.240 ;
        RECT 4.400 248.560 346.000 249.920 ;
        RECT 4.400 248.520 345.600 248.560 ;
        RECT 3.950 247.200 345.600 248.520 ;
        RECT 4.400 247.160 345.600 247.200 ;
        RECT 4.400 245.800 346.000 247.160 ;
        RECT 3.950 244.480 346.000 245.800 ;
        RECT 4.400 243.120 346.000 244.480 ;
        RECT 4.400 243.080 345.600 243.120 ;
        RECT 3.950 241.760 345.600 243.080 ;
        RECT 4.400 241.720 345.600 241.760 ;
        RECT 4.400 240.360 346.000 241.720 ;
        RECT 3.950 239.040 346.000 240.360 ;
        RECT 4.400 237.680 346.000 239.040 ;
        RECT 4.400 237.640 345.600 237.680 ;
        RECT 3.950 236.320 345.600 237.640 ;
        RECT 4.400 236.280 345.600 236.320 ;
        RECT 4.400 234.920 346.000 236.280 ;
        RECT 3.950 233.600 346.000 234.920 ;
        RECT 4.400 232.240 346.000 233.600 ;
        RECT 4.400 232.200 345.600 232.240 ;
        RECT 3.950 230.880 345.600 232.200 ;
        RECT 4.400 230.840 345.600 230.880 ;
        RECT 4.400 229.480 346.000 230.840 ;
        RECT 3.950 228.160 346.000 229.480 ;
        RECT 4.400 226.800 346.000 228.160 ;
        RECT 4.400 226.760 345.600 226.800 ;
        RECT 3.950 225.440 345.600 226.760 ;
        RECT 4.400 225.400 345.600 225.440 ;
        RECT 4.400 224.040 346.000 225.400 ;
        RECT 3.950 222.720 346.000 224.040 ;
        RECT 4.400 221.360 346.000 222.720 ;
        RECT 4.400 221.320 345.600 221.360 ;
        RECT 3.950 220.000 345.600 221.320 ;
        RECT 4.400 219.960 345.600 220.000 ;
        RECT 4.400 218.600 346.000 219.960 ;
        RECT 3.950 217.280 346.000 218.600 ;
        RECT 4.400 215.920 346.000 217.280 ;
        RECT 4.400 215.880 345.600 215.920 ;
        RECT 3.950 214.560 345.600 215.880 ;
        RECT 4.400 214.520 345.600 214.560 ;
        RECT 4.400 213.160 346.000 214.520 ;
        RECT 3.950 211.840 346.000 213.160 ;
        RECT 4.400 210.480 346.000 211.840 ;
        RECT 4.400 210.440 345.600 210.480 ;
        RECT 3.950 209.120 345.600 210.440 ;
        RECT 4.400 209.080 345.600 209.120 ;
        RECT 4.400 207.720 346.000 209.080 ;
        RECT 3.950 206.400 346.000 207.720 ;
        RECT 4.400 205.040 346.000 206.400 ;
        RECT 4.400 205.000 345.600 205.040 ;
        RECT 3.950 203.680 345.600 205.000 ;
        RECT 4.400 203.640 345.600 203.680 ;
        RECT 4.400 202.280 346.000 203.640 ;
        RECT 3.950 200.960 346.000 202.280 ;
        RECT 4.400 199.600 346.000 200.960 ;
        RECT 4.400 199.560 345.600 199.600 ;
        RECT 3.950 198.240 345.600 199.560 ;
        RECT 4.400 198.200 345.600 198.240 ;
        RECT 4.400 196.840 346.000 198.200 ;
        RECT 3.950 195.520 346.000 196.840 ;
        RECT 4.400 194.160 346.000 195.520 ;
        RECT 4.400 194.120 345.600 194.160 ;
        RECT 3.950 192.800 345.600 194.120 ;
        RECT 4.400 192.760 345.600 192.800 ;
        RECT 4.400 191.400 346.000 192.760 ;
        RECT 3.950 190.080 346.000 191.400 ;
        RECT 4.400 188.720 346.000 190.080 ;
        RECT 4.400 188.680 345.600 188.720 ;
        RECT 3.950 187.360 345.600 188.680 ;
        RECT 4.400 187.320 345.600 187.360 ;
        RECT 4.400 185.960 346.000 187.320 ;
        RECT 3.950 184.640 346.000 185.960 ;
        RECT 4.400 183.280 346.000 184.640 ;
        RECT 4.400 183.240 345.600 183.280 ;
        RECT 3.950 181.920 345.600 183.240 ;
        RECT 4.400 181.880 345.600 181.920 ;
        RECT 4.400 180.520 346.000 181.880 ;
        RECT 3.950 179.200 346.000 180.520 ;
        RECT 4.400 177.840 346.000 179.200 ;
        RECT 4.400 177.800 345.600 177.840 ;
        RECT 3.950 176.480 345.600 177.800 ;
        RECT 4.400 176.440 345.600 176.480 ;
        RECT 4.400 175.080 346.000 176.440 ;
        RECT 3.950 173.760 346.000 175.080 ;
        RECT 4.400 172.400 346.000 173.760 ;
        RECT 4.400 172.360 345.600 172.400 ;
        RECT 3.950 171.040 345.600 172.360 ;
        RECT 4.400 171.000 345.600 171.040 ;
        RECT 4.400 169.640 346.000 171.000 ;
        RECT 3.950 168.320 346.000 169.640 ;
        RECT 4.400 166.960 346.000 168.320 ;
        RECT 4.400 166.920 345.600 166.960 ;
        RECT 3.950 165.600 345.600 166.920 ;
        RECT 4.400 165.560 345.600 165.600 ;
        RECT 4.400 164.200 346.000 165.560 ;
        RECT 3.950 162.880 346.000 164.200 ;
        RECT 4.400 161.520 346.000 162.880 ;
        RECT 4.400 161.480 345.600 161.520 ;
        RECT 3.950 160.160 345.600 161.480 ;
        RECT 4.400 160.120 345.600 160.160 ;
        RECT 4.400 158.760 346.000 160.120 ;
        RECT 3.950 157.440 346.000 158.760 ;
        RECT 4.400 156.080 346.000 157.440 ;
        RECT 4.400 156.040 345.600 156.080 ;
        RECT 3.950 154.720 345.600 156.040 ;
        RECT 4.400 154.680 345.600 154.720 ;
        RECT 4.400 153.320 346.000 154.680 ;
        RECT 3.950 152.000 346.000 153.320 ;
        RECT 4.400 150.640 346.000 152.000 ;
        RECT 4.400 150.600 345.600 150.640 ;
        RECT 3.950 149.280 345.600 150.600 ;
        RECT 4.400 149.240 345.600 149.280 ;
        RECT 4.400 147.880 346.000 149.240 ;
        RECT 3.950 146.560 346.000 147.880 ;
        RECT 4.400 145.200 346.000 146.560 ;
        RECT 4.400 145.160 345.600 145.200 ;
        RECT 3.950 143.840 345.600 145.160 ;
        RECT 4.400 143.800 345.600 143.840 ;
        RECT 4.400 142.440 346.000 143.800 ;
        RECT 3.950 141.120 346.000 142.440 ;
        RECT 4.400 139.760 346.000 141.120 ;
        RECT 4.400 139.720 345.600 139.760 ;
        RECT 3.950 138.400 345.600 139.720 ;
        RECT 4.400 138.360 345.600 138.400 ;
        RECT 4.400 137.000 346.000 138.360 ;
        RECT 3.950 135.680 346.000 137.000 ;
        RECT 4.400 134.320 346.000 135.680 ;
        RECT 4.400 134.280 345.600 134.320 ;
        RECT 3.950 132.960 345.600 134.280 ;
        RECT 4.400 132.920 345.600 132.960 ;
        RECT 4.400 131.560 346.000 132.920 ;
        RECT 3.950 130.240 346.000 131.560 ;
        RECT 4.400 128.880 346.000 130.240 ;
        RECT 4.400 128.840 345.600 128.880 ;
        RECT 3.950 127.520 345.600 128.840 ;
        RECT 4.400 127.480 345.600 127.520 ;
        RECT 4.400 126.120 346.000 127.480 ;
        RECT 3.950 124.800 346.000 126.120 ;
        RECT 4.400 123.440 346.000 124.800 ;
        RECT 4.400 123.400 345.600 123.440 ;
        RECT 3.950 122.080 345.600 123.400 ;
        RECT 4.400 122.040 345.600 122.080 ;
        RECT 4.400 120.680 346.000 122.040 ;
        RECT 3.950 119.360 346.000 120.680 ;
        RECT 4.400 118.000 346.000 119.360 ;
        RECT 4.400 117.960 345.600 118.000 ;
        RECT 3.950 116.640 345.600 117.960 ;
        RECT 4.400 116.600 345.600 116.640 ;
        RECT 4.400 115.240 346.000 116.600 ;
        RECT 3.950 113.920 346.000 115.240 ;
        RECT 4.400 112.560 346.000 113.920 ;
        RECT 4.400 112.520 345.600 112.560 ;
        RECT 3.950 111.200 345.600 112.520 ;
        RECT 4.400 111.160 345.600 111.200 ;
        RECT 4.400 109.800 346.000 111.160 ;
        RECT 3.950 108.480 346.000 109.800 ;
        RECT 4.400 107.120 346.000 108.480 ;
        RECT 4.400 107.080 345.600 107.120 ;
        RECT 3.950 105.760 345.600 107.080 ;
        RECT 4.400 105.720 345.600 105.760 ;
        RECT 4.400 104.360 346.000 105.720 ;
        RECT 3.950 103.040 346.000 104.360 ;
        RECT 4.400 101.680 346.000 103.040 ;
        RECT 4.400 101.640 345.600 101.680 ;
        RECT 3.950 100.320 345.600 101.640 ;
        RECT 4.400 100.280 345.600 100.320 ;
        RECT 4.400 98.920 346.000 100.280 ;
        RECT 3.950 97.600 346.000 98.920 ;
        RECT 4.400 96.240 346.000 97.600 ;
        RECT 4.400 96.200 345.600 96.240 ;
        RECT 3.950 94.880 345.600 96.200 ;
        RECT 4.400 94.840 345.600 94.880 ;
        RECT 4.400 93.480 346.000 94.840 ;
        RECT 3.950 92.160 346.000 93.480 ;
        RECT 4.400 90.800 346.000 92.160 ;
        RECT 4.400 90.760 345.600 90.800 ;
        RECT 3.950 89.440 345.600 90.760 ;
        RECT 4.400 89.400 345.600 89.440 ;
        RECT 4.400 88.040 346.000 89.400 ;
        RECT 3.950 86.720 346.000 88.040 ;
        RECT 4.400 85.360 346.000 86.720 ;
        RECT 4.400 85.320 345.600 85.360 ;
        RECT 3.950 84.000 345.600 85.320 ;
        RECT 4.400 83.960 345.600 84.000 ;
        RECT 4.400 82.600 346.000 83.960 ;
        RECT 3.950 81.280 346.000 82.600 ;
        RECT 4.400 79.920 346.000 81.280 ;
        RECT 4.400 79.880 345.600 79.920 ;
        RECT 3.950 78.560 345.600 79.880 ;
        RECT 4.400 78.520 345.600 78.560 ;
        RECT 4.400 77.160 346.000 78.520 ;
        RECT 3.950 75.840 346.000 77.160 ;
        RECT 4.400 74.480 346.000 75.840 ;
        RECT 4.400 74.440 345.600 74.480 ;
        RECT 3.950 73.120 345.600 74.440 ;
        RECT 4.400 73.080 345.600 73.120 ;
        RECT 4.400 71.720 346.000 73.080 ;
        RECT 3.950 70.400 346.000 71.720 ;
        RECT 4.400 69.040 346.000 70.400 ;
        RECT 4.400 69.000 345.600 69.040 ;
        RECT 3.950 67.680 345.600 69.000 ;
        RECT 4.400 67.640 345.600 67.680 ;
        RECT 4.400 66.280 346.000 67.640 ;
        RECT 3.950 64.960 346.000 66.280 ;
        RECT 4.400 63.600 346.000 64.960 ;
        RECT 4.400 63.560 345.600 63.600 ;
        RECT 3.950 62.240 345.600 63.560 ;
        RECT 4.400 62.200 345.600 62.240 ;
        RECT 4.400 60.840 346.000 62.200 ;
        RECT 3.950 59.520 346.000 60.840 ;
        RECT 4.400 58.160 346.000 59.520 ;
        RECT 4.400 58.120 345.600 58.160 ;
        RECT 3.950 56.800 345.600 58.120 ;
        RECT 4.400 56.760 345.600 56.800 ;
        RECT 4.400 55.400 346.000 56.760 ;
        RECT 3.950 54.080 346.000 55.400 ;
        RECT 4.400 52.720 346.000 54.080 ;
        RECT 4.400 52.680 345.600 52.720 ;
        RECT 3.950 51.360 345.600 52.680 ;
        RECT 4.400 51.320 345.600 51.360 ;
        RECT 4.400 49.960 346.000 51.320 ;
        RECT 3.950 48.640 346.000 49.960 ;
        RECT 4.400 47.280 346.000 48.640 ;
        RECT 4.400 47.240 345.600 47.280 ;
        RECT 3.950 45.920 345.600 47.240 ;
        RECT 4.400 45.880 345.600 45.920 ;
        RECT 4.400 44.520 346.000 45.880 ;
        RECT 3.950 43.200 346.000 44.520 ;
        RECT 4.400 41.840 346.000 43.200 ;
        RECT 4.400 41.800 345.600 41.840 ;
        RECT 3.950 40.480 345.600 41.800 ;
        RECT 4.400 40.440 345.600 40.480 ;
        RECT 4.400 39.080 346.000 40.440 ;
        RECT 3.950 37.760 346.000 39.080 ;
        RECT 4.400 36.400 346.000 37.760 ;
        RECT 4.400 36.360 345.600 36.400 ;
        RECT 3.950 35.040 345.600 36.360 ;
        RECT 4.400 35.000 345.600 35.040 ;
        RECT 4.400 33.640 346.000 35.000 ;
        RECT 3.950 32.320 346.000 33.640 ;
        RECT 4.400 30.960 346.000 32.320 ;
        RECT 4.400 30.920 345.600 30.960 ;
        RECT 3.950 29.600 345.600 30.920 ;
        RECT 4.400 29.560 345.600 29.600 ;
        RECT 4.400 28.200 346.000 29.560 ;
        RECT 3.950 26.880 346.000 28.200 ;
        RECT 4.400 25.520 346.000 26.880 ;
        RECT 4.400 25.480 345.600 25.520 ;
        RECT 3.950 24.160 345.600 25.480 ;
        RECT 4.400 24.120 345.600 24.160 ;
        RECT 4.400 22.760 346.000 24.120 ;
        RECT 3.950 21.440 346.000 22.760 ;
        RECT 4.400 20.080 346.000 21.440 ;
        RECT 4.400 20.040 345.600 20.080 ;
        RECT 3.950 18.720 345.600 20.040 ;
        RECT 4.400 18.680 345.600 18.720 ;
        RECT 4.400 17.320 346.000 18.680 ;
        RECT 3.950 16.000 346.000 17.320 ;
        RECT 4.400 14.600 346.000 16.000 ;
        RECT 3.950 13.280 346.000 14.600 ;
        RECT 4.400 11.880 346.000 13.280 ;
        RECT 3.950 10.560 346.000 11.880 ;
        RECT 4.400 9.160 346.000 10.560 ;
        RECT 3.950 7.840 346.000 9.160 ;
        RECT 4.400 6.975 346.000 7.840 ;
      LAYER met4 ;
        RECT 3.975 19.895 20.640 1087.145 ;
        RECT 23.040 19.895 97.440 1087.145 ;
        RECT 99.840 19.895 174.240 1087.145 ;
        RECT 176.640 19.895 251.040 1087.145 ;
        RECT 253.440 19.895 322.625 1087.145 ;
  END
END WishboneInterconnect
END LIBRARY

