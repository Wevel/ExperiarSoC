// This is the unpowered netlist.
module Video (sram0_clk0,
    sram0_clk1,
    sram0_web0,
    sram1_clk0,
    sram1_clk1,
    sram1_web0,
    vga_hsync,
    vga_vsync,
    wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_error_o,
    wb_rst_i,
    wb_stall_o,
    wb_stb_i,
    wb_we_i,
    sram0_addr0,
    sram0_addr1,
    sram0_csb0,
    sram0_csb1,
    sram0_din0,
    sram0_dout0,
    sram0_dout1,
    sram0_wmask0,
    sram1_addr0,
    sram1_addr1,
    sram1_csb0,
    sram1_csb1,
    sram1_din0,
    sram1_dout0,
    sram1_dout1,
    sram1_wmask0,
    vga_b,
    vga_g,
    vga_r,
    video_irq,
    wb_adr_i,
    wb_data_i,
    wb_data_o,
    wb_sel_i);
 output sram0_clk0;
 output sram0_clk1;
 output sram0_web0;
 output sram1_clk0;
 output sram1_clk1;
 output sram1_web0;
 output vga_hsync;
 output vga_vsync;
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 output wb_error_o;
 input wb_rst_i;
 output wb_stall_o;
 input wb_stb_i;
 input wb_we_i;
 output [8:0] sram0_addr0;
 output [8:0] sram0_addr1;
 output [1:0] sram0_csb0;
 output [1:0] sram0_csb1;
 output [31:0] sram0_din0;
 input [63:0] sram0_dout0;
 input [63:0] sram0_dout1;
 output [3:0] sram0_wmask0;
 output [8:0] sram1_addr0;
 output [8:0] sram1_addr1;
 output [1:0] sram1_csb0;
 output [1:0] sram1_csb1;
 output [31:0] sram1_din0;
 input [63:0] sram1_dout0;
 input [63:0] sram1_dout1;
 output [3:0] sram1_wmask0;
 output [1:0] vga_b;
 output [1:0] vga_g;
 output [1:0] vga_r;
 output [1:0] video_irq;
 input [23:0] wb_adr_i;
 input [31:0] wb_data_i;
 output [31:0] wb_data_o;
 input [3:0] wb_sel_i;

 wire net619;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \vga.configuration[0] ;
 wire \vga.configuration[10] ;
 wire \vga.configuration[11] ;
 wire \vga.configuration[12] ;
 wire \vga.configuration[1] ;
 wire \vga.configuration[2] ;
 wire \vga.configuration[3] ;
 wire \vga.configuration[4] ;
 wire \vga.configuration[5] ;
 wire \vga.configuration[6] ;
 wire \vga.configuration[7] ;
 wire \vga.configuration[8] ;
 wire \vga.configuration[9] ;
 wire \vga.currentPixelData[0] ;
 wire \vga.currentPixelData[10] ;
 wire \vga.currentPixelData[11] ;
 wire \vga.currentPixelData[12] ;
 wire \vga.currentPixelData[13] ;
 wire \vga.currentPixelData[14] ;
 wire \vga.currentPixelData[15] ;
 wire \vga.currentPixelData[16] ;
 wire \vga.currentPixelData[17] ;
 wire \vga.currentPixelData[18] ;
 wire \vga.currentPixelData[19] ;
 wire \vga.currentPixelData[1] ;
 wire \vga.currentPixelData[20] ;
 wire \vga.currentPixelData[21] ;
 wire \vga.currentPixelData[22] ;
 wire \vga.currentPixelData[23] ;
 wire \vga.currentPixelData[24] ;
 wire \vga.currentPixelData[25] ;
 wire \vga.currentPixelData[26] ;
 wire \vga.currentPixelData[27] ;
 wire \vga.currentPixelData[28] ;
 wire \vga.currentPixelData[29] ;
 wire \vga.currentPixelData[2] ;
 wire \vga.currentPixelData[3] ;
 wire \vga.currentPixelData[4] ;
 wire \vga.currentPixelData[5] ;
 wire \vga.currentPixelData[6] ;
 wire \vga.currentPixelData[7] ;
 wire \vga.currentPixelData[8] ;
 wire \vga.currentPixelData[9] ;
 wire \vga.horizontalCounter[0] ;
 wire \vga.horizontalCounter[10] ;
 wire \vga.horizontalCounter[1] ;
 wire \vga.horizontalCounter[2] ;
 wire \vga.horizontalCounter[3] ;
 wire \vga.horizontalCounter[4] ;
 wire \vga.horizontalCounter[5] ;
 wire \vga.horizontalCounter[6] ;
 wire \vga.horizontalCounter[7] ;
 wire \vga.horizontalCounter[8] ;
 wire \vga.horizontalCounter[9] ;
 wire \vga.horizontalFrontPorchCompare[0] ;
 wire \vga.horizontalFrontPorchCompare[10] ;
 wire \vga.horizontalFrontPorchCompare[1] ;
 wire \vga.horizontalFrontPorchCompare[2] ;
 wire \vga.horizontalFrontPorchCompare[3] ;
 wire \vga.horizontalFrontPorchCompare[4] ;
 wire \vga.horizontalFrontPorchCompare[5] ;
 wire \vga.horizontalFrontPorchCompare[6] ;
 wire \vga.horizontalFrontPorchCompare[7] ;
 wire \vga.horizontalFrontPorchCompare[8] ;
 wire \vga.horizontalFrontPorchCompare[9] ;
 wire \vga.horizontalSyncPulseCompare[0] ;
 wire \vga.horizontalSyncPulseCompare[10] ;
 wire \vga.horizontalSyncPulseCompare[1] ;
 wire \vga.horizontalSyncPulseCompare[2] ;
 wire \vga.horizontalSyncPulseCompare[3] ;
 wire \vga.horizontalSyncPulseCompare[4] ;
 wire \vga.horizontalSyncPulseCompare[5] ;
 wire \vga.horizontalSyncPulseCompare[6] ;
 wire \vga.horizontalSyncPulseCompare[7] ;
 wire \vga.horizontalSyncPulseCompare[8] ;
 wire \vga.horizontalSyncPulseCompare[9] ;
 wire \vga.horizontalVisibleAreaCompare[0] ;
 wire \vga.horizontalVisibleAreaCompare[10] ;
 wire \vga.horizontalVisibleAreaCompare[1] ;
 wire \vga.horizontalVisibleAreaCompare[2] ;
 wire \vga.horizontalVisibleAreaCompare[3] ;
 wire \vga.horizontalVisibleAreaCompare[4] ;
 wire \vga.horizontalVisibleAreaCompare[5] ;
 wire \vga.horizontalVisibleAreaCompare[6] ;
 wire \vga.horizontalVisibleAreaCompare[7] ;
 wire \vga.horizontalVisibleAreaCompare[8] ;
 wire \vga.horizontalVisibleAreaCompare[9] ;
 wire \vga.horizontalWholeLineCompare[0] ;
 wire \vga.horizontalWholeLineCompare[10] ;
 wire \vga.horizontalWholeLineCompare[1] ;
 wire \vga.horizontalWholeLineCompare[2] ;
 wire \vga.horizontalWholeLineCompare[3] ;
 wire \vga.horizontalWholeLineCompare[4] ;
 wire \vga.horizontalWholeLineCompare[5] ;
 wire \vga.horizontalWholeLineCompare[6] ;
 wire \vga.horizontalWholeLineCompare[7] ;
 wire \vga.horizontalWholeLineCompare[8] ;
 wire \vga.horizontalWholeLineCompare[9] ;
 wire \vga.hsync ;
 wire \vga.inHorizontalVisibleArea ;
 wire \vga.inVerticalVisibleArea ;
 wire \vga.lastHSync ;
 wire \vga.lastVSync ;
 wire \vga.loadPixelData ;
 wire \vga.raw_directPixelCounterVertical[0] ;
 wire \vga.raw_directPixelCounterVertical[10] ;
 wire \vga.raw_directPixelCounterVertical[1] ;
 wire \vga.raw_directPixelCounterVertical[2] ;
 wire \vga.raw_directPixelCounterVertical[3] ;
 wire \vga.raw_directPixelCounterVertical[4] ;
 wire \vga.raw_directPixelCounterVertical[5] ;
 wire \vga.raw_directPixelCounterVertical[6] ;
 wire \vga.raw_directPixelCounterVertical[7] ;
 wire \vga.raw_directPixelCounterVertical[8] ;
 wire \vga.raw_directPixelCounterVertical[9] ;
 wire \vga.raw_horizontalPixelCounter[0] ;
 wire \vga.raw_horizontalPixelCounter[1] ;
 wire \vga.raw_horizontalPixelCounter[2] ;
 wire \vga.raw_horizontalPixelCounter[3] ;
 wire \vga.raw_horizontalPixelCounter[4] ;
 wire \vga.raw_horizontalPixelCounter[5] ;
 wire \vga.raw_horizontalPixelCounter[6] ;
 wire \vga.raw_horizontalPixelCounter[7] ;
 wire \vga.raw_horizontalPixelCounter[8] ;
 wire \vga.raw_horizontalPixelStretchCounter[0] ;
 wire \vga.raw_horizontalPixelStretchCounter[1] ;
 wire \vga.raw_horizontalPixelStretchCounter[2] ;
 wire \vga.raw_horizontalPixelStretchCounter[3] ;
 wire \vga.raw_subPixelCounter[0] ;
 wire \vga.raw_subPixelCounter[1] ;
 wire \vga.raw_subPixelCounter[2] ;
 wire \vga.raw_subPixelCounter_buffered[0] ;
 wire \vga.raw_subPixelCounter_buffered[1] ;
 wire \vga.raw_subPixelCounter_buffered[2] ;
 wire \vga.raw_verticalPixelCounter[0] ;
 wire \vga.raw_verticalPixelCounter[1] ;
 wire \vga.raw_verticalPixelCounter[2] ;
 wire \vga.raw_verticalPixelCounter[3] ;
 wire \vga.raw_verticalPixelCounter[4] ;
 wire \vga.raw_verticalPixelCounter[5] ;
 wire \vga.raw_verticalPixelCounter[6] ;
 wire \vga.raw_verticalPixelCounter[7] ;
 wire \vga.raw_verticalPixelCounter[8] ;
 wire \vga.raw_verticalPixelCounter[9] ;
 wire \vga.raw_verticalPixelStretchCounter[0] ;
 wire \vga.raw_verticalPixelStretchCounter[1] ;
 wire \vga.raw_verticalPixelStretchCounter[2] ;
 wire \vga.raw_verticalPixelStretchCounter[3] ;
 wire \vga.stateRegister.baseReadData[0] ;
 wire \vga.stateRegister.baseReadData[1] ;
 wire \vga.stateRegister.baseReadData[2] ;
 wire \vga.stateRegister.baseReadData[3] ;
 wire \vga.stateRegister.baseReadData[4] ;
 wire \vga.verticalCounter[0] ;
 wire \vga.verticalCounter[1] ;
 wire \vga.verticalCounter[2] ;
 wire \vga.verticalCounter[3] ;
 wire \vga.verticalCounter[4] ;
 wire \vga.verticalCounter[5] ;
 wire \vga.verticalCounter[6] ;
 wire \vga.verticalCounter[7] ;
 wire \vga.verticalCounter[8] ;
 wire \vga.verticalCounter[9] ;
 wire \vga.verticalFrontPorchCompare[0] ;
 wire \vga.verticalFrontPorchCompare[1] ;
 wire \vga.verticalFrontPorchCompare[2] ;
 wire \vga.verticalFrontPorchCompare[3] ;
 wire \vga.verticalFrontPorchCompare[4] ;
 wire \vga.verticalFrontPorchCompare[5] ;
 wire \vga.verticalFrontPorchCompare[6] ;
 wire \vga.verticalFrontPorchCompare[7] ;
 wire \vga.verticalFrontPorchCompare[8] ;
 wire \vga.verticalFrontPorchCompare[9] ;
 wire \vga.verticalSyncPulseCompare[0] ;
 wire \vga.verticalSyncPulseCompare[1] ;
 wire \vga.verticalSyncPulseCompare[2] ;
 wire \vga.verticalSyncPulseCompare[3] ;
 wire \vga.verticalSyncPulseCompare[4] ;
 wire \vga.verticalSyncPulseCompare[5] ;
 wire \vga.verticalSyncPulseCompare[6] ;
 wire \vga.verticalSyncPulseCompare[7] ;
 wire \vga.verticalSyncPulseCompare[8] ;
 wire \vga.verticalSyncPulseCompare[9] ;
 wire \vga.verticalVisibleAreaCompare[0] ;
 wire \vga.verticalVisibleAreaCompare[1] ;
 wire \vga.verticalVisibleAreaCompare[2] ;
 wire \vga.verticalVisibleAreaCompare[3] ;
 wire \vga.verticalVisibleAreaCompare[4] ;
 wire \vga.verticalVisibleAreaCompare[5] ;
 wire \vga.verticalVisibleAreaCompare[6] ;
 wire \vga.verticalVisibleAreaCompare[7] ;
 wire \vga.verticalVisibleAreaCompare[8] ;
 wire \vga.verticalVisibleAreaCompare[9] ;
 wire \vga.verticalWholeLineCompare[0] ;
 wire \vga.verticalWholeLineCompare[1] ;
 wire \vga.verticalWholeLineCompare[2] ;
 wire \vga.verticalWholeLineCompare[3] ;
 wire \vga.verticalWholeLineCompare[4] ;
 wire \vga.verticalWholeLineCompare[5] ;
 wire \vga.verticalWholeLineCompare[6] ;
 wire \vga.verticalWholeLineCompare[7] ;
 wire \vga.verticalWholeLineCompare[8] ;
 wire \vga.verticalWholeLineCompare[9] ;
 wire \vga.vsync ;
 wire \videoMemory.wbReadReady ;
 wire \wbPeripheralBusInterface.currentAddress[10] ;
 wire \wbPeripheralBusInterface.currentAddress[11] ;
 wire \wbPeripheralBusInterface.currentAddress[12] ;
 wire \wbPeripheralBusInterface.currentAddress[13] ;
 wire \wbPeripheralBusInterface.currentAddress[14] ;
 wire \wbPeripheralBusInterface.currentAddress[15] ;
 wire \wbPeripheralBusInterface.currentAddress[16] ;
 wire \wbPeripheralBusInterface.currentAddress[17] ;
 wire \wbPeripheralBusInterface.currentAddress[18] ;
 wire \wbPeripheralBusInterface.currentAddress[19] ;
 wire \wbPeripheralBusInterface.currentAddress[20] ;
 wire \wbPeripheralBusInterface.currentAddress[21] ;
 wire \wbPeripheralBusInterface.currentAddress[22] ;
 wire \wbPeripheralBusInterface.currentAddress[23] ;
 wire \wbPeripheralBusInterface.currentAddress[2] ;
 wire \wbPeripheralBusInterface.currentAddress[3] ;
 wire \wbPeripheralBusInterface.currentAddress[4] ;
 wire \wbPeripheralBusInterface.currentAddress[5] ;
 wire \wbPeripheralBusInterface.currentAddress[6] ;
 wire \wbPeripheralBusInterface.currentAddress[7] ;
 wire \wbPeripheralBusInterface.currentAddress[8] ;
 wire \wbPeripheralBusInterface.currentAddress[9] ;
 wire \wbPeripheralBusInterface.currentByteSelect[0] ;
 wire \wbPeripheralBusInterface.currentByteSelect[1] ;
 wire \wbPeripheralBusInterface.currentByteSelect[2] ;
 wire \wbPeripheralBusInterface.currentByteSelect[3] ;
 wire \wbPeripheralBusInterface.state[0] ;
 wire \wbPeripheralBusInterface.state[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net366));
 sky130_fd_sc_hd__decap_4 FILLER_0_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_94 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__conb_1 Video_619 (.LO(net619));
 sky130_fd_sc_hd__inv_2 _1358_ (.A(\vga.verticalWholeLineCompare[0] ),
    .Y(_1291_));
 sky130_fd_sc_hd__inv_2 _1359_ (.A(\vga.verticalWholeLineCompare[1] ),
    .Y(_1292_));
 sky130_fd_sc_hd__inv_2 _1360_ (.A(\vga.verticalWholeLineCompare[4] ),
    .Y(_1293_));
 sky130_fd_sc_hd__inv_2 _1361_ (.A(\vga.verticalWholeLineCompare[5] ),
    .Y(_1294_));
 sky130_fd_sc_hd__inv_2 _1362_ (.A(\vga.verticalWholeLineCompare[6] ),
    .Y(_1295_));
 sky130_fd_sc_hd__inv_2 _1363_ (.A(\vga.verticalWholeLineCompare[7] ),
    .Y(_1296_));
 sky130_fd_sc_hd__inv_2 _1364_ (.A(\vga.verticalSyncPulseCompare[1] ),
    .Y(_1297_));
 sky130_fd_sc_hd__inv_2 _1365_ (.A(\vga.verticalSyncPulseCompare[2] ),
    .Y(_1298_));
 sky130_fd_sc_hd__inv_2 _1366_ (.A(\vga.verticalSyncPulseCompare[3] ),
    .Y(_1299_));
 sky130_fd_sc_hd__inv_2 _1367_ (.A(\vga.verticalSyncPulseCompare[6] ),
    .Y(_1300_));
 sky130_fd_sc_hd__inv_2 _1368_ (.A(\vga.verticalFrontPorchCompare[0] ),
    .Y(_1301_));
 sky130_fd_sc_hd__inv_2 _1369_ (.A(\vga.verticalFrontPorchCompare[2] ),
    .Y(_1302_));
 sky130_fd_sc_hd__inv_2 _1370_ (.A(\vga.verticalVisibleAreaCompare[5] ),
    .Y(_1303_));
 sky130_fd_sc_hd__inv_2 _1371_ (.A(\vga.verticalVisibleAreaCompare[8] ),
    .Y(_1304_));
 sky130_fd_sc_hd__inv_2 _1372_ (.A(\vga.horizontalWholeLineCompare[5] ),
    .Y(_1305_));
 sky130_fd_sc_hd__inv_2 _1373_ (.A(\vga.horizontalWholeLineCompare[6] ),
    .Y(_1306_));
 sky130_fd_sc_hd__inv_2 _1374_ (.A(\vga.horizontalWholeLineCompare[7] ),
    .Y(_1307_));
 sky130_fd_sc_hd__inv_2 _1375_ (.A(\vga.horizontalSyncPulseCompare[0] ),
    .Y(_1308_));
 sky130_fd_sc_hd__inv_2 _1376_ (.A(\vga.horizontalSyncPulseCompare[3] ),
    .Y(_1309_));
 sky130_fd_sc_hd__inv_2 _1377_ (.A(\vga.horizontalSyncPulseCompare[6] ),
    .Y(_1310_));
 sky130_fd_sc_hd__inv_2 _1378_ (.A(\vga.horizontalSyncPulseCompare[9] ),
    .Y(_1311_));
 sky130_fd_sc_hd__inv_2 _1379_ (.A(\vga.horizontalFrontPorchCompare[2] ),
    .Y(_1312_));
 sky130_fd_sc_hd__inv_2 _1380_ (.A(\vga.horizontalFrontPorchCompare[4] ),
    .Y(_1313_));
 sky130_fd_sc_hd__inv_2 _1381_ (.A(\vga.horizontalFrontPorchCompare[6] ),
    .Y(_1314_));
 sky130_fd_sc_hd__inv_2 _1382_ (.A(\vga.horizontalVisibleAreaCompare[7] ),
    .Y(_1315_));
 sky130_fd_sc_hd__inv_2 _1383_ (.A(\vga.horizontalVisibleAreaCompare[8] ),
    .Y(_1316_));
 sky130_fd_sc_hd__inv_2 _1384_ (.A(\vga.horizontalVisibleAreaCompare[9] ),
    .Y(_1317_));
 sky130_fd_sc_hd__inv_2 _1385_ (.A(\vga.verticalCounter[9] ),
    .Y(_1318_));
 sky130_fd_sc_hd__clkinv_4 _1386_ (.A(\vga.verticalCounter[8] ),
    .Y(_1319_));
 sky130_fd_sc_hd__clkinv_2 _1387_ (.A(\vga.verticalCounter[7] ),
    .Y(_1320_));
 sky130_fd_sc_hd__clkinv_2 _1388_ (.A(\vga.verticalCounter[6] ),
    .Y(_1321_));
 sky130_fd_sc_hd__inv_2 _1389_ (.A(\vga.verticalCounter[5] ),
    .Y(_1322_));
 sky130_fd_sc_hd__clkinv_2 _1390_ (.A(\vga.verticalCounter[4] ),
    .Y(_1323_));
 sky130_fd_sc_hd__clkinv_2 _1391_ (.A(\vga.verticalCounter[3] ),
    .Y(_1324_));
 sky130_fd_sc_hd__clkinv_4 _1392_ (.A(\vga.verticalCounter[2] ),
    .Y(_1325_));
 sky130_fd_sc_hd__inv_2 _1393_ (.A(\vga.verticalCounter[1] ),
    .Y(_1326_));
 sky130_fd_sc_hd__inv_2 _1394_ (.A(\vga.verticalCounter[0] ),
    .Y(_1327_));
 sky130_fd_sc_hd__inv_2 _1395_ (.A(net593),
    .Y(_1328_));
 sky130_fd_sc_hd__inv_2 _1396_ (.A(\vga.raw_subPixelCounter[0] ),
    .Y(_1329_));
 sky130_fd_sc_hd__inv_2 _1397_ (.A(net443),
    .Y(_1330_));
 sky130_fd_sc_hd__inv_2 _1398_ (.A(net610),
    .Y(_1331_));
 sky130_fd_sc_hd__clkinv_4 _1399_ (.A(\vga.horizontalCounter[0] ),
    .Y(_1332_));
 sky130_fd_sc_hd__inv_2 _1400_ (.A(\vga.horizontalCounter[1] ),
    .Y(_1333_));
 sky130_fd_sc_hd__clkinv_2 _1401_ (.A(\vga.horizontalCounter[2] ),
    .Y(_1334_));
 sky130_fd_sc_hd__inv_2 _1402_ (.A(\vga.horizontalCounter[3] ),
    .Y(_1335_));
 sky130_fd_sc_hd__inv_2 _1403_ (.A(\vga.horizontalCounter[4] ),
    .Y(_1336_));
 sky130_fd_sc_hd__inv_2 _1404_ (.A(\vga.horizontalCounter[5] ),
    .Y(_1337_));
 sky130_fd_sc_hd__inv_2 _1405_ (.A(\vga.horizontalCounter[6] ),
    .Y(_1338_));
 sky130_fd_sc_hd__clkinv_4 _1406_ (.A(\vga.horizontalCounter[7] ),
    .Y(_1339_));
 sky130_fd_sc_hd__inv_2 _1407_ (.A(\vga.horizontalCounter[8] ),
    .Y(_1340_));
 sky130_fd_sc_hd__inv_2 _1408_ (.A(\vga.horizontalCounter[9] ),
    .Y(_1341_));
 sky130_fd_sc_hd__clkinv_4 _1409_ (.A(\vga.horizontalCounter[10] ),
    .Y(_1342_));
 sky130_fd_sc_hd__inv_6 _1410_ (.A(net302),
    .Y(_1343_));
 sky130_fd_sc_hd__inv_6 _1411_ (.A(net303),
    .Y(_1344_));
 sky130_fd_sc_hd__clkinv_2 _1412_ (.A(net595),
    .Y(_1345_));
 sky130_fd_sc_hd__clkinv_4 _1413_ (.A(\vga.raw_horizontalPixelCounter[4] ),
    .Y(_1346_));
 sky130_fd_sc_hd__inv_2 _1414_ (.A(\vga.raw_directPixelCounterVertical[9] ),
    .Y(_1347_));
 sky130_fd_sc_hd__inv_2 _1415_ (.A(\vga.raw_directPixelCounterVertical[5] ),
    .Y(_1348_));
 sky130_fd_sc_hd__inv_2 _1416_ (.A(\vga.raw_directPixelCounterVertical[1] ),
    .Y(_1349_));
 sky130_fd_sc_hd__inv_2 _1417_ (.A(\vga.raw_directPixelCounterVertical[0] ),
    .Y(_1350_));
 sky130_fd_sc_hd__and2b_4 _1418_ (.A_N(\wbPeripheralBusInterface.state[1] ),
    .B(\wbPeripheralBusInterface.state[0] ),
    .X(_1351_));
 sky130_fd_sc_hd__nand2b_4 _1419_ (.A_N(\wbPeripheralBusInterface.state[1] ),
    .B(\wbPeripheralBusInterface.state[0] ),
    .Y(_1352_));
 sky130_fd_sc_hd__and2_4 _1420_ (.A(net272),
    .B(net582),
    .X(net335));
 sky130_fd_sc_hd__and2_4 _1421_ (.A(net283),
    .B(net582),
    .X(net346));
 sky130_fd_sc_hd__and2_4 _1422_ (.A(net294),
    .B(net582),
    .X(net357));
 sky130_fd_sc_hd__and2_4 _1423_ (.A(net297),
    .B(net582),
    .X(net360));
 sky130_fd_sc_hd__and2_4 _1424_ (.A(net298),
    .B(net582),
    .X(net361));
 sky130_fd_sc_hd__and2_4 _1425_ (.A(net299),
    .B(net582),
    .X(net362));
 sky130_fd_sc_hd__and2_4 _1426_ (.A(net300),
    .B(net582),
    .X(net363));
 sky130_fd_sc_hd__and2_4 _1427_ (.A(net301),
    .B(net582),
    .X(net364));
 sky130_fd_sc_hd__nor2_8 _1428_ (.A(_1343_),
    .B(_1352_),
    .Y(net365));
 sky130_fd_sc_hd__nor2_8 _1429_ (.A(_1344_),
    .B(_1352_),
    .Y(net366));
 sky130_fd_sc_hd__and2_4 _1430_ (.A(net273),
    .B(net584),
    .X(net336));
 sky130_fd_sc_hd__and2_4 _1431_ (.A(net274),
    .B(net582),
    .X(net337));
 sky130_fd_sc_hd__and2_4 _1432_ (.A(net275),
    .B(net584),
    .X(net338));
 sky130_fd_sc_hd__nor2_1 _1433_ (.A(\wbPeripheralBusInterface.state[1] ),
    .B(\wbPeripheralBusInterface.state[0] ),
    .Y(_1353_));
 sky130_fd_sc_hd__or2_4 _1434_ (.A(\wbPeripheralBusInterface.state[1] ),
    .B(\wbPeripheralBusInterface.state[0] ),
    .X(_1354_));
 sky130_fd_sc_hd__nand2_4 _1435_ (.A(\wbPeripheralBusInterface.currentAddress[4] ),
    .B(net580),
    .Y(_1355_));
 sky130_fd_sc_hd__clkinv_4 _1436_ (.A(_1355_),
    .Y(net313));
 sky130_fd_sc_hd__nand2_2 _1437_ (.A(\wbPeripheralBusInterface.currentAddress[2] ),
    .B(net580),
    .Y(_1356_));
 sky130_fd_sc_hd__clkinv_4 _1438_ (.A(_1356_),
    .Y(net311));
 sky130_fd_sc_hd__nand2_2 _1439_ (.A(\wbPeripheralBusInterface.currentAddress[3] ),
    .B(net580),
    .Y(_1357_));
 sky130_fd_sc_hd__clkinv_4 _1440_ (.A(_1357_),
    .Y(net312));
 sky130_fd_sc_hd__nand2_8 _1441_ (.A(\wbPeripheralBusInterface.currentAddress[5] ),
    .B(net580),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_4 _1442_ (.A(_0267_),
    .Y(net314));
 sky130_fd_sc_hd__and2_4 _1443_ (.A(\wbPeripheralBusInterface.currentAddress[6] ),
    .B(net581),
    .X(net315));
 sky130_fd_sc_hd__and2_4 _1444_ (.A(\wbPeripheralBusInterface.currentAddress[7] ),
    .B(net581),
    .X(net316));
 sky130_fd_sc_hd__and2_4 _1445_ (.A(\wbPeripheralBusInterface.currentAddress[8] ),
    .B(net581),
    .X(net317));
 sky130_fd_sc_hd__and2_4 _1446_ (.A(\wbPeripheralBusInterface.currentAddress[9] ),
    .B(net581),
    .X(net318));
 sky130_fd_sc_hd__and2_4 _1447_ (.A(\wbPeripheralBusInterface.currentAddress[10] ),
    .B(net581),
    .X(net319));
 sky130_fd_sc_hd__or3_1 _1448_ (.A(\wbPeripheralBusInterface.currentAddress[13] ),
    .B(\wbPeripheralBusInterface.currentAddress[19] ),
    .C(\wbPeripheralBusInterface.currentAddress[21] ),
    .X(_0268_));
 sky130_fd_sc_hd__or3_2 _1449_ (.A(\wbPeripheralBusInterface.currentAddress[20] ),
    .B(\wbPeripheralBusInterface.currentAddress[22] ),
    .C(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__or3_4 _1450_ (.A(\wbPeripheralBusInterface.currentAddress[14] ),
    .B(\wbPeripheralBusInterface.currentAddress[15] ),
    .C(\wbPeripheralBusInterface.currentAddress[18] ),
    .X(_0270_));
 sky130_fd_sc_hd__or2_1 _1451_ (.A(\wbPeripheralBusInterface.currentAddress[16] ),
    .B(\wbPeripheralBusInterface.currentAddress[17] ),
    .X(_0271_));
 sky130_fd_sc_hd__or4_4 _1452_ (.A(\wbPeripheralBusInterface.currentAddress[23] ),
    .B(_0269_),
    .C(_0270_),
    .D(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__or2_4 _1453_ (.A(_1352_),
    .B(_0272_),
    .X(net367));
 sky130_fd_sc_hd__nand2b_4 _1454_ (.A_N(\vga.vsync ),
    .B(\vga.configuration[10] ),
    .Y(net440));
 sky130_fd_sc_hd__nand2b_4 _1455_ (.A_N(\vga.hsync ),
    .B(\vga.configuration[10] ),
    .Y(net437));
 sky130_fd_sc_hd__and2_4 _1456_ (.A(\wbPeripheralBusInterface.currentByteSelect[3] ),
    .B(net581),
    .X(net371));
 sky130_fd_sc_hd__and2_4 _1457_ (.A(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .B(net581),
    .X(net370));
 sky130_fd_sc_hd__and2_1 _1458_ (.A(net596),
    .B(net580),
    .X(net369));
 sky130_fd_sc_hd__and2_1 _1459_ (.A(net602),
    .B(net580),
    .X(net368));
 sky130_fd_sc_hd__and3b_4 _1460_ (.A_N(\vga.vsync ),
    .B(\vga.lastVSync ),
    .C(\vga.configuration[12] ),
    .X(net442));
 sky130_fd_sc_hd__and3b_2 _1461_ (.A_N(\vga.hsync ),
    .B(\vga.lastHSync ),
    .C(\vga.configuration[11] ),
    .X(net441));
 sky130_fd_sc_hd__and2_4 _1462_ (.A(net276),
    .B(net583),
    .X(net339));
 sky130_fd_sc_hd__and2_4 _1463_ (.A(net277),
    .B(net582),
    .X(net340));
 sky130_fd_sc_hd__and2_4 _1464_ (.A(net278),
    .B(net585),
    .X(net341));
 sky130_fd_sc_hd__and2_4 _1465_ (.A(net279),
    .B(net585),
    .X(net342));
 sky130_fd_sc_hd__and2_4 _1466_ (.A(net280),
    .B(net585),
    .X(net343));
 sky130_fd_sc_hd__and2_4 _1467_ (.A(net281),
    .B(net585),
    .X(net344));
 sky130_fd_sc_hd__and2_4 _1468_ (.A(net282),
    .B(net585),
    .X(net345));
 sky130_fd_sc_hd__and2_4 _1469_ (.A(net284),
    .B(net585),
    .X(net347));
 sky130_fd_sc_hd__and2_4 _1470_ (.A(net285),
    .B(net585),
    .X(net348));
 sky130_fd_sc_hd__and2_4 _1471_ (.A(net286),
    .B(net586),
    .X(net349));
 sky130_fd_sc_hd__and2_4 _1472_ (.A(net287),
    .B(net586),
    .X(net350));
 sky130_fd_sc_hd__and2_4 _1473_ (.A(net288),
    .B(net586),
    .X(net351));
 sky130_fd_sc_hd__and2_4 _1474_ (.A(net289),
    .B(net586),
    .X(net352));
 sky130_fd_sc_hd__and2_4 _1475_ (.A(net290),
    .B(net585),
    .X(net353));
 sky130_fd_sc_hd__and2_4 _1476_ (.A(net291),
    .B(net585),
    .X(net354));
 sky130_fd_sc_hd__and2_4 _1477_ (.A(net292),
    .B(net585),
    .X(net355));
 sky130_fd_sc_hd__and2_4 _1478_ (.A(net293),
    .B(net586),
    .X(net356));
 sky130_fd_sc_hd__and2_4 _1479_ (.A(net295),
    .B(net586),
    .X(net358));
 sky130_fd_sc_hd__and2_4 _1480_ (.A(net296),
    .B(net586),
    .X(net359));
 sky130_fd_sc_hd__o21ai_4 _1481_ (.A1(\wbPeripheralBusInterface.currentAddress[12] ),
    .A2(\wbPeripheralBusInterface.currentAddress[11] ),
    .B1(_1354_),
    .Y(_0273_));
 sky130_fd_sc_hd__o21a_1 _1482_ (.A1(\wbPeripheralBusInterface.currentAddress[12] ),
    .A2(\wbPeripheralBusInterface.currentAddress[11] ),
    .B1(net580),
    .X(_0274_));
 sky130_fd_sc_hd__and2b_4 _1483_ (.A_N(\wbPeripheralBusInterface.state[0] ),
    .B(\wbPeripheralBusInterface.state[1] ),
    .X(_0275_));
 sky130_fd_sc_hd__nand2b_2 _1484_ (.A_N(\wbPeripheralBusInterface.state[0] ),
    .B(\wbPeripheralBusInterface.state[1] ),
    .Y(_0276_));
 sky130_fd_sc_hd__or2_2 _1485_ (.A(_0272_),
    .B(net578),
    .X(_0277_));
 sky130_fd_sc_hd__inv_2 _1486_ (.A(net530),
    .Y(_0278_));
 sky130_fd_sc_hd__nand2_8 _1487_ (.A(net367),
    .B(net530),
    .Y(_0279_));
 sky130_fd_sc_hd__nand2_1 _1488_ (.A(net564),
    .B(_0279_),
    .Y(net331));
 sky130_fd_sc_hd__and3b_4 _1489_ (.A_N(\wbPeripheralBusInterface.currentAddress[12] ),
    .B(\wbPeripheralBusInterface.currentAddress[11] ),
    .C(net580),
    .X(_0280_));
 sky130_fd_sc_hd__nand2_1 _1490_ (.A(_0279_),
    .B(net554),
    .Y(net332));
 sky130_fd_sc_hd__and3b_4 _1491_ (.A_N(\wbPeripheralBusInterface.currentAddress[11] ),
    .B(_1354_),
    .C(\wbPeripheralBusInterface.currentAddress[12] ),
    .X(_0281_));
 sky130_fd_sc_hd__nand2_1 _1492_ (.A(_0279_),
    .B(_0281_),
    .Y(net392));
 sky130_fd_sc_hd__and3_4 _1493_ (.A(\wbPeripheralBusInterface.currentAddress[12] ),
    .B(\wbPeripheralBusInterface.currentAddress[11] ),
    .C(_1354_),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _1494_ (.A(_0279_),
    .B(_0282_),
    .Y(net393));
 sky130_fd_sc_hd__nand2_8 _1495_ (.A(\vga.configuration[10] ),
    .B(net606),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_2 _1496_ (.A(_0283_),
    .Y(_0059_));
 sky130_fd_sc_hd__and2_1 _1497_ (.A(\vga.inHorizontalVisibleArea ),
    .B(net608),
    .X(_0062_));
 sky130_fd_sc_hd__and3_4 _1498_ (.A(\vga.configuration[10] ),
    .B(\vga.inHorizontalVisibleArea ),
    .C(\vga.inVerticalVisibleArea ),
    .X(_0284_));
 sky130_fd_sc_hd__and2_4 _1499_ (.A(net608),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__nand2_4 _1500_ (.A(net606),
    .B(_0284_),
    .Y(_0286_));
 sky130_fd_sc_hd__and3b_2 _1501_ (.A_N(\vga.raw_subPixelCounter[1] ),
    .B(_1329_),
    .C(\vga.raw_subPixelCounter[2] ),
    .X(_0287_));
 sky130_fd_sc_hd__nand3_4 _1502_ (.A(\vga.raw_horizontalPixelStretchCounter[0] ),
    .B(\vga.raw_horizontalPixelStretchCounter[1] ),
    .C(\vga.raw_horizontalPixelStretchCounter[2] ),
    .Y(_0288_));
 sky130_fd_sc_hd__xor2_4 _1503_ (.A(\vga.raw_horizontalPixelStretchCounter[3] ),
    .B(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__xor2_4 _1504_ (.A(\vga.configuration[3] ),
    .B(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__xnor2_2 _1505_ (.A(\vga.raw_horizontalPixelStretchCounter[0] ),
    .B(\vga.raw_horizontalPixelStretchCounter[1] ),
    .Y(_0291_));
 sky130_fd_sc_hd__xor2_1 _1506_ (.A(\vga.configuration[1] ),
    .B(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__nand2_1 _1507_ (.A(\vga.configuration[0] ),
    .B(\vga.raw_horizontalPixelStretchCounter[0] ),
    .Y(_0293_));
 sky130_fd_sc_hd__or2_1 _1508_ (.A(\vga.configuration[0] ),
    .B(\vga.raw_horizontalPixelStretchCounter[0] ),
    .X(_0294_));
 sky130_fd_sc_hd__a21o_1 _1509_ (.A1(\vga.raw_horizontalPixelStretchCounter[0] ),
    .A2(\vga.raw_horizontalPixelStretchCounter[1] ),
    .B1(\vga.raw_horizontalPixelStretchCounter[2] ),
    .X(_0295_));
 sky130_fd_sc_hd__a21oi_1 _1510_ (.A1(_0288_),
    .A2(_0295_),
    .B1(\vga.configuration[2] ),
    .Y(_0296_));
 sky130_fd_sc_hd__and3_1 _1511_ (.A(\vga.configuration[2] ),
    .B(_0288_),
    .C(_0295_),
    .X(_0297_));
 sky130_fd_sc_hd__o2111a_2 _1512_ (.A1(_0296_),
    .A2(_0297_),
    .B1(_0292_),
    .C1(_0293_),
    .D1(_0294_),
    .X(_0298_));
 sky130_fd_sc_hd__nand2_2 _1513_ (.A(_0290_),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__and3_4 _1514_ (.A(_0287_),
    .B(_0290_),
    .C(_0298_),
    .X(_0300_));
 sky130_fd_sc_hd__and3_4 _1515_ (.A(net595),
    .B(\vga.raw_horizontalPixelCounter[1] ),
    .C(\vga.raw_horizontalPixelCounter[2] ),
    .X(_0301_));
 sky130_fd_sc_hd__and4_4 _1516_ (.A(net595),
    .B(\vga.raw_horizontalPixelCounter[1] ),
    .C(\vga.raw_horizontalPixelCounter[2] ),
    .D(\vga.raw_horizontalPixelCounter[3] ),
    .X(_0302_));
 sky130_fd_sc_hd__and3_2 _1517_ (.A(\vga.raw_horizontalPixelCounter[4] ),
    .B(\vga.raw_horizontalPixelCounter[5] ),
    .C(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__a21oi_2 _1518_ (.A1(\vga.raw_horizontalPixelCounter[4] ),
    .A2(_0302_),
    .B1(\vga.raw_horizontalPixelCounter[5] ),
    .Y(_0304_));
 sky130_fd_sc_hd__nor2_4 _1519_ (.A(_0303_),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__nor2_8 _1520_ (.A(_0286_),
    .B(_0300_),
    .Y(_0306_));
 sky130_fd_sc_hd__or2_2 _1521_ (.A(_0286_),
    .B(_0300_),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_2 _1522_ (.A(_0285_),
    .B(_0305_),
    .Y(_0308_));
 sky130_fd_sc_hd__and2_4 _1523_ (.A(_0285_),
    .B(_0300_),
    .X(_0309_));
 sky130_fd_sc_hd__or4_1 _1524_ (.A(net595),
    .B(\vga.raw_horizontalPixelCounter[1] ),
    .C(\vga.raw_horizontalPixelCounter[2] ),
    .D(\vga.raw_horizontalPixelCounter[3] ),
    .X(_0310_));
 sky130_fd_sc_hd__o41a_1 _1525_ (.A1(\vga.raw_horizontalPixelCounter[6] ),
    .A2(\vga.raw_horizontalPixelCounter[7] ),
    .A3(\vga.raw_horizontalPixelCounter[8] ),
    .A4(_0310_),
    .B1(_0286_),
    .X(_0311_));
 sky130_fd_sc_hd__and3_4 _1526_ (.A(\vga.configuration[10] ),
    .B(\vga.inVerticalVisibleArea ),
    .C(net605),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_2 _1527_ (.A(\vga.inVerticalVisibleArea ),
    .B(net543),
    .Y(_0313_));
 sky130_fd_sc_hd__nand2_1 _1528_ (.A(\vga.horizontalVisibleAreaCompare[3] ),
    .B(\vga.horizontalCounter[3] ),
    .Y(_0314_));
 sky130_fd_sc_hd__or2_1 _1529_ (.A(\vga.horizontalVisibleAreaCompare[3] ),
    .B(\vga.horizontalCounter[3] ),
    .X(_0315_));
 sky130_fd_sc_hd__nor2_1 _1530_ (.A(\vga.horizontalVisibleAreaCompare[6] ),
    .B(_1338_),
    .Y(_0316_));
 sky130_fd_sc_hd__xor2_1 _1531_ (.A(\vga.horizontalVisibleAreaCompare[10] ),
    .B(\vga.horizontalCounter[10] ),
    .X(_0317_));
 sky130_fd_sc_hd__a22o_1 _1532_ (.A1(\vga.horizontalVisibleAreaCompare[0] ),
    .A2(_1332_),
    .B1(_1339_),
    .B2(\vga.horizontalVisibleAreaCompare[7] ),
    .X(_0318_));
 sky130_fd_sc_hd__xor2_1 _1533_ (.A(\vga.horizontalVisibleAreaCompare[1] ),
    .B(\vga.horizontalCounter[1] ),
    .X(_0319_));
 sky130_fd_sc_hd__a21o_1 _1534_ (.A1(_0314_),
    .A2(_0315_),
    .B1(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__xor2_1 _1535_ (.A(\vga.horizontalVisibleAreaCompare[2] ),
    .B(\vga.horizontalCounter[2] ),
    .X(_0321_));
 sky130_fd_sc_hd__a221o_2 _1536_ (.A1(_1315_),
    .A2(\vga.horizontalCounter[7] ),
    .B1(_1341_),
    .B2(\vga.horizontalVisibleAreaCompare[9] ),
    .C1(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__o22a_1 _1537_ (.A1(\vga.horizontalVisibleAreaCompare[0] ),
    .A2(_1332_),
    .B1(_1341_),
    .B2(\vga.horizontalVisibleAreaCompare[9] ),
    .X(_0323_));
 sky130_fd_sc_hd__or3b_4 _1538_ (.A(_0317_),
    .B(_0318_),
    .C_N(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__xor2_1 _1539_ (.A(\vga.horizontalVisibleAreaCompare[4] ),
    .B(\vga.horizontalCounter[4] ),
    .X(_0325_));
 sky130_fd_sc_hd__a221o_1 _1540_ (.A1(\vga.horizontalVisibleAreaCompare[5] ),
    .A2(_1337_),
    .B1(\vga.horizontalCounter[8] ),
    .B2(_1316_),
    .C1(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nor2_1 _1541_ (.A(\vga.horizontalVisibleAreaCompare[5] ),
    .B(_1337_),
    .Y(_0327_));
 sky130_fd_sc_hd__a22o_1 _1542_ (.A1(\vga.horizontalVisibleAreaCompare[6] ),
    .A2(_1338_),
    .B1(_1340_),
    .B2(\vga.horizontalVisibleAreaCompare[8] ),
    .X(_0328_));
 sky130_fd_sc_hd__or4_2 _1543_ (.A(_0316_),
    .B(_0326_),
    .C(_0327_),
    .D(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__nor4_4 _1544_ (.A(_0320_),
    .B(_0322_),
    .C(_0324_),
    .D(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__xor2_1 _1545_ (.A(\vga.configuration[5] ),
    .B(\vga.raw_verticalPixelStretchCounter[1] ),
    .X(_0331_));
 sky130_fd_sc_hd__or3b_1 _1546_ (.A(\vga.raw_verticalPixelStretchCounter[0] ),
    .B(_0331_),
    .C_N(\vga.configuration[4] ),
    .X(_0332_));
 sky130_fd_sc_hd__and2b_1 _1547_ (.A_N(\vga.configuration[4] ),
    .B(\vga.raw_verticalPixelStretchCounter[0] ),
    .X(_0333_));
 sky130_fd_sc_hd__a21bo_1 _1548_ (.A1(_0331_),
    .A2(_0333_),
    .B1_N(_0332_),
    .X(_0334_));
 sky130_fd_sc_hd__and3_2 _1549_ (.A(\vga.raw_verticalPixelStretchCounter[2] ),
    .B(\vga.raw_verticalPixelStretchCounter[1] ),
    .C(\vga.raw_verticalPixelStretchCounter[0] ),
    .X(_0335_));
 sky130_fd_sc_hd__a21oi_1 _1550_ (.A1(\vga.raw_verticalPixelStretchCounter[1] ),
    .A2(\vga.raw_verticalPixelStretchCounter[0] ),
    .B1(\vga.raw_verticalPixelStretchCounter[2] ),
    .Y(_0336_));
 sky130_fd_sc_hd__nor2_1 _1551_ (.A(_0335_),
    .B(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__xnor2_1 _1552_ (.A(\vga.configuration[6] ),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__xnor2_2 _1553_ (.A(\vga.raw_verticalPixelStretchCounter[3] ),
    .B(_0335_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand2_1 _1554_ (.A(\vga.configuration[7] ),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__or2_1 _1555_ (.A(\vga.configuration[7] ),
    .B(_0339_),
    .X(_0341_));
 sky130_fd_sc_hd__and4_4 _1556_ (.A(_0334_),
    .B(_0338_),
    .C(_0340_),
    .D(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__and2_4 _1557_ (.A(net528),
    .B(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__nand2_4 _1558_ (.A(net528),
    .B(_0342_),
    .Y(_0344_));
 sky130_fd_sc_hd__nor2_2 _1559_ (.A(net532),
    .B(_0343_),
    .Y(_0345_));
 sky130_fd_sc_hd__nand2_2 _1560_ (.A(net576),
    .B(_0344_),
    .Y(_0346_));
 sky130_fd_sc_hd__or4_2 _1561_ (.A(\vga.raw_verticalPixelCounter[7] ),
    .B(\vga.raw_verticalPixelCounter[8] ),
    .C(\vga.raw_verticalPixelCounter[9] ),
    .D(net576),
    .X(_0347_));
 sky130_fd_sc_hd__or4_1 _1562_ (.A(\vga.raw_verticalPixelCounter[3] ),
    .B(\vga.raw_verticalPixelCounter[4] ),
    .C(\vga.raw_verticalPixelCounter[5] ),
    .D(\vga.raw_verticalPixelCounter[6] ),
    .X(_0348_));
 sky130_fd_sc_hd__o41a_2 _1563_ (.A1(\vga.raw_verticalPixelCounter[0] ),
    .A2(\vga.raw_verticalPixelCounter[1] ),
    .A3(_0347_),
    .A4(_0348_),
    .B1(_0346_),
    .X(_0349_));
 sky130_fd_sc_hd__nor2_1 _1564_ (.A(net532),
    .B(_0344_),
    .Y(_0350_));
 sky130_fd_sc_hd__xnor2_4 _1565_ (.A(_1346_),
    .B(_0302_),
    .Y(_0351_));
 sky130_fd_sc_hd__and2_1 _1566_ (.A(_0285_),
    .B(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__and3b_1 _1567_ (.A_N(_0352_),
    .B(\vga.raw_horizontalPixelCounter[4] ),
    .C(_0307_),
    .X(_0353_));
 sky130_fd_sc_hd__xor2_4 _1568_ (.A(\vga.raw_horizontalPixelCounter[3] ),
    .B(_0301_),
    .X(_0354_));
 sky130_fd_sc_hd__or4_1 _1569_ (.A(_0309_),
    .B(_0311_),
    .C(_0349_),
    .D(_0353_),
    .X(_0355_));
 sky130_fd_sc_hd__a31o_2 _1570_ (.A1(\vga.raw_horizontalPixelCounter[5] ),
    .A2(_0307_),
    .A3(_0308_),
    .B1(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__o22a_4 _1571_ (.A1(\vga.raw_horizontalPixelCounter[4] ),
    .A2(_0300_),
    .B1(_0306_),
    .B2(_0352_),
    .X(_0103_));
 sky130_fd_sc_hd__a31o_1 _1572_ (.A1(\vga.raw_verticalPixelCounter[0] ),
    .A2(\vga.raw_verticalPixelCounter[1] ),
    .A3(_0343_),
    .B1(net532),
    .X(_0357_));
 sky130_fd_sc_hd__a21oi_2 _1573_ (.A1(net595),
    .A2(\vga.raw_horizontalPixelCounter[1] ),
    .B1(\vga.raw_horizontalPixelCounter[2] ),
    .Y(_0358_));
 sky130_fd_sc_hd__nor2_4 _1574_ (.A(_0301_),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__and4_1 _1575_ (.A(\vga.raw_verticalPixelCounter[0] ),
    .B(\vga.raw_verticalPixelCounter[1] ),
    .C(\vga.raw_verticalPixelCounter[2] ),
    .D(_0343_),
    .X(_0360_));
 sky130_fd_sc_hd__and2_1 _1576_ (.A(\vga.raw_verticalPixelCounter[3] ),
    .B(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__and3_2 _1577_ (.A(\vga.raw_verticalPixelCounter[3] ),
    .B(\vga.raw_verticalPixelCounter[4] ),
    .C(_0360_),
    .X(_0362_));
 sky130_fd_sc_hd__and2_1 _1578_ (.A(\vga.raw_verticalPixelCounter[5] ),
    .B(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__a21oi_1 _1579_ (.A1(\vga.raw_verticalPixelCounter[6] ),
    .A2(_0363_),
    .B1(net532),
    .Y(_0364_));
 sky130_fd_sc_hd__nor2_1 _1580_ (.A(net532),
    .B(_0362_),
    .Y(_0365_));
 sky130_fd_sc_hd__a22o_4 _1581_ (.A1(\vga.raw_horizontalPixelCounter[2] ),
    .A2(_0306_),
    .B1(_0309_),
    .B2(_0359_),
    .X(_0101_));
 sky130_fd_sc_hd__a22o_2 _1582_ (.A1(\vga.raw_horizontalPixelCounter[3] ),
    .A2(_0306_),
    .B1(_0309_),
    .B2(_0354_),
    .X(_0102_));
 sky130_fd_sc_hd__a221o_2 _1583_ (.A1(_1346_),
    .A2(_0103_),
    .B1(_0357_),
    .B2(\vga.raw_verticalPixelCounter[2] ),
    .C1(_0356_),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _1584_ (.A(net539),
    .B(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__inv_2 _1585_ (.A(_0367_),
    .Y(_0157_));
 sky130_fd_sc_hd__and2_4 _1586_ (.A(\vga.raw_horizontalPixelCounter[6] ),
    .B(_0303_),
    .X(_0368_));
 sky130_fd_sc_hd__nand2_2 _1587_ (.A(\vga.raw_horizontalPixelCounter[7] ),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__xnor2_4 _1588_ (.A(\vga.raw_horizontalPixelCounter[8] ),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__a22o_4 _1589_ (.A1(\vga.raw_horizontalPixelCounter[8] ),
    .A2(_0306_),
    .B1(_0309_),
    .B2(_0370_),
    .X(_0107_));
 sky130_fd_sc_hd__xnor2_1 _1590_ (.A(\vga.raw_directPixelCounterVertical[8] ),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__xor2_4 _1591_ (.A(\vga.raw_horizontalPixelCounter[7] ),
    .B(_0368_),
    .X(_0372_));
 sky130_fd_sc_hd__nand2_1 _1592_ (.A(\vga.raw_directPixelCounterVertical[7] ),
    .B(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__or2_1 _1593_ (.A(\vga.raw_directPixelCounterVertical[7] ),
    .B(_0372_),
    .X(_0374_));
 sky130_fd_sc_hd__nor2_1 _1594_ (.A(\vga.raw_horizontalPixelCounter[6] ),
    .B(_0303_),
    .Y(_0375_));
 sky130_fd_sc_hd__nor2_2 _1595_ (.A(_0368_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__and2_1 _1596_ (.A(\vga.raw_directPixelCounterVertical[6] ),
    .B(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__nand2_1 _1597_ (.A(\vga.raw_directPixelCounterVertical[6] ),
    .B(_0376_),
    .Y(_0378_));
 sky130_fd_sc_hd__nor2_1 _1598_ (.A(\vga.raw_directPixelCounterVertical[6] ),
    .B(_0376_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _1599_ (.A(\vga.raw_directPixelCounterVertical[4] ),
    .B(_0351_),
    .Y(_0380_));
 sky130_fd_sc_hd__xnor2_2 _1600_ (.A(\vga.raw_directPixelCounterVertical[4] ),
    .B(_0351_),
    .Y(_0381_));
 sky130_fd_sc_hd__and2_1 _1601_ (.A(\vga.raw_directPixelCounterVertical[3] ),
    .B(_0354_),
    .X(_0382_));
 sky130_fd_sc_hd__nand2_1 _1602_ (.A(\vga.raw_directPixelCounterVertical[3] ),
    .B(_0354_),
    .Y(_0383_));
 sky130_fd_sc_hd__nor2_2 _1603_ (.A(\vga.raw_directPixelCounterVertical[3] ),
    .B(_0354_),
    .Y(_0384_));
 sky130_fd_sc_hd__nand2_1 _1604_ (.A(\vga.raw_directPixelCounterVertical[2] ),
    .B(_0359_),
    .Y(_0385_));
 sky130_fd_sc_hd__xnor2_2 _1605_ (.A(\vga.raw_directPixelCounterVertical[2] ),
    .B(_0359_),
    .Y(_0386_));
 sky130_fd_sc_hd__xor2_4 _1606_ (.A(\vga.raw_horizontalPixelCounter[0] ),
    .B(\vga.raw_horizontalPixelCounter[1] ),
    .X(_0387_));
 sky130_fd_sc_hd__xnor2_1 _1607_ (.A(net595),
    .B(\vga.raw_horizontalPixelCounter[1] ),
    .Y(_0388_));
 sky130_fd_sc_hd__nand2_1 _1608_ (.A(\vga.raw_directPixelCounterVertical[1] ),
    .B(_0387_),
    .Y(_0389_));
 sky130_fd_sc_hd__xnor2_1 _1609_ (.A(\vga.raw_directPixelCounterVertical[1] ),
    .B(_0387_),
    .Y(_0390_));
 sky130_fd_sc_hd__or3_1 _1610_ (.A(net595),
    .B(_1350_),
    .C(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__o31a_2 _1611_ (.A1(net595),
    .A2(_1350_),
    .A3(_0390_),
    .B1(_0389_),
    .X(_0392_));
 sky130_fd_sc_hd__o21a_1 _1612_ (.A1(_0386_),
    .A2(_0392_),
    .B1(_0385_),
    .X(_0393_));
 sky130_fd_sc_hd__o211a_1 _1613_ (.A1(_0386_),
    .A2(_0392_),
    .B1(_0383_),
    .C1(_0385_),
    .X(_0394_));
 sky130_fd_sc_hd__nor2_1 _1614_ (.A(_0384_),
    .B(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__o31a_1 _1615_ (.A1(_0381_),
    .A2(_0384_),
    .A3(_0394_),
    .B1(_0380_),
    .X(_0396_));
 sky130_fd_sc_hd__o211a_1 _1616_ (.A1(\vga.raw_directPixelCounterVertical[5] ),
    .A2(_0305_),
    .B1(_0351_),
    .C1(\vga.raw_directPixelCounterVertical[4] ),
    .X(_0397_));
 sky130_fd_sc_hd__a21oi_1 _1617_ (.A1(\vga.raw_directPixelCounterVertical[5] ),
    .A2(_0305_),
    .B1(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__xnor2_2 _1618_ (.A(\vga.raw_directPixelCounterVertical[5] ),
    .B(_0305_),
    .Y(_0399_));
 sky130_fd_sc_hd__or4_1 _1619_ (.A(_0381_),
    .B(_0384_),
    .C(_0394_),
    .D(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__nand2_1 _1620_ (.A(_0398_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__a31o_2 _1621_ (.A1(_0378_),
    .A2(_0398_),
    .A3(_0400_),
    .B1(_0379_),
    .X(_0402_));
 sky130_fd_sc_hd__a21boi_2 _1622_ (.A1(_0373_),
    .A2(_0402_),
    .B1_N(_0374_),
    .Y(_0403_));
 sky130_fd_sc_hd__xnor2_1 _1623_ (.A(_0371_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__or2_1 _1624_ (.A(\vga.raw_directPixelCounterVertical[8] ),
    .B(_0343_),
    .X(_0405_));
 sky130_fd_sc_hd__o211a_2 _1625_ (.A1(_0344_),
    .A2(_0404_),
    .B1(_0405_),
    .C1(_0312_),
    .X(_0072_));
 sky130_fd_sc_hd__and2_2 _1626_ (.A(_0107_),
    .B(_0072_),
    .X(_0406_));
 sky130_fd_sc_hd__xor2_2 _1627_ (.A(_0107_),
    .B(_0072_),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_2 _1628_ (.A1(\vga.raw_horizontalPixelCounter[7] ),
    .A2(_0306_),
    .B1(_0309_),
    .B2(_0372_),
    .X(_0106_));
 sky130_fd_sc_hd__nand2_1 _1629_ (.A(_0373_),
    .B(_0374_),
    .Y(_0408_));
 sky130_fd_sc_hd__nor2_1 _1630_ (.A(_0402_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__a21bo_1 _1631_ (.A1(_0402_),
    .A2(_0408_),
    .B1_N(_0350_),
    .X(_0410_));
 sky130_fd_sc_hd__o2bb2a_1 _1632_ (.A1_N(\vga.raw_directPixelCounterVertical[7] ),
    .A2_N(_0345_),
    .B1(_0409_),
    .B2(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__inv_2 _1633_ (.A(_0411_),
    .Y(_0071_));
 sky130_fd_sc_hd__or2_2 _1634_ (.A(_0106_),
    .B(_0071_),
    .X(_0412_));
 sky130_fd_sc_hd__inv_2 _1635_ (.A(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__and2_2 _1636_ (.A(_0106_),
    .B(_0071_),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_4 _1637_ (.A1(\vga.raw_horizontalPixelCounter[6] ),
    .A2(_0306_),
    .B1(_0309_),
    .B2(_0376_),
    .X(_0105_));
 sky130_fd_sc_hd__nor2_1 _1638_ (.A(_0377_),
    .B(_0379_),
    .Y(_0415_));
 sky130_fd_sc_hd__xnor2_2 _1639_ (.A(_0401_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__o21ai_2 _1640_ (.A1(\vga.raw_directPixelCounterVertical[6] ),
    .A2(_0343_),
    .B1(_0312_),
    .Y(_0417_));
 sky130_fd_sc_hd__a21oi_4 _1641_ (.A1(_0343_),
    .A2(_0416_),
    .B1(_0417_),
    .Y(_0070_));
 sky130_fd_sc_hd__and2_2 _1642_ (.A(_0105_),
    .B(_0070_),
    .X(_0418_));
 sky130_fd_sc_hd__xor2_2 _1643_ (.A(_0105_),
    .B(_0070_),
    .X(_0419_));
 sky130_fd_sc_hd__a2bb2oi_4 _1644_ (.A1_N(\vga.raw_horizontalPixelCounter[5] ),
    .A2_N(_0300_),
    .B1(_0307_),
    .B2(_0308_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand2_1 _1645_ (.A(_0396_),
    .B(_0399_),
    .Y(_0420_));
 sky130_fd_sc_hd__or2_1 _1646_ (.A(_0396_),
    .B(_0399_),
    .X(_0421_));
 sky130_fd_sc_hd__o21ai_1 _1647_ (.A1(_1348_),
    .A2(_0342_),
    .B1(net528),
    .Y(_0422_));
 sky130_fd_sc_hd__a31o_1 _1648_ (.A1(_0342_),
    .A2(_0420_),
    .A3(_0421_),
    .B1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__o211a_1 _1649_ (.A1(\vga.raw_directPixelCounterVertical[5] ),
    .A2(net529),
    .B1(_0423_),
    .C1(_0312_),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _1650_ (.A(_0104_),
    .B(_0069_),
    .X(_0424_));
 sky130_fd_sc_hd__or2_2 _1651_ (.A(_0104_),
    .B(_0069_),
    .X(_0425_));
 sky130_fd_sc_hd__xnor2_1 _1652_ (.A(_0381_),
    .B(_0395_),
    .Y(_0426_));
 sky130_fd_sc_hd__a22o_2 _1653_ (.A1(\vga.raw_directPixelCounterVertical[4] ),
    .A2(_0345_),
    .B1(_0350_),
    .B2(_0426_),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _1654_ (.A(_0103_),
    .B(_0068_),
    .X(_0427_));
 sky130_fd_sc_hd__xor2_1 _1655_ (.A(_0103_),
    .B(_0068_),
    .X(_0428_));
 sky130_fd_sc_hd__or3_1 _1656_ (.A(_0382_),
    .B(_0384_),
    .C(_0393_),
    .X(_0429_));
 sky130_fd_sc_hd__o21ai_1 _1657_ (.A1(_0382_),
    .A2(_0384_),
    .B1(_0393_),
    .Y(_0430_));
 sky130_fd_sc_hd__a32o_1 _1658_ (.A1(_0350_),
    .A2(_0429_),
    .A3(_0430_),
    .B1(_0345_),
    .B2(\vga.raw_directPixelCounterVertical[3] ),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _1659_ (.A(_0102_),
    .B(_0067_),
    .X(_0431_));
 sky130_fd_sc_hd__or2_1 _1660_ (.A(_0102_),
    .B(_0067_),
    .X(_0432_));
 sky130_fd_sc_hd__xor2_1 _1661_ (.A(_0386_),
    .B(_0392_),
    .X(_0433_));
 sky130_fd_sc_hd__a21o_1 _1662_ (.A1(net529),
    .A2(_0342_),
    .B1(\vga.raw_directPixelCounterVertical[2] ),
    .X(_0434_));
 sky130_fd_sc_hd__o211a_2 _1663_ (.A1(_0344_),
    .A2(_0433_),
    .B1(_0434_),
    .C1(net576),
    .X(_0066_));
 sky130_fd_sc_hd__nand2_2 _1664_ (.A(_0101_),
    .B(_0066_),
    .Y(_0435_));
 sky130_fd_sc_hd__or2_1 _1665_ (.A(_0101_),
    .B(_0066_),
    .X(_0436_));
 sky130_fd_sc_hd__a211oi_2 _1666_ (.A1(net528),
    .A2(_0342_),
    .B1(_1349_),
    .C1(_0313_),
    .Y(_0437_));
 sky130_fd_sc_hd__o21ai_1 _1667_ (.A1(net595),
    .A2(_1350_),
    .B1(_0390_),
    .Y(_0438_));
 sky130_fd_sc_hd__and2_1 _1668_ (.A(_0391_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__and4_1 _1669_ (.A(net576),
    .B(net528),
    .C(_0342_),
    .D(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__or2_1 _1670_ (.A(_0437_),
    .B(_0440_),
    .X(_0065_));
 sky130_fd_sc_hd__a31o_1 _1671_ (.A1(_0287_),
    .A2(_0290_),
    .A3(_0298_),
    .B1(\vga.raw_horizontalPixelCounter[1] ),
    .X(_0441_));
 sky130_fd_sc_hd__and4_1 _1672_ (.A(_0287_),
    .B(_0290_),
    .C(_0298_),
    .D(_0388_),
    .X(_0442_));
 sky130_fd_sc_hd__and3b_4 _1673_ (.A_N(_0442_),
    .B(_0285_),
    .C(_0441_),
    .X(_0100_));
 sky130_fd_sc_hd__o21a_1 _1674_ (.A1(_0437_),
    .A2(_0440_),
    .B1(_0100_),
    .X(_0443_));
 sky130_fd_sc_hd__a31o_1 _1675_ (.A1(_1345_),
    .A2(net528),
    .A3(_0342_),
    .B1(\vga.raw_directPixelCounterVertical[0] ),
    .X(_0444_));
 sky130_fd_sc_hd__o311a_4 _1676_ (.A1(net595),
    .A2(_1350_),
    .A3(_0344_),
    .B1(_0444_),
    .C1(net576),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_8 _1677_ (.A0(_0306_),
    .A1(_0309_),
    .S(_1345_),
    .X(_0099_));
 sky130_fd_sc_hd__nand2_1 _1678_ (.A(_0064_),
    .B(_0099_),
    .Y(_0445_));
 sky130_fd_sc_hd__or3_4 _1679_ (.A(_0437_),
    .B(_0440_),
    .C(_0100_),
    .X(_0446_));
 sky130_fd_sc_hd__nand2b_1 _1680_ (.A_N(_0443_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__a31oi_4 _1681_ (.A1(_0064_),
    .A2(_0099_),
    .A3(_0446_),
    .B1(_0443_),
    .Y(_0448_));
 sky130_fd_sc_hd__a21boi_4 _1682_ (.A1(_0435_),
    .A2(_0448_),
    .B1_N(_0436_),
    .Y(_0449_));
 sky130_fd_sc_hd__o21a_1 _1683_ (.A1(_0431_),
    .A2(_0449_),
    .B1(_0432_),
    .X(_0450_));
 sky130_fd_sc_hd__o211a_2 _1684_ (.A1(_0431_),
    .A2(_0449_),
    .B1(_0432_),
    .C1(_0428_),
    .X(_0451_));
 sky130_fd_sc_hd__or2_2 _1685_ (.A(_0427_),
    .B(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__o311a_4 _1686_ (.A1(_0424_),
    .A2(_0427_),
    .A3(_0451_),
    .B1(_0425_),
    .C1(_0419_),
    .X(_0453_));
 sky130_fd_sc_hd__o31a_1 _1687_ (.A1(_0414_),
    .A2(_0418_),
    .A3(_0453_),
    .B1(_0412_),
    .X(_0454_));
 sky130_fd_sc_hd__o311a_4 _1688_ (.A1(_0414_),
    .A2(_0418_),
    .A3(_0453_),
    .B1(_0412_),
    .C1(_0407_),
    .X(_0455_));
 sky130_fd_sc_hd__a21o_1 _1689_ (.A1(\vga.raw_directPixelCounterVertical[8] ),
    .A2(_0370_),
    .B1(_0403_),
    .X(_0456_));
 sky130_fd_sc_hd__o211ai_4 _1690_ (.A1(\vga.raw_directPixelCounterVertical[8] ),
    .A2(_0370_),
    .B1(_0456_),
    .C1(_0343_),
    .Y(_0457_));
 sky130_fd_sc_hd__or2_1 _1691_ (.A(_1347_),
    .B(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__a21oi_1 _1692_ (.A1(_1347_),
    .A2(_0457_),
    .B1(net532),
    .Y(_0459_));
 sky130_fd_sc_hd__and2_2 _1693_ (.A(_0458_),
    .B(_0459_),
    .X(_0073_));
 sky130_fd_sc_hd__o21ai_4 _1694_ (.A1(_0406_),
    .A2(_0455_),
    .B1(_0073_),
    .Y(_0460_));
 sky130_fd_sc_hd__xor2_1 _1695_ (.A(\vga.raw_directPixelCounterVertical[10] ),
    .B(_0458_),
    .X(_0461_));
 sky130_fd_sc_hd__o211a_1 _1696_ (.A1(_0406_),
    .A2(_0455_),
    .B1(_0073_),
    .C1(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__and2b_2 _1697_ (.A_N(\vga.configuration[9] ),
    .B(\vga.configuration[8] ),
    .X(_0463_));
 sky130_fd_sc_hd__nand2b_4 _1698_ (.A_N(\vga.configuration[9] ),
    .B(\vga.configuration[8] ),
    .Y(_0464_));
 sky130_fd_sc_hd__nor2_1 _1699_ (.A(net532),
    .B(_0461_),
    .Y(_0074_));
 sky130_fd_sc_hd__a211oi_2 _1700_ (.A1(_0460_),
    .A2(_0074_),
    .B1(_0464_),
    .C1(_0462_),
    .Y(_0465_));
 sky130_fd_sc_hd__a211o_1 _1701_ (.A1(_0460_),
    .A2(_0074_),
    .B1(_0464_),
    .C1(_0462_),
    .X(_0466_));
 sky130_fd_sc_hd__o21a_1 _1702_ (.A1(\vga.raw_verticalPixelCounter[6] ),
    .A2(_0363_),
    .B1(_0364_),
    .X(_0092_));
 sky130_fd_sc_hd__nor2_1 _1703_ (.A(net575),
    .B(_0092_),
    .Y(_0467_));
 sky130_fd_sc_hd__or2_1 _1704_ (.A(net575),
    .B(_0092_),
    .X(_0468_));
 sky130_fd_sc_hd__nand2_2 _1705_ (.A(net493),
    .B(net501),
    .Y(_0469_));
 sky130_fd_sc_hd__nor2_1 _1706_ (.A(net532),
    .B(_0363_),
    .Y(_0470_));
 sky130_fd_sc_hd__o21a_1 _1707_ (.A1(\vga.raw_verticalPixelCounter[5] ),
    .A2(_0362_),
    .B1(_0470_),
    .X(_0091_));
 sky130_fd_sc_hd__o31a_2 _1708_ (.A1(_0406_),
    .A2(_0455_),
    .A3(_0073_),
    .B1(net575),
    .X(_0471_));
 sky130_fd_sc_hd__and2_2 _1709_ (.A(_0464_),
    .B(_0091_),
    .X(_0472_));
 sky130_fd_sc_hd__a21o_1 _1710_ (.A1(_0460_),
    .A2(_0471_),
    .B1(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__a21oi_4 _1711_ (.A1(_0460_),
    .A2(_0471_),
    .B1(_0472_),
    .Y(_0474_));
 sky130_fd_sc_hd__a21o_1 _1712_ (.A1(net493),
    .A2(net501),
    .B1(net492),
    .X(_0475_));
 sky130_fd_sc_hd__or2_4 _1713_ (.A(_0367_),
    .B(net477),
    .X(net333));
 sky130_fd_sc_hd__nand2_1 _1714_ (.A(_0366_),
    .B(net492),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2b_4 _1715_ (.A_N(_0476_),
    .B(_0469_),
    .Y(net334));
 sky130_fd_sc_hd__or3_2 _1716_ (.A(_0367_),
    .B(_0469_),
    .C(net492),
    .X(net394));
 sky130_fd_sc_hd__or2_1 _1717_ (.A(_0469_),
    .B(_0476_),
    .X(net395));
 sky130_fd_sc_hd__nand2_2 _1718_ (.A(_0064_),
    .B(net575),
    .Y(_0477_));
 sky130_fd_sc_hd__xnor2_4 _1719_ (.A(_0099_),
    .B(_0477_),
    .Y(net320));
 sky130_fd_sc_hd__xor2_1 _1720_ (.A(_0445_),
    .B(_0447_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_8 _1721_ (.A0(_0100_),
    .A1(_0478_),
    .S(net575),
    .X(net321));
 sky130_fd_sc_hd__nand2_1 _1722_ (.A(_0435_),
    .B(_0436_),
    .Y(_0479_));
 sky130_fd_sc_hd__xor2_1 _1723_ (.A(_0448_),
    .B(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_8 _1724_ (.A0(_0101_),
    .A1(_0480_),
    .S(net575),
    .X(net322));
 sky130_fd_sc_hd__nand2b_1 _1725_ (.A_N(_0431_),
    .B(_0432_),
    .Y(_0481_));
 sky130_fd_sc_hd__xnor2_1 _1726_ (.A(_0449_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__mux2_8 _1727_ (.A0(_0102_),
    .A1(_0482_),
    .S(net575),
    .X(net323));
 sky130_fd_sc_hd__o21ai_1 _1728_ (.A1(\vga.raw_verticalPixelCounter[0] ),
    .A2(_0343_),
    .B1(net576),
    .Y(_0483_));
 sky130_fd_sc_hd__a21oi_2 _1729_ (.A1(\vga.raw_verticalPixelCounter[0] ),
    .A2(_0343_),
    .B1(_0483_),
    .Y(_0086_));
 sky130_fd_sc_hd__o21ai_1 _1730_ (.A1(_0428_),
    .A2(_0450_),
    .B1(net575),
    .Y(_0484_));
 sky130_fd_sc_hd__a2bb2o_4 _1731_ (.A1_N(_0451_),
    .A2_N(_0484_),
    .B1(_0464_),
    .B2(_0086_),
    .X(net324));
 sky130_fd_sc_hd__and2b_1 _1732_ (.A_N(_0424_),
    .B(_0425_),
    .X(_0485_));
 sky130_fd_sc_hd__xor2_2 _1733_ (.A(_0452_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__a31o_1 _1734_ (.A1(\vga.raw_verticalPixelCounter[0] ),
    .A2(net528),
    .A3(_0342_),
    .B1(\vga.raw_verticalPixelCounter[1] ),
    .X(_0487_));
 sky130_fd_sc_hd__and2b_1 _1735_ (.A_N(_0357_),
    .B(_0487_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_8 _1736_ (.A0(_0486_),
    .A1(_0087_),
    .S(_0464_),
    .X(net325));
 sky130_fd_sc_hd__a211oi_1 _1737_ (.A1(_0425_),
    .A2(_0452_),
    .B1(_0419_),
    .C1(_0424_),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2_1 _1738_ (.A(_0453_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__a31o_1 _1739_ (.A1(\vga.raw_verticalPixelCounter[0] ),
    .A2(\vga.raw_verticalPixelCounter[1] ),
    .A3(_0343_),
    .B1(\vga.raw_verticalPixelCounter[2] ),
    .X(_0490_));
 sky130_fd_sc_hd__and3b_1 _1740_ (.A_N(_0360_),
    .B(_0490_),
    .C(net576),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_8 _1741_ (.A0(_0489_),
    .A1(_0088_),
    .S(_0464_),
    .X(net326));
 sky130_fd_sc_hd__o22ai_4 _1742_ (.A1(_0413_),
    .A2(_0414_),
    .B1(_0418_),
    .B2(_0453_),
    .Y(_0491_));
 sky130_fd_sc_hd__o41a_1 _1743_ (.A1(_0413_),
    .A2(_0414_),
    .A3(_0418_),
    .A4(_0453_),
    .B1(net575),
    .X(_0492_));
 sky130_fd_sc_hd__o21ai_1 _1744_ (.A1(\vga.raw_verticalPixelCounter[3] ),
    .A2(_0360_),
    .B1(net576),
    .Y(_0493_));
 sky130_fd_sc_hd__nor2_1 _1745_ (.A(_0361_),
    .B(_0493_),
    .Y(_0089_));
 sky130_fd_sc_hd__o2bb2a_4 _1746_ (.A1_N(_0491_),
    .A2_N(_0492_),
    .B1(_0089_),
    .B2(_0463_),
    .X(net327));
 sky130_fd_sc_hd__o21a_1 _1747_ (.A1(\vga.raw_verticalPixelCounter[4] ),
    .A2(_0361_),
    .B1(_0365_),
    .X(_0090_));
 sky130_fd_sc_hd__o21ai_1 _1748_ (.A1(_0407_),
    .A2(_0454_),
    .B1(net575),
    .Y(_0494_));
 sky130_fd_sc_hd__a2bb2o_4 _1749_ (.A1_N(_0455_),
    .A2_N(_0494_),
    .B1(_0464_),
    .B2(_0090_),
    .X(net328));
 sky130_fd_sc_hd__nor3b_4 _1750_ (.A(\vga.raw_subPixelCounter_buffered[0] ),
    .B(\vga.raw_subPixelCounter_buffered[2] ),
    .C_N(\vga.raw_subPixelCounter_buffered[1] ),
    .Y(_0495_));
 sky130_fd_sc_hd__nor3b_4 _1751_ (.A(\vga.raw_subPixelCounter_buffered[0] ),
    .B(\vga.raw_subPixelCounter_buffered[1] ),
    .C_N(\vga.raw_subPixelCounter_buffered[2] ),
    .Y(_0496_));
 sky130_fd_sc_hd__nor3b_4 _1752_ (.A(\vga.raw_subPixelCounter_buffered[1] ),
    .B(\vga.raw_subPixelCounter_buffered[2] ),
    .C_N(\vga.raw_subPixelCounter_buffered[0] ),
    .Y(_0497_));
 sky130_fd_sc_hd__and3b_4 _1753_ (.A_N(\vga.raw_subPixelCounter_buffered[2] ),
    .B(\vga.raw_subPixelCounter_buffered[1] ),
    .C(\vga.raw_subPixelCounter_buffered[0] ),
    .X(_0498_));
 sky130_fd_sc_hd__nor4_4 _1754_ (.A(_0495_),
    .B(_0496_),
    .C(_0497_),
    .D(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__or4_4 _1755_ (.A(_0495_),
    .B(_0496_),
    .C(_0497_),
    .D(_0498_),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_2 _1756_ (.A1(\vga.currentPixelData[28] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(\vga.currentPixelData[22] ),
    .X(_0501_));
 sky130_fd_sc_hd__a22o_1 _1757_ (.A1(\vga.currentPixelData[16] ),
    .A2(_0495_),
    .B1(_0497_),
    .B2(\vga.currentPixelData[10] ),
    .X(_0502_));
 sky130_fd_sc_hd__or3_2 _1758_ (.A(_0499_),
    .B(_0501_),
    .C(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__o211a_1 _1759_ (.A1(\vga.currentPixelData[4] ),
    .A2(_0500_),
    .B1(_0503_),
    .C1(_0284_),
    .X(net433));
 sky130_fd_sc_hd__a22o_1 _1760_ (.A1(\vga.currentPixelData[29] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(\vga.currentPixelData[23] ),
    .X(_0504_));
 sky130_fd_sc_hd__a22o_1 _1761_ (.A1(\vga.currentPixelData[17] ),
    .A2(_0495_),
    .B1(_0497_),
    .B2(\vga.currentPixelData[11] ),
    .X(_0505_));
 sky130_fd_sc_hd__or3_4 _1762_ (.A(_0499_),
    .B(_0504_),
    .C(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__o211a_1 _1763_ (.A1(\vga.currentPixelData[5] ),
    .A2(_0500_),
    .B1(_0506_),
    .C1(_0284_),
    .X(net434));
 sky130_fd_sc_hd__a22o_1 _1764_ (.A1(\vga.currentPixelData[26] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(\vga.currentPixelData[20] ),
    .X(_0507_));
 sky130_fd_sc_hd__a22o_1 _1765_ (.A1(\vga.currentPixelData[14] ),
    .A2(_0495_),
    .B1(_0497_),
    .B2(\vga.currentPixelData[8] ),
    .X(_0508_));
 sky130_fd_sc_hd__or3_2 _1766_ (.A(_0499_),
    .B(_0507_),
    .C(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__o211a_1 _1767_ (.A1(\vga.currentPixelData[2] ),
    .A2(_0500_),
    .B1(_0509_),
    .C1(_0284_),
    .X(net435));
 sky130_fd_sc_hd__a22o_2 _1768_ (.A1(\vga.currentPixelData[27] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(\vga.currentPixelData[21] ),
    .X(_0510_));
 sky130_fd_sc_hd__a22o_1 _1769_ (.A1(\vga.currentPixelData[15] ),
    .A2(_0495_),
    .B1(_0497_),
    .B2(\vga.currentPixelData[9] ),
    .X(_0511_));
 sky130_fd_sc_hd__or3_2 _1770_ (.A(_0499_),
    .B(_0510_),
    .C(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__o211a_1 _1771_ (.A1(\vga.currentPixelData[3] ),
    .A2(_0500_),
    .B1(_0512_),
    .C1(_0284_),
    .X(net436));
 sky130_fd_sc_hd__a22o_2 _1772_ (.A1(\vga.currentPixelData[24] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(\vga.currentPixelData[18] ),
    .X(_0513_));
 sky130_fd_sc_hd__a22o_1 _1773_ (.A1(\vga.currentPixelData[12] ),
    .A2(_0495_),
    .B1(_0497_),
    .B2(\vga.currentPixelData[6] ),
    .X(_0514_));
 sky130_fd_sc_hd__or3_1 _1774_ (.A(_0499_),
    .B(_0513_),
    .C(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__o211a_1 _1775_ (.A1(\vga.currentPixelData[0] ),
    .A2(_0500_),
    .B1(_0515_),
    .C1(_0284_),
    .X(net438));
 sky130_fd_sc_hd__a22o_2 _1776_ (.A1(\vga.currentPixelData[25] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(\vga.currentPixelData[19] ),
    .X(_0516_));
 sky130_fd_sc_hd__a22o_1 _1777_ (.A1(\vga.currentPixelData[13] ),
    .A2(_0495_),
    .B1(_0497_),
    .B2(\vga.currentPixelData[7] ),
    .X(_0517_));
 sky130_fd_sc_hd__or3_1 _1778_ (.A(_0499_),
    .B(_0516_),
    .C(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__o211a_1 _1779_ (.A1(\vga.currentPixelData[1] ),
    .A2(_0500_),
    .B1(_0518_),
    .C1(_0284_),
    .X(net439));
 sky130_fd_sc_hd__nor2_8 _1780_ (.A(\videoMemory.wbReadReady ),
    .B(net531),
    .Y(_0519_));
 sky130_fd_sc_hd__nor2_8 _1781_ (.A(net578),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__or2_1 _1782_ (.A(net578),
    .B(_0519_),
    .X(_0521_));
 sky130_fd_sc_hd__nand2_1 _1783_ (.A(\wbPeripheralBusInterface.currentAddress[23] ),
    .B(net581),
    .Y(_0522_));
 sky130_fd_sc_hd__or4_2 _1784_ (.A(\wbPeripheralBusInterface.currentAddress[12] ),
    .B(_0269_),
    .C(_0271_),
    .D(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__a2111oi_4 _1785_ (.A1(\wbPeripheralBusInterface.currentAddress[11] ),
    .A2(net581),
    .B1(net319),
    .C1(_0270_),
    .D1(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__nor4_4 _1786_ (.A(net315),
    .B(net316),
    .C(net317),
    .D(net318),
    .Y(_0525_));
 sky130_fd_sc_hd__and4_4 _1787_ (.A(_1356_),
    .B(_1357_),
    .C(_0524_),
    .D(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__and3_2 _1788_ (.A(_1355_),
    .B(_0267_),
    .C(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__and2_2 _1789_ (.A(net579),
    .B(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__nand2_1 _1790_ (.A(net579),
    .B(_0527_),
    .Y(_0529_));
 sky130_fd_sc_hd__a21o_1 _1791_ (.A1(\vga.configuration[0] ),
    .A2(net565),
    .B1(net521),
    .X(_0530_));
 sky130_fd_sc_hd__a221o_2 _1792_ (.A1(net26),
    .A2(net556),
    .B1(net545),
    .B2(net150),
    .C1(net563),
    .X(_0531_));
 sky130_fd_sc_hd__a21o_4 _1793_ (.A1(net125),
    .A2(net548),
    .B1(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__and3_4 _1794_ (.A(\videoMemory.wbReadReady ),
    .B(net599),
    .C(net580),
    .X(_0533_));
 sky130_fd_sc_hd__o211a_2 _1795_ (.A1(net1),
    .A2(net559),
    .B1(_0532_),
    .C1(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__nor2_2 _1796_ (.A(\wbPeripheralBusInterface.currentAddress[5] ),
    .B(_1355_),
    .Y(_0535_));
 sky130_fd_sc_hd__and2_4 _1797_ (.A(_0526_),
    .B(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__and3_2 _1798_ (.A(net579),
    .B(_0526_),
    .C(_0535_),
    .X(_0537_));
 sky130_fd_sc_hd__nand2_2 _1799_ (.A(net579),
    .B(_0536_),
    .Y(_0538_));
 sky130_fd_sc_hd__and2_1 _1800_ (.A(_0524_),
    .B(_0535_),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_2 _1801_ (.A(_0524_),
    .B(_0535_),
    .Y(_0540_));
 sky130_fd_sc_hd__or3b_4 _1802_ (.A(\wbPeripheralBusInterface.currentAddress[3] ),
    .B(_1356_),
    .C_N(_0525_),
    .X(_0541_));
 sky130_fd_sc_hd__nor2_4 _1803_ (.A(_0540_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__and2_2 _1804_ (.A(net579),
    .B(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__nand2_2 _1805_ (.A(_0275_),
    .B(_0542_),
    .Y(_0544_));
 sky130_fd_sc_hd__or3b_4 _1806_ (.A(\wbPeripheralBusInterface.currentAddress[2] ),
    .B(_1357_),
    .C_N(_0525_),
    .X(_0545_));
 sky130_fd_sc_hd__nor2_2 _1807_ (.A(_0540_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__and2_2 _1808_ (.A(net579),
    .B(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__nand2_2 _1809_ (.A(net579),
    .B(_0546_),
    .Y(_0548_));
 sky130_fd_sc_hd__and3_1 _1810_ (.A(\wbPeripheralBusInterface.currentAddress[3] ),
    .B(net311),
    .C(_0525_),
    .X(_0549_));
 sky130_fd_sc_hd__or3b_4 _1811_ (.A(\wbPeripheralBusInterface.currentAddress[4] ),
    .B(_0267_),
    .C_N(_0524_),
    .X(_0550_));
 sky130_fd_sc_hd__or4bb_4 _1812_ (.A(\wbPeripheralBusInterface.currentAddress[4] ),
    .B(_0267_),
    .C_N(_0524_),
    .D_N(_0549_),
    .X(_0551_));
 sky130_fd_sc_hd__nor2_8 _1813_ (.A(net577),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__a211o_1 _1814_ (.A1(\vga.verticalWholeLineCompare[0] ),
    .A2(net570),
    .B1(net578),
    .C1(_0551_),
    .X(_0553_));
 sky130_fd_sc_hd__nor3_4 _1815_ (.A(net577),
    .B(_0545_),
    .C(_0550_),
    .Y(_0554_));
 sky130_fd_sc_hd__or3_4 _1816_ (.A(net577),
    .B(_0545_),
    .C(_0550_),
    .X(_0555_));
 sky130_fd_sc_hd__or2_4 _1817_ (.A(_0541_),
    .B(_0550_),
    .X(_0556_));
 sky130_fd_sc_hd__nor2_2 _1818_ (.A(net577),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__or2_2 _1819_ (.A(net578),
    .B(_0556_),
    .X(_0558_));
 sky130_fd_sc_hd__or3b_4 _1820_ (.A(\wbPeripheralBusInterface.currentAddress[4] ),
    .B(_0267_),
    .C_N(_0526_),
    .X(_0559_));
 sky130_fd_sc_hd__nor2_2 _1821_ (.A(net578),
    .B(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__or2_4 _1822_ (.A(net577),
    .B(_0559_),
    .X(_0561_));
 sky130_fd_sc_hd__nand2_1 _1823_ (.A(_0539_),
    .B(_0549_),
    .Y(_0562_));
 sky130_fd_sc_hd__nor2_2 _1824_ (.A(net577),
    .B(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__or2_2 _1825_ (.A(net577),
    .B(_0562_),
    .X(_0564_));
 sky130_fd_sc_hd__a21o_1 _1826_ (.A1(\vga.verticalFrontPorchCompare[0] ),
    .A2(net571),
    .B1(_0558_),
    .X(_0565_));
 sky130_fd_sc_hd__and3_1 _1827_ (.A(net602),
    .B(net579),
    .C(_0536_),
    .X(_0566_));
 sky130_fd_sc_hd__and4_1 _1828_ (.A(_1356_),
    .B(_1357_),
    .C(_0524_),
    .D(_0525_),
    .X(_0567_));
 sky130_fd_sc_hd__or3b_2 _1829_ (.A(\wbPeripheralBusInterface.currentAddress[4] ),
    .B(_0267_),
    .C_N(_0524_),
    .X(_0568_));
 sky130_fd_sc_hd__inv_2 _1830_ (.A(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__nor2_2 _1831_ (.A(_0545_),
    .B(_0568_),
    .Y(_0570_));
 sky130_fd_sc_hd__and3_1 _1832_ (.A(\wbPeripheralBusInterface.currentAddress[2] ),
    .B(net312),
    .C(_0525_),
    .X(_0571_));
 sky130_fd_sc_hd__a21o_1 _1833_ (.A1(\vga.horizontalSyncPulseCompare[0] ),
    .A2(net567),
    .B1(net517),
    .X(_0572_));
 sky130_fd_sc_hd__or4b_4 _1834_ (.A(_1355_),
    .B(_0267_),
    .C(net577),
    .D_N(_0526_),
    .X(_0573_));
 sky130_fd_sc_hd__a21o_1 _1835_ (.A1(\vga.stateRegister.baseReadData[0] ),
    .A2(net570),
    .B1(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__and3_1 _1836_ (.A(\vga.verticalSyncPulseCompare[0] ),
    .B(net570),
    .C(_0554_),
    .X(_0575_));
 sky130_fd_sc_hd__a31o_1 _1837_ (.A1(_0553_),
    .A2(_0555_),
    .A3(_0574_),
    .B1(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__or3b_4 _1838_ (.A(\wbPeripheralBusInterface.currentAddress[4] ),
    .B(_0267_),
    .C_N(_0526_),
    .X(_0577_));
 sky130_fd_sc_hd__nor2_2 _1839_ (.A(net577),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__or2_4 _1840_ (.A(net577),
    .B(_0577_),
    .X(_0579_));
 sky130_fd_sc_hd__a21o_1 _1841_ (.A1(\vga.verticalVisibleAreaCompare[0] ),
    .A2(net571),
    .B1(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__a31o_1 _1842_ (.A1(\vga.horizontalWholeLineCompare[0] ),
    .A2(net568),
    .A3(net515),
    .B1(net518),
    .X(_0581_));
 sky130_fd_sc_hd__a41o_2 _1843_ (.A1(net514),
    .A2(_0565_),
    .A3(_0576_),
    .A4(_0580_),
    .B1(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__and3_1 _1844_ (.A(net519),
    .B(_0572_),
    .C(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__and3_2 _1845_ (.A(net565),
    .B(net579),
    .C(_0542_),
    .X(_0584_));
 sky130_fd_sc_hd__a21o_1 _1846_ (.A1(\vga.horizontalFrontPorchCompare[0] ),
    .A2(_0584_),
    .B1(_0583_),
    .X(_0585_));
 sky130_fd_sc_hd__a31o_1 _1847_ (.A1(\vga.horizontalVisibleAreaCompare[0] ),
    .A2(net565),
    .A3(_0537_),
    .B1(_0528_),
    .X(_0586_));
 sky130_fd_sc_hd__a21o_1 _1848_ (.A1(_0538_),
    .A2(_0585_),
    .B1(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__o211a_2 _1849_ (.A1(net530),
    .A2(_0534_),
    .B1(_0587_),
    .C1(_0530_),
    .X(_0588_));
 sky130_fd_sc_hd__a21o_2 _1850_ (.A1(_1352_),
    .A2(net578),
    .B1(net527),
    .X(_0589_));
 sky130_fd_sc_hd__o22a_1 _1851_ (.A1(net522),
    .A2(_0588_),
    .B1(net513),
    .B2(net444),
    .X(_0590_));
 sky130_fd_sc_hd__or2_1 _1852_ (.A(net610),
    .B(_0590_),
    .X(_0000_));
 sky130_fd_sc_hd__a21o_1 _1853_ (.A1(\vga.configuration[1] ),
    .A2(net565),
    .B1(net521),
    .X(_0591_));
 sky130_fd_sc_hd__a221o_1 _1854_ (.A1(net27),
    .A2(net555),
    .B1(net548),
    .B2(net136),
    .C1(net561),
    .X(_0592_));
 sky130_fd_sc_hd__a21o_2 _1855_ (.A1(net151),
    .A2(net544),
    .B1(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__or2_1 _1856_ (.A(net12),
    .B(net557),
    .X(_0594_));
 sky130_fd_sc_hd__a31o_2 _1857_ (.A1(_0533_),
    .A2(_0593_),
    .A3(_0594_),
    .B1(net530),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _1858_ (.A0(\vga.stateRegister.baseReadData[1] ),
    .A1(\vga.verticalWholeLineCompare[1] ),
    .S(_0552_),
    .X(_0596_));
 sky130_fd_sc_hd__a41o_1 _1859_ (.A1(\wbPeripheralBusInterface.currentAddress[4] ),
    .A2(net314),
    .A3(_0275_),
    .A4(_0526_),
    .B1(_0552_),
    .X(_0597_));
 sky130_fd_sc_hd__a21o_1 _1860_ (.A1(\vga.verticalSyncPulseCompare[1] ),
    .A2(net569),
    .B1(_0555_),
    .X(_0598_));
 sky130_fd_sc_hd__a21o_1 _1861_ (.A1(\vga.horizontalSyncPulseCompare[1] ),
    .A2(net567),
    .B1(net517),
    .X(_0599_));
 sky130_fd_sc_hd__and3_1 _1862_ (.A(\vga.horizontalVisibleAreaCompare[1] ),
    .B(net567),
    .C(_0537_),
    .X(_0600_));
 sky130_fd_sc_hd__a21o_1 _1863_ (.A1(\vga.verticalVisibleAreaCompare[1] ),
    .A2(net568),
    .B1(_0579_),
    .X(_0601_));
 sky130_fd_sc_hd__o21a_2 _1864_ (.A1(net578),
    .A2(_0551_),
    .B1(_0573_),
    .X(_0602_));
 sky130_fd_sc_hd__a21o_1 _1865_ (.A1(net569),
    .A2(_0596_),
    .B1(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__a31o_1 _1866_ (.A1(\vga.verticalFrontPorchCompare[1] ),
    .A2(net569),
    .A3(_0557_),
    .B1(_0578_),
    .X(_0604_));
 sky130_fd_sc_hd__a31o_1 _1867_ (.A1(net516),
    .A2(_0598_),
    .A3(_0603_),
    .B1(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__a31o_1 _1868_ (.A1(\vga.horizontalWholeLineCompare[1] ),
    .A2(net568),
    .A3(net515),
    .B1(net518),
    .X(_0606_));
 sky130_fd_sc_hd__a31o_2 _1869_ (.A1(net514),
    .A2(_0601_),
    .A3(_0605_),
    .B1(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__a32o_1 _1870_ (.A1(net519),
    .A2(_0599_),
    .A3(_0607_),
    .B1(_0584_),
    .B2(\vga.horizontalFrontPorchCompare[1] ),
    .X(_0608_));
 sky130_fd_sc_hd__a21o_1 _1871_ (.A1(net520),
    .A2(_0608_),
    .B1(_0600_),
    .X(_0609_));
 sky130_fd_sc_hd__and3_2 _1872_ (.A(_0591_),
    .B(_0595_),
    .C(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__o22a_1 _1873_ (.A1(net455),
    .A2(net513),
    .B1(_0610_),
    .B2(net522),
    .X(_0611_));
 sky130_fd_sc_hd__or2_1 _1874_ (.A(net610),
    .B(_0611_),
    .X(_0001_));
 sky130_fd_sc_hd__a21o_1 _1875_ (.A1(\vga.configuration[2] ),
    .A2(net565),
    .B1(_0529_),
    .X(_0612_));
 sky130_fd_sc_hd__a221o_1 _1876_ (.A1(net28),
    .A2(net555),
    .B1(net548),
    .B2(net147),
    .C1(net561),
    .X(_0613_));
 sky130_fd_sc_hd__a21o_4 _1877_ (.A1(net152),
    .A2(net544),
    .B1(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__or2_1 _1878_ (.A(net23),
    .B(net557),
    .X(_0615_));
 sky130_fd_sc_hd__a31o_2 _1879_ (.A1(_0533_),
    .A2(_0614_),
    .A3(_0615_),
    .B1(net530),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _1880_ (.A0(\vga.stateRegister.baseReadData[2] ),
    .A1(\vga.verticalWholeLineCompare[2] ),
    .S(_0552_),
    .X(_0617_));
 sky130_fd_sc_hd__a21o_1 _1881_ (.A1(\vga.verticalSyncPulseCompare[2] ),
    .A2(net569),
    .B1(_0555_),
    .X(_0618_));
 sky130_fd_sc_hd__a21o_1 _1882_ (.A1(\vga.horizontalSyncPulseCompare[2] ),
    .A2(net567),
    .B1(net517),
    .X(_0619_));
 sky130_fd_sc_hd__and3_1 _1883_ (.A(\vga.horizontalVisibleAreaCompare[2] ),
    .B(net567),
    .C(_0537_),
    .X(_0620_));
 sky130_fd_sc_hd__a21o_1 _1884_ (.A1(\vga.verticalVisibleAreaCompare[2] ),
    .A2(net568),
    .B1(_0579_),
    .X(_0621_));
 sky130_fd_sc_hd__a21o_1 _1885_ (.A1(net570),
    .A2(_0617_),
    .B1(_0602_),
    .X(_0622_));
 sky130_fd_sc_hd__a31o_1 _1886_ (.A1(\vga.verticalFrontPorchCompare[2] ),
    .A2(net569),
    .A3(_0557_),
    .B1(_0578_),
    .X(_0623_));
 sky130_fd_sc_hd__a31o_1 _1887_ (.A1(net516),
    .A2(_0618_),
    .A3(_0622_),
    .B1(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__a31o_1 _1888_ (.A1(\vga.horizontalWholeLineCompare[2] ),
    .A2(net568),
    .A3(net515),
    .B1(net518),
    .X(_0625_));
 sky130_fd_sc_hd__a31o_2 _1889_ (.A1(net514),
    .A2(_0621_),
    .A3(_0624_),
    .B1(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__a32o_1 _1890_ (.A1(net519),
    .A2(_0619_),
    .A3(_0626_),
    .B1(_0584_),
    .B2(\vga.horizontalFrontPorchCompare[2] ),
    .X(_0627_));
 sky130_fd_sc_hd__a21o_1 _1891_ (.A1(net520),
    .A2(_0627_),
    .B1(_0620_),
    .X(_0628_));
 sky130_fd_sc_hd__and3_2 _1892_ (.A(_0612_),
    .B(_0616_),
    .C(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__o22a_1 _1893_ (.A1(net466),
    .A2(net513),
    .B1(_0629_),
    .B2(net522),
    .X(_0630_));
 sky130_fd_sc_hd__or2_1 _1894_ (.A(net610),
    .B(_0630_),
    .X(_0002_));
 sky130_fd_sc_hd__a21o_1 _1895_ (.A1(\vga.configuration[3] ),
    .A2(net565),
    .B1(net521),
    .X(_0631_));
 sky130_fd_sc_hd__a221o_1 _1896_ (.A1(net29),
    .A2(net555),
    .B1(net552),
    .B2(net158),
    .C1(net561),
    .X(_0632_));
 sky130_fd_sc_hd__a21o_4 _1897_ (.A1(net153),
    .A2(net544),
    .B1(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__or2_1 _1898_ (.A(net34),
    .B(net557),
    .X(_0634_));
 sky130_fd_sc_hd__a31o_2 _1899_ (.A1(_0533_),
    .A2(_0633_),
    .A3(_0634_),
    .B1(net530),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _1900_ (.A0(\vga.stateRegister.baseReadData[3] ),
    .A1(\vga.verticalWholeLineCompare[3] ),
    .S(_0552_),
    .X(_0636_));
 sky130_fd_sc_hd__a21o_1 _1901_ (.A1(\vga.verticalSyncPulseCompare[3] ),
    .A2(net570),
    .B1(_0555_),
    .X(_0637_));
 sky130_fd_sc_hd__a21o_1 _1902_ (.A1(\vga.horizontalSyncPulseCompare[3] ),
    .A2(net567),
    .B1(net517),
    .X(_0638_));
 sky130_fd_sc_hd__and3_1 _1903_ (.A(\vga.horizontalVisibleAreaCompare[3] ),
    .B(net567),
    .C(_0537_),
    .X(_0639_));
 sky130_fd_sc_hd__a21o_1 _1904_ (.A1(\vga.verticalVisibleAreaCompare[3] ),
    .A2(net568),
    .B1(_0579_),
    .X(_0640_));
 sky130_fd_sc_hd__a21o_1 _1905_ (.A1(net570),
    .A2(_0636_),
    .B1(_0602_),
    .X(_0641_));
 sky130_fd_sc_hd__a31o_1 _1906_ (.A1(\vga.verticalFrontPorchCompare[3] ),
    .A2(net569),
    .A3(_0557_),
    .B1(_0578_),
    .X(_0642_));
 sky130_fd_sc_hd__a31o_1 _1907_ (.A1(net516),
    .A2(_0637_),
    .A3(_0641_),
    .B1(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__a31o_1 _1908_ (.A1(\vga.horizontalWholeLineCompare[3] ),
    .A2(net568),
    .A3(net515),
    .B1(net518),
    .X(_0644_));
 sky130_fd_sc_hd__a31o_2 _1909_ (.A1(net514),
    .A2(_0640_),
    .A3(_0643_),
    .B1(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__a32o_1 _1910_ (.A1(net519),
    .A2(_0638_),
    .A3(_0645_),
    .B1(_0584_),
    .B2(\vga.horizontalFrontPorchCompare[3] ),
    .X(_0646_));
 sky130_fd_sc_hd__a21o_1 _1911_ (.A1(net520),
    .A2(_0646_),
    .B1(_0639_),
    .X(_0647_));
 sky130_fd_sc_hd__and3_2 _1912_ (.A(_0631_),
    .B(_0635_),
    .C(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__o22a_1 _1913_ (.A1(net469),
    .A2(net513),
    .B1(_0648_),
    .B2(net522),
    .X(_0649_));
 sky130_fd_sc_hd__or2_1 _1914_ (.A(net611),
    .B(_0649_),
    .X(_0003_));
 sky130_fd_sc_hd__a21o_1 _1915_ (.A1(\vga.configuration[4] ),
    .A2(net565),
    .B1(_0529_),
    .X(_0650_));
 sky130_fd_sc_hd__a221o_1 _1916_ (.A1(net30),
    .A2(net555),
    .B1(net552),
    .B2(net169),
    .C1(net561),
    .X(_0651_));
 sky130_fd_sc_hd__a21o_2 _1917_ (.A1(net154),
    .A2(net544),
    .B1(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__or2_2 _1918_ (.A(net45),
    .B(net557),
    .X(_0653_));
 sky130_fd_sc_hd__a31o_2 _1919_ (.A1(_0533_),
    .A2(_0652_),
    .A3(_0653_),
    .B1(net530),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _1920_ (.A0(\vga.stateRegister.baseReadData[4] ),
    .A1(\vga.verticalWholeLineCompare[4] ),
    .S(_0552_),
    .X(_0655_));
 sky130_fd_sc_hd__a21o_1 _1921_ (.A1(\vga.verticalSyncPulseCompare[4] ),
    .A2(net570),
    .B1(_0555_),
    .X(_0656_));
 sky130_fd_sc_hd__a21o_1 _1922_ (.A1(\vga.horizontalSyncPulseCompare[4] ),
    .A2(net565),
    .B1(net517),
    .X(_0657_));
 sky130_fd_sc_hd__a31o_1 _1923_ (.A1(\vga.horizontalVisibleAreaCompare[4] ),
    .A2(net565),
    .A3(_0537_),
    .B1(_0528_),
    .X(_0658_));
 sky130_fd_sc_hd__a21o_1 _1924_ (.A1(\vga.verticalVisibleAreaCompare[4] ),
    .A2(net571),
    .B1(_0579_),
    .X(_0659_));
 sky130_fd_sc_hd__a21o_1 _1925_ (.A1(net570),
    .A2(_0655_),
    .B1(_0602_),
    .X(_0660_));
 sky130_fd_sc_hd__a31o_1 _1926_ (.A1(\vga.verticalFrontPorchCompare[4] ),
    .A2(net569),
    .A3(_0557_),
    .B1(_0578_),
    .X(_0661_));
 sky130_fd_sc_hd__a31o_1 _1927_ (.A1(net516),
    .A2(_0656_),
    .A3(_0660_),
    .B1(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__a31o_1 _1928_ (.A1(\vga.horizontalWholeLineCompare[4] ),
    .A2(net568),
    .A3(_0563_),
    .B1(_0547_),
    .X(_0663_));
 sky130_fd_sc_hd__a31o_2 _1929_ (.A1(net514),
    .A2(_0659_),
    .A3(_0662_),
    .B1(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__a32o_1 _1930_ (.A1(_0544_),
    .A2(_0657_),
    .A3(_0664_),
    .B1(_0584_),
    .B2(\vga.horizontalFrontPorchCompare[4] ),
    .X(_0665_));
 sky130_fd_sc_hd__a21o_1 _1931_ (.A1(_0538_),
    .A2(_0665_),
    .B1(_0658_),
    .X(_0666_));
 sky130_fd_sc_hd__and3_2 _1932_ (.A(_0650_),
    .B(_0654_),
    .C(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__o22a_1 _1933_ (.A1(net470),
    .A2(net513),
    .B1(_0667_),
    .B2(net522),
    .X(_0668_));
 sky130_fd_sc_hd__or2_1 _1934_ (.A(net612),
    .B(_0668_),
    .X(_0004_));
 sky130_fd_sc_hd__a21o_1 _1935_ (.A1(\vga.configuration[5] ),
    .A2(net566),
    .B1(net521),
    .X(_0669_));
 sky130_fd_sc_hd__a221o_1 _1936_ (.A1(net31),
    .A2(net555),
    .B1(net548),
    .B2(net180),
    .C1(net561),
    .X(_0670_));
 sky130_fd_sc_hd__a21o_2 _1937_ (.A1(net155),
    .A2(net544),
    .B1(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__or2_2 _1938_ (.A(net56),
    .B(net557),
    .X(_0672_));
 sky130_fd_sc_hd__a31o_2 _1939_ (.A1(_0533_),
    .A2(_0671_),
    .A3(_0672_),
    .B1(net530),
    .X(_0673_));
 sky130_fd_sc_hd__a31o_1 _1940_ (.A1(\vga.horizontalSyncPulseCompare[5] ),
    .A2(net601),
    .A3(net518),
    .B1(_0543_),
    .X(_0674_));
 sky130_fd_sc_hd__a22o_1 _1941_ (.A1(\vga.verticalWholeLineCompare[5] ),
    .A2(_0552_),
    .B1(_0554_),
    .B2(\vga.verticalSyncPulseCompare[5] ),
    .X(_0675_));
 sky130_fd_sc_hd__nor2_4 _1942_ (.A(_0554_),
    .B(_0597_),
    .Y(_0676_));
 sky130_fd_sc_hd__a21o_1 _1943_ (.A1(net569),
    .A2(_0675_),
    .B1(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__a21o_1 _1944_ (.A1(\vga.verticalFrontPorchCompare[5] ),
    .A2(net571),
    .B1(net516),
    .X(_0678_));
 sky130_fd_sc_hd__a31o_1 _1945_ (.A1(\vga.verticalVisibleAreaCompare[5] ),
    .A2(net599),
    .A3(_0560_),
    .B1(net515),
    .X(_0679_));
 sky130_fd_sc_hd__a31o_2 _1946_ (.A1(_0561_),
    .A2(_0677_),
    .A3(_0678_),
    .B1(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__a21o_1 _1947_ (.A1(\vga.horizontalWholeLineCompare[5] ),
    .A2(net572),
    .B1(_0564_),
    .X(_0681_));
 sky130_fd_sc_hd__a31o_1 _1948_ (.A1(net517),
    .A2(_0680_),
    .A3(_0681_),
    .B1(_0674_),
    .X(_0682_));
 sky130_fd_sc_hd__a21o_1 _1949_ (.A1(\vga.horizontalFrontPorchCompare[5] ),
    .A2(net565),
    .B1(net519),
    .X(_0683_));
 sky130_fd_sc_hd__a32o_1 _1950_ (.A1(net520),
    .A2(_0682_),
    .A3(_0683_),
    .B1(_0566_),
    .B2(\vga.horizontalVisibleAreaCompare[5] ),
    .X(_0684_));
 sky130_fd_sc_hd__and3_2 _1951_ (.A(_0669_),
    .B(_0673_),
    .C(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__o22a_1 _1952_ (.A1(net471),
    .A2(_0589_),
    .B1(_0685_),
    .B2(net522),
    .X(_0686_));
 sky130_fd_sc_hd__or2_1 _1953_ (.A(net612),
    .B(_0686_),
    .X(_0005_));
 sky130_fd_sc_hd__a221o_1 _1954_ (.A1(net32),
    .A2(net555),
    .B1(net552),
    .B2(net185),
    .C1(net561),
    .X(_0687_));
 sky130_fd_sc_hd__a21o_2 _1955_ (.A1(net156),
    .A2(_0282_),
    .B1(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__or2_2 _1956_ (.A(net61),
    .B(net557),
    .X(_0689_));
 sky130_fd_sc_hd__a31o_2 _1957_ (.A1(_0533_),
    .A2(_0688_),
    .A3(_0689_),
    .B1(net531),
    .X(_0690_));
 sky130_fd_sc_hd__a21o_1 _1958_ (.A1(\vga.configuration[6] ),
    .A2(net566),
    .B1(net521),
    .X(_0691_));
 sky130_fd_sc_hd__a31o_1 _1959_ (.A1(\vga.horizontalSyncPulseCompare[6] ),
    .A2(net601),
    .A3(net518),
    .B1(_0543_),
    .X(_0692_));
 sky130_fd_sc_hd__a22o_1 _1960_ (.A1(\vga.verticalWholeLineCompare[6] ),
    .A2(_0552_),
    .B1(_0554_),
    .B2(\vga.verticalSyncPulseCompare[6] ),
    .X(_0693_));
 sky130_fd_sc_hd__a21o_1 _1961_ (.A1(net569),
    .A2(_0693_),
    .B1(_0676_),
    .X(_0694_));
 sky130_fd_sc_hd__a21o_1 _1962_ (.A1(\vga.verticalFrontPorchCompare[6] ),
    .A2(net571),
    .B1(net516),
    .X(_0695_));
 sky130_fd_sc_hd__a31o_1 _1963_ (.A1(\vga.verticalVisibleAreaCompare[6] ),
    .A2(net600),
    .A3(_0560_),
    .B1(net515),
    .X(_0696_));
 sky130_fd_sc_hd__a31o_2 _1964_ (.A1(_0561_),
    .A2(_0694_),
    .A3(_0695_),
    .B1(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__a21o_1 _1965_ (.A1(\vga.horizontalWholeLineCompare[6] ),
    .A2(net568),
    .B1(net514),
    .X(_0698_));
 sky130_fd_sc_hd__a31o_1 _1966_ (.A1(net517),
    .A2(_0697_),
    .A3(_0698_),
    .B1(_0692_),
    .X(_0699_));
 sky130_fd_sc_hd__a21o_1 _1967_ (.A1(\vga.horizontalFrontPorchCompare[6] ),
    .A2(net567),
    .B1(net519),
    .X(_0700_));
 sky130_fd_sc_hd__a32o_1 _1968_ (.A1(net520),
    .A2(_0699_),
    .A3(_0700_),
    .B1(_0566_),
    .B2(\vga.horizontalVisibleAreaCompare[6] ),
    .X(_0701_));
 sky130_fd_sc_hd__and3_2 _1969_ (.A(_0690_),
    .B(_0691_),
    .C(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__o22a_1 _1970_ (.A1(net472),
    .A2(net513),
    .B1(_0702_),
    .B2(net523),
    .X(_0703_));
 sky130_fd_sc_hd__or2_1 _1971_ (.A(net612),
    .B(_0703_),
    .X(_0006_));
 sky130_fd_sc_hd__a221o_1 _1972_ (.A1(net33),
    .A2(net556),
    .B1(net548),
    .B2(net186),
    .C1(net564),
    .X(_0704_));
 sky130_fd_sc_hd__a21o_2 _1973_ (.A1(net157),
    .A2(net544),
    .B1(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__or2_2 _1974_ (.A(net62),
    .B(net557),
    .X(_0706_));
 sky130_fd_sc_hd__a31o_2 _1975_ (.A1(_0533_),
    .A2(_0705_),
    .A3(_0706_),
    .B1(net531),
    .X(_0707_));
 sky130_fd_sc_hd__a21o_1 _1976_ (.A1(\vga.configuration[7] ),
    .A2(net566),
    .B1(net521),
    .X(_0708_));
 sky130_fd_sc_hd__a31o_1 _1977_ (.A1(\vga.horizontalSyncPulseCompare[7] ),
    .A2(net601),
    .A3(net518),
    .B1(_0543_),
    .X(_0709_));
 sky130_fd_sc_hd__a22o_1 _1978_ (.A1(\vga.verticalWholeLineCompare[7] ),
    .A2(_0552_),
    .B1(_0554_),
    .B2(\vga.verticalSyncPulseCompare[7] ),
    .X(_0710_));
 sky130_fd_sc_hd__a21o_1 _1979_ (.A1(net569),
    .A2(_0710_),
    .B1(_0676_),
    .X(_0711_));
 sky130_fd_sc_hd__a21o_1 _1980_ (.A1(\vga.verticalFrontPorchCompare[7] ),
    .A2(net571),
    .B1(net516),
    .X(_0712_));
 sky130_fd_sc_hd__a31o_1 _1981_ (.A1(\vga.verticalVisibleAreaCompare[7] ),
    .A2(net600),
    .A3(_0560_),
    .B1(net515),
    .X(_0713_));
 sky130_fd_sc_hd__a31o_2 _1982_ (.A1(_0561_),
    .A2(_0711_),
    .A3(_0712_),
    .B1(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__a21o_1 _1983_ (.A1(\vga.horizontalWholeLineCompare[7] ),
    .A2(net568),
    .B1(net514),
    .X(_0715_));
 sky130_fd_sc_hd__a31o_1 _1984_ (.A1(_0548_),
    .A2(_0714_),
    .A3(_0715_),
    .B1(_0709_),
    .X(_0716_));
 sky130_fd_sc_hd__a21o_1 _1985_ (.A1(\vga.horizontalFrontPorchCompare[7] ),
    .A2(net567),
    .B1(net519),
    .X(_0717_));
 sky130_fd_sc_hd__a32o_1 _1986_ (.A1(net520),
    .A2(_0716_),
    .A3(_0717_),
    .B1(_0566_),
    .B2(\vga.horizontalVisibleAreaCompare[7] ),
    .X(_0718_));
 sky130_fd_sc_hd__and3_2 _1987_ (.A(_0707_),
    .B(_0708_),
    .C(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__o22a_1 _1988_ (.A1(net473),
    .A2(net513),
    .B1(_0719_),
    .B2(net522),
    .X(_0720_));
 sky130_fd_sc_hd__or2_1 _1989_ (.A(net612),
    .B(_0720_),
    .X(_0007_));
 sky130_fd_sc_hd__or2_1 _1990_ (.A(net474),
    .B(net513),
    .X(_0721_));
 sky130_fd_sc_hd__and3_1 _1991_ (.A(net597),
    .B(net579),
    .C(_0536_),
    .X(_0722_));
 sky130_fd_sc_hd__a31o_1 _1992_ (.A1(\vga.horizontalSyncPulseCompare[8] ),
    .A2(net596),
    .A3(net518),
    .B1(_0543_),
    .X(_0723_));
 sky130_fd_sc_hd__a22o_1 _1993_ (.A1(\vga.verticalWholeLineCompare[8] ),
    .A2(_0552_),
    .B1(_0554_),
    .B2(\vga.verticalSyncPulseCompare[8] ),
    .X(_0724_));
 sky130_fd_sc_hd__a21o_1 _1994_ (.A1(net573),
    .A2(_0724_),
    .B1(_0676_),
    .X(_0725_));
 sky130_fd_sc_hd__a21o_1 _1995_ (.A1(\vga.verticalFrontPorchCompare[8] ),
    .A2(net573),
    .B1(net516),
    .X(_0726_));
 sky130_fd_sc_hd__a31o_1 _1996_ (.A1(\vga.verticalVisibleAreaCompare[8] ),
    .A2(net596),
    .A3(_0560_),
    .B1(net515),
    .X(_0727_));
 sky130_fd_sc_hd__a31o_1 _1997_ (.A1(_0561_),
    .A2(_0725_),
    .A3(_0726_),
    .B1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__a21o_1 _1998_ (.A1(\vga.horizontalWholeLineCompare[8] ),
    .A2(net574),
    .B1(net514),
    .X(_0729_));
 sky130_fd_sc_hd__a31o_1 _1999_ (.A1(_0548_),
    .A2(_0728_),
    .A3(_0729_),
    .B1(_0723_),
    .X(_0730_));
 sky130_fd_sc_hd__a21o_1 _2000_ (.A1(\vga.horizontalFrontPorchCompare[8] ),
    .A2(net573),
    .B1(net519),
    .X(_0731_));
 sky130_fd_sc_hd__a32o_1 _2001_ (.A1(net520),
    .A2(_0730_),
    .A3(_0731_),
    .B1(_0722_),
    .B2(\vga.horizontalVisibleAreaCompare[8] ),
    .X(_0732_));
 sky130_fd_sc_hd__a21o_1 _2002_ (.A1(\vga.configuration[8] ),
    .A2(net573),
    .B1(net521),
    .X(_0733_));
 sky130_fd_sc_hd__a221o_1 _2003_ (.A1(net35),
    .A2(net556),
    .B1(net547),
    .B2(net159),
    .C1(net562),
    .X(_0734_));
 sky130_fd_sc_hd__a21o_2 _2004_ (.A1(net187),
    .A2(net548),
    .B1(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__and3_4 _2005_ (.A(\videoMemory.wbReadReady ),
    .B(net596),
    .C(net580),
    .X(_0736_));
 sky130_fd_sc_hd__or2_2 _2006_ (.A(net63),
    .B(net557),
    .X(_0737_));
 sky130_fd_sc_hd__a31o_2 _2007_ (.A1(_0735_),
    .A2(_0736_),
    .A3(_0737_),
    .B1(net530),
    .X(_0738_));
 sky130_fd_sc_hd__a31o_1 _2008_ (.A1(_0732_),
    .A2(_0733_),
    .A3(_0738_),
    .B1(net525),
    .X(_0739_));
 sky130_fd_sc_hd__a21o_1 _2009_ (.A1(_0721_),
    .A2(_0739_),
    .B1(net612),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _2010_ (.A(net475),
    .B(net513),
    .X(_0740_));
 sky130_fd_sc_hd__a21o_1 _2011_ (.A1(\vga.configuration[9] ),
    .A2(net573),
    .B1(net521),
    .X(_0741_));
 sky130_fd_sc_hd__a221o_4 _2012_ (.A1(net188),
    .A2(net549),
    .B1(net545),
    .B2(net160),
    .C1(net562),
    .X(_0742_));
 sky130_fd_sc_hd__a21o_1 _2013_ (.A1(net36),
    .A2(net553),
    .B1(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__or2_1 _2014_ (.A(net64),
    .B(net557),
    .X(_0744_));
 sky130_fd_sc_hd__a31o_2 _2015_ (.A1(_0736_),
    .A2(_0743_),
    .A3(_0744_),
    .B1(net530),
    .X(_0745_));
 sky130_fd_sc_hd__a31o_1 _2016_ (.A1(\vga.horizontalSyncPulseCompare[9] ),
    .A2(net596),
    .A3(net518),
    .B1(_0543_),
    .X(_0746_));
 sky130_fd_sc_hd__a22o_1 _2017_ (.A1(\vga.verticalWholeLineCompare[9] ),
    .A2(_0552_),
    .B1(_0554_),
    .B2(\vga.verticalSyncPulseCompare[9] ),
    .X(_0747_));
 sky130_fd_sc_hd__a21o_1 _2018_ (.A1(net574),
    .A2(_0747_),
    .B1(_0676_),
    .X(_0748_));
 sky130_fd_sc_hd__a21o_1 _2019_ (.A1(\vga.verticalFrontPorchCompare[9] ),
    .A2(net574),
    .B1(net516),
    .X(_0749_));
 sky130_fd_sc_hd__a31o_1 _2020_ (.A1(\vga.verticalVisibleAreaCompare[9] ),
    .A2(net596),
    .A3(_0560_),
    .B1(net515),
    .X(_0750_));
 sky130_fd_sc_hd__a31o_1 _2021_ (.A1(_0561_),
    .A2(_0748_),
    .A3(_0749_),
    .B1(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__a21o_1 _2022_ (.A1(\vga.horizontalWholeLineCompare[9] ),
    .A2(net574),
    .B1(net514),
    .X(_0752_));
 sky130_fd_sc_hd__a31o_1 _2023_ (.A1(net517),
    .A2(_0751_),
    .A3(_0752_),
    .B1(_0746_),
    .X(_0753_));
 sky130_fd_sc_hd__a21o_1 _2024_ (.A1(\vga.horizontalFrontPorchCompare[9] ),
    .A2(net573),
    .B1(net519),
    .X(_0754_));
 sky130_fd_sc_hd__a32o_1 _2025_ (.A1(net520),
    .A2(_0753_),
    .A3(_0754_),
    .B1(_0722_),
    .B2(\vga.horizontalVisibleAreaCompare[9] ),
    .X(_0755_));
 sky130_fd_sc_hd__a31o_2 _2026_ (.A1(_0741_),
    .A2(_0745_),
    .A3(_0755_),
    .B1(net525),
    .X(_0756_));
 sky130_fd_sc_hd__a21o_1 _2027_ (.A1(_0740_),
    .A2(_0756_),
    .B1(net612),
    .X(_0009_));
 sky130_fd_sc_hd__a221o_1 _2028_ (.A1(net37),
    .A2(net555),
    .B1(net548),
    .B2(net126),
    .C1(net561),
    .X(_0757_));
 sky130_fd_sc_hd__a21o_4 _2029_ (.A1(net161),
    .A2(net544),
    .B1(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__o211a_2 _2030_ (.A1(net2),
    .A2(net559),
    .B1(_0736_),
    .C1(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__and3_1 _2031_ (.A(net516),
    .B(_0561_),
    .C(net514),
    .X(_0760_));
 sky130_fd_sc_hd__a31o_1 _2032_ (.A1(\vga.horizontalWholeLineCompare[10] ),
    .A2(net574),
    .A3(net515),
    .B1(net518),
    .X(_0761_));
 sky130_fd_sc_hd__a21o_1 _2033_ (.A1(_0676_),
    .A2(_0760_),
    .B1(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__a21o_1 _2034_ (.A1(\vga.horizontalSyncPulseCompare[10] ),
    .A2(net573),
    .B1(net517),
    .X(_0763_));
 sky130_fd_sc_hd__a21o_1 _2035_ (.A1(\vga.horizontalFrontPorchCompare[10] ),
    .A2(net573),
    .B1(net519),
    .X(_0764_));
 sky130_fd_sc_hd__and3_1 _2036_ (.A(net520),
    .B(_0763_),
    .C(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__a22o_1 _2037_ (.A1(\vga.horizontalVisibleAreaCompare[10] ),
    .A2(_0722_),
    .B1(_0762_),
    .B2(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__and4_1 _2038_ (.A(net521),
    .B(net520),
    .C(_0544_),
    .D(net517),
    .X(_0767_));
 sky130_fd_sc_hd__and3_4 _2039_ (.A(_0676_),
    .B(_0760_),
    .C(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__a31o_1 _2040_ (.A1(\vga.configuration[10] ),
    .A2(net597),
    .A3(_0528_),
    .B1(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__a21o_1 _2041_ (.A1(net521),
    .A2(_0766_),
    .B1(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__o21a_2 _2042_ (.A1(net531),
    .A2(_0759_),
    .B1(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__o22a_1 _2043_ (.A1(net445),
    .A2(net513),
    .B1(_0771_),
    .B2(net523),
    .X(_0772_));
 sky130_fd_sc_hd__or2_1 _2044_ (.A(net612),
    .B(_0772_),
    .X(_0010_));
 sky130_fd_sc_hd__a221o_4 _2045_ (.A1(net127),
    .A2(net549),
    .B1(net546),
    .B2(net162),
    .C1(net562),
    .X(_0773_));
 sky130_fd_sc_hd__a21o_1 _2046_ (.A1(net38),
    .A2(net553),
    .B1(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__o211a_4 _2047_ (.A1(net3),
    .A2(net557),
    .B1(_0736_),
    .C1(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__and3_1 _2048_ (.A(\vga.configuration[11] ),
    .B(net598),
    .C(_0528_),
    .X(_0776_));
 sky130_fd_sc_hd__o22a_1 _2049_ (.A1(net531),
    .A2(_0775_),
    .B1(_0776_),
    .B2(_0768_),
    .X(_0777_));
 sky130_fd_sc_hd__o22a_1 _2050_ (.A1(net446),
    .A2(_0589_),
    .B1(_0777_),
    .B2(net523),
    .X(_0778_));
 sky130_fd_sc_hd__or2_1 _2051_ (.A(net612),
    .B(_0778_),
    .X(_0011_));
 sky130_fd_sc_hd__a221o_4 _2052_ (.A1(net128),
    .A2(net550),
    .B1(net546),
    .B2(net163),
    .C1(net563),
    .X(_0779_));
 sky130_fd_sc_hd__a21o_1 _2053_ (.A1(net39),
    .A2(net553),
    .B1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__o211a_4 _2054_ (.A1(net4),
    .A2(net558),
    .B1(_0736_),
    .C1(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__and3_1 _2055_ (.A(\vga.configuration[12] ),
    .B(net598),
    .C(_0528_),
    .X(_0782_));
 sky130_fd_sc_hd__o22a_1 _2056_ (.A1(net531),
    .A2(_0781_),
    .B1(_0782_),
    .B2(_0768_),
    .X(_0783_));
 sky130_fd_sc_hd__o22a_1 _2057_ (.A1(net447),
    .A2(_0589_),
    .B1(_0783_),
    .B2(net522),
    .X(_0784_));
 sky130_fd_sc_hd__or2_1 _2058_ (.A(net612),
    .B(_0784_),
    .X(_0012_));
 sky130_fd_sc_hd__and2_1 _2059_ (.A(net531),
    .B(_0768_),
    .X(_0785_));
 sky130_fd_sc_hd__a221o_4 _2060_ (.A1(net129),
    .A2(net550),
    .B1(net546),
    .B2(net164),
    .C1(net563),
    .X(_0786_));
 sky130_fd_sc_hd__a21o_1 _2061_ (.A1(net40),
    .A2(net553),
    .B1(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__and2_2 _2062_ (.A(_0278_),
    .B(_0736_),
    .X(_0788_));
 sky130_fd_sc_hd__o211a_4 _2063_ (.A1(net5),
    .A2(net559),
    .B1(_0787_),
    .C1(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__o21a_2 _2064_ (.A1(net510),
    .A2(_0789_),
    .B1(net527),
    .X(_0790_));
 sky130_fd_sc_hd__a21o_2 _2065_ (.A1(_1352_),
    .A2(net578),
    .B1(net611),
    .X(_0791_));
 sky130_fd_sc_hd__a211o_1 _2066_ (.A1(net448),
    .A2(net524),
    .B1(_0790_),
    .C1(net536),
    .X(_0013_));
 sky130_fd_sc_hd__a221o_1 _2067_ (.A1(net41),
    .A2(net555),
    .B1(net548),
    .B2(net130),
    .C1(net561),
    .X(_0792_));
 sky130_fd_sc_hd__a21o_4 _2068_ (.A1(net165),
    .A2(net544),
    .B1(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__o211a_4 _2069_ (.A1(net6),
    .A2(net559),
    .B1(_0788_),
    .C1(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__o21a_1 _2070_ (.A1(net510),
    .A2(_0794_),
    .B1(net527),
    .X(_0795_));
 sky130_fd_sc_hd__a211o_1 _2071_ (.A1(net449),
    .A2(net523),
    .B1(net536),
    .C1(_0795_),
    .X(_0014_));
 sky130_fd_sc_hd__a221o_4 _2072_ (.A1(net131),
    .A2(net550),
    .B1(net546),
    .B2(net166),
    .C1(net562),
    .X(_0796_));
 sky130_fd_sc_hd__a21o_1 _2073_ (.A1(net42),
    .A2(net554),
    .B1(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__o211a_2 _2074_ (.A1(net7),
    .A2(net559),
    .B1(_0788_),
    .C1(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__o21a_4 _2075_ (.A1(net509),
    .A2(_0798_),
    .B1(net526),
    .X(_0799_));
 sky130_fd_sc_hd__a211o_1 _2076_ (.A1(net450),
    .A2(net524),
    .B1(net537),
    .C1(_0799_),
    .X(_0015_));
 sky130_fd_sc_hd__and3_4 _2077_ (.A(\videoMemory.wbReadReady ),
    .B(net370),
    .C(_0278_),
    .X(_0800_));
 sky130_fd_sc_hd__a221o_1 _2078_ (.A1(net43),
    .A2(net555),
    .B1(net548),
    .B2(net132),
    .C1(net561),
    .X(_0801_));
 sky130_fd_sc_hd__a21o_2 _2079_ (.A1(net167),
    .A2(net544),
    .B1(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__o211a_1 _2080_ (.A1(net8),
    .A2(net560),
    .B1(_0800_),
    .C1(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__o21a_4 _2081_ (.A1(net509),
    .A2(_0803_),
    .B1(net526),
    .X(_0804_));
 sky130_fd_sc_hd__a211o_1 _2082_ (.A1(net451),
    .A2(net524),
    .B1(net537),
    .C1(_0804_),
    .X(_0016_));
 sky130_fd_sc_hd__a221o_1 _2083_ (.A1(net44),
    .A2(net556),
    .B1(net551),
    .B2(net133),
    .C1(net562),
    .X(_0805_));
 sky130_fd_sc_hd__a21o_2 _2084_ (.A1(net168),
    .A2(net547),
    .B1(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__o211a_1 _2085_ (.A1(net9),
    .A2(net560),
    .B1(_0800_),
    .C1(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__o21a_4 _2086_ (.A1(net509),
    .A2(_0807_),
    .B1(net526),
    .X(_0808_));
 sky130_fd_sc_hd__a211o_1 _2087_ (.A1(net452),
    .A2(net524),
    .B1(net537),
    .C1(_0808_),
    .X(_0017_));
 sky130_fd_sc_hd__a221o_1 _2088_ (.A1(net46),
    .A2(net556),
    .B1(net551),
    .B2(net134),
    .C1(net562),
    .X(_0809_));
 sky130_fd_sc_hd__a21o_2 _2089_ (.A1(net170),
    .A2(net547),
    .B1(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__o211a_1 _2090_ (.A1(net10),
    .A2(net560),
    .B1(_0800_),
    .C1(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__o21a_4 _2091_ (.A1(net510),
    .A2(_0811_),
    .B1(net527),
    .X(_0812_));
 sky130_fd_sc_hd__a211o_1 _2092_ (.A1(net453),
    .A2(net524),
    .B1(net536),
    .C1(_0812_),
    .X(_0018_));
 sky130_fd_sc_hd__a221o_1 _2093_ (.A1(net47),
    .A2(net555),
    .B1(net548),
    .B2(net135),
    .C1(net561),
    .X(_0813_));
 sky130_fd_sc_hd__a21o_2 _2094_ (.A1(net171),
    .A2(net544),
    .B1(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__o211a_1 _2095_ (.A1(net11),
    .A2(net560),
    .B1(_0800_),
    .C1(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__o21a_1 _2096_ (.A1(net509),
    .A2(_0815_),
    .B1(net526),
    .X(_0816_));
 sky130_fd_sc_hd__a211o_1 _2097_ (.A1(net454),
    .A2(net525),
    .B1(net538),
    .C1(_0816_),
    .X(_0019_));
 sky130_fd_sc_hd__a221o_1 _2098_ (.A1(net48),
    .A2(net556),
    .B1(net550),
    .B2(net137),
    .C1(net562),
    .X(_0817_));
 sky130_fd_sc_hd__a21o_2 _2099_ (.A1(net172),
    .A2(net546),
    .B1(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__o211a_1 _2100_ (.A1(net13),
    .A2(net560),
    .B1(_0800_),
    .C1(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__o21a_1 _2101_ (.A1(net509),
    .A2(_0819_),
    .B1(net526),
    .X(_0820_));
 sky130_fd_sc_hd__a211o_1 _2102_ (.A1(net456),
    .A2(net525),
    .B1(net538),
    .C1(_0820_),
    .X(_0020_));
 sky130_fd_sc_hd__a221o_4 _2103_ (.A1(net138),
    .A2(net550),
    .B1(net546),
    .B2(net173),
    .C1(net562),
    .X(_0821_));
 sky130_fd_sc_hd__a21o_1 _2104_ (.A1(net49),
    .A2(net554),
    .B1(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__o211a_2 _2105_ (.A1(net14),
    .A2(net559),
    .B1(_0800_),
    .C1(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__o21a_4 _2106_ (.A1(net509),
    .A2(_0823_),
    .B1(net526),
    .X(_0824_));
 sky130_fd_sc_hd__a211o_1 _2107_ (.A1(net457),
    .A2(net524),
    .B1(net537),
    .C1(_0824_),
    .X(_0021_));
 sky130_fd_sc_hd__a221o_4 _2108_ (.A1(net139),
    .A2(net550),
    .B1(net546),
    .B2(net174),
    .C1(net562),
    .X(_0825_));
 sky130_fd_sc_hd__a21o_1 _2109_ (.A1(net50),
    .A2(net554),
    .B1(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__o211a_4 _2110_ (.A1(net15),
    .A2(net559),
    .B1(_0800_),
    .C1(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__o21a_4 _2111_ (.A1(net509),
    .A2(_0827_),
    .B1(net526),
    .X(_0828_));
 sky130_fd_sc_hd__a211o_1 _2112_ (.A1(net458),
    .A2(net524),
    .B1(net537),
    .C1(_0828_),
    .X(_0022_));
 sky130_fd_sc_hd__a221o_1 _2113_ (.A1(net51),
    .A2(net556),
    .B1(net551),
    .B2(net140),
    .C1(net562),
    .X(_0829_));
 sky130_fd_sc_hd__a21o_2 _2114_ (.A1(net175),
    .A2(net547),
    .B1(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__o211a_1 _2115_ (.A1(net16),
    .A2(net560),
    .B1(_0800_),
    .C1(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__o21a_1 _2116_ (.A1(net509),
    .A2(_0831_),
    .B1(net526),
    .X(_0832_));
 sky130_fd_sc_hd__a211o_1 _2117_ (.A1(net459),
    .A2(net525),
    .B1(net538),
    .C1(_0832_),
    .X(_0023_));
 sky130_fd_sc_hd__and3_4 _2118_ (.A(\videoMemory.wbReadReady ),
    .B(net371),
    .C(_0278_),
    .X(_0833_));
 sky130_fd_sc_hd__a221o_1 _2119_ (.A1(net52),
    .A2(net556),
    .B1(net549),
    .B2(net141),
    .C1(net563),
    .X(_0834_));
 sky130_fd_sc_hd__a21o_1 _2120_ (.A1(net176),
    .A2(net545),
    .B1(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__o211a_1 _2121_ (.A1(net17),
    .A2(net560),
    .B1(_0833_),
    .C1(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__o21a_1 _2122_ (.A1(net509),
    .A2(_0836_),
    .B1(net526),
    .X(_0837_));
 sky130_fd_sc_hd__a211o_1 _2123_ (.A1(net460),
    .A2(net525),
    .B1(net538),
    .C1(_0837_),
    .X(_0024_));
 sky130_fd_sc_hd__a221o_4 _2124_ (.A1(net142),
    .A2(net549),
    .B1(net545),
    .B2(net177),
    .C1(net563),
    .X(_0838_));
 sky130_fd_sc_hd__a21o_1 _2125_ (.A1(net53),
    .A2(net553),
    .B1(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__o211a_4 _2126_ (.A1(net18),
    .A2(net558),
    .B1(_0833_),
    .C1(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__o21a_1 _2127_ (.A1(net510),
    .A2(_0840_),
    .B1(net527),
    .X(_0841_));
 sky130_fd_sc_hd__a211o_1 _2128_ (.A1(net461),
    .A2(net523),
    .B1(net536),
    .C1(_0841_),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_4 _2129_ (.A1(net143),
    .A2(net549),
    .B1(net545),
    .B2(net178),
    .X(_0842_));
 sky130_fd_sc_hd__a211o_1 _2130_ (.A1(net54),
    .A2(net553),
    .B1(_0842_),
    .C1(net564),
    .X(_0843_));
 sky130_fd_sc_hd__o211a_4 _2131_ (.A1(net19),
    .A2(net558),
    .B1(_0833_),
    .C1(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__o21a_4 _2132_ (.A1(net510),
    .A2(_0844_),
    .B1(net527),
    .X(_0845_));
 sky130_fd_sc_hd__a211o_1 _2133_ (.A1(net462),
    .A2(net525),
    .B1(net536),
    .C1(_0845_),
    .X(_0026_));
 sky130_fd_sc_hd__a22o_4 _2134_ (.A1(net144),
    .A2(net549),
    .B1(net545),
    .B2(net179),
    .X(_0846_));
 sky130_fd_sc_hd__a211o_1 _2135_ (.A1(net55),
    .A2(net553),
    .B1(_0846_),
    .C1(net564),
    .X(_0847_));
 sky130_fd_sc_hd__o211a_4 _2136_ (.A1(net20),
    .A2(net558),
    .B1(_0833_),
    .C1(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__o21a_2 _2137_ (.A1(net510),
    .A2(_0848_),
    .B1(net527),
    .X(_0849_));
 sky130_fd_sc_hd__a211o_1 _2138_ (.A1(net463),
    .A2(net525),
    .B1(net536),
    .C1(_0849_),
    .X(_0027_));
 sky130_fd_sc_hd__a22o_4 _2139_ (.A1(net145),
    .A2(net549),
    .B1(net545),
    .B2(net181),
    .X(_0850_));
 sky130_fd_sc_hd__a211o_1 _2140_ (.A1(net57),
    .A2(net553),
    .B1(_0850_),
    .C1(net564),
    .X(_0851_));
 sky130_fd_sc_hd__o211a_4 _2141_ (.A1(net21),
    .A2(net558),
    .B1(_0833_),
    .C1(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__o21a_1 _2142_ (.A1(net510),
    .A2(_0852_),
    .B1(net527),
    .X(_0853_));
 sky130_fd_sc_hd__a211o_1 _2143_ (.A1(net464),
    .A2(net522),
    .B1(net536),
    .C1(_0853_),
    .X(_0028_));
 sky130_fd_sc_hd__a221o_4 _2144_ (.A1(net146),
    .A2(net549),
    .B1(net545),
    .B2(net182),
    .C1(net563),
    .X(_0854_));
 sky130_fd_sc_hd__a21o_1 _2145_ (.A1(net58),
    .A2(net553),
    .B1(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__o211a_4 _2146_ (.A1(net22),
    .A2(net558),
    .B1(_0833_),
    .C1(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__o21a_1 _2147_ (.A1(net510),
    .A2(_0856_),
    .B1(net527),
    .X(_0857_));
 sky130_fd_sc_hd__a211o_1 _2148_ (.A1(net465),
    .A2(net523),
    .B1(net536),
    .C1(_0857_),
    .X(_0029_));
 sky130_fd_sc_hd__a221o_4 _2149_ (.A1(net148),
    .A2(net549),
    .B1(net545),
    .B2(net183),
    .C1(net563),
    .X(_0858_));
 sky130_fd_sc_hd__a21o_1 _2150_ (.A1(net59),
    .A2(net553),
    .B1(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__o211a_4 _2151_ (.A1(net24),
    .A2(net558),
    .B1(_0833_),
    .C1(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__o21a_1 _2152_ (.A1(net510),
    .A2(_0860_),
    .B1(net527),
    .X(_0861_));
 sky130_fd_sc_hd__a211o_1 _2153_ (.A1(net467),
    .A2(net522),
    .B1(net536),
    .C1(_0861_),
    .X(_0030_));
 sky130_fd_sc_hd__a221o_1 _2154_ (.A1(net60),
    .A2(net556),
    .B1(net549),
    .B2(net149),
    .C1(net563),
    .X(_0862_));
 sky130_fd_sc_hd__a21o_1 _2155_ (.A1(net184),
    .A2(net545),
    .B1(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__o211a_1 _2156_ (.A1(net25),
    .A2(net560),
    .B1(_0833_),
    .C1(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__o21a_4 _2157_ (.A1(net509),
    .A2(_0864_),
    .B1(net526),
    .X(_0865_));
 sky130_fd_sc_hd__a211o_1 _2158_ (.A1(net468),
    .A2(net524),
    .B1(net536),
    .C1(_0865_),
    .X(_0031_));
 sky130_fd_sc_hd__a21oi_1 _2159_ (.A1(_1330_),
    .A2(_0519_),
    .B1(net538),
    .Y(_0032_));
 sky130_fd_sc_hd__nand2_2 _2160_ (.A(net271),
    .B(net309),
    .Y(_0866_));
 sky130_fd_sc_hd__o31ai_4 _2161_ (.A1(\wbPeripheralBusInterface.state[1] ),
    .A2(net610),
    .A3(_0866_),
    .B1(net538),
    .Y(_0867_));
 sky130_fd_sc_hd__o21a_1 _2162_ (.A1(net476),
    .A2(_1353_),
    .B1(_0867_),
    .X(_0033_));
 sky130_fd_sc_hd__and3b_1 _2163_ (.A_N(_0866_),
    .B(net603),
    .C(_1353_),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_1 _2164_ (.A0(\wbPeripheralBusInterface.currentAddress[2] ),
    .A1(net263),
    .S(net533),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2165_ (.A0(\wbPeripheralBusInterface.currentAddress[3] ),
    .A1(net264),
    .S(net533),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2166_ (.A0(\wbPeripheralBusInterface.currentAddress[4] ),
    .A1(net265),
    .S(net533),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2167_ (.A0(\wbPeripheralBusInterface.currentAddress[5] ),
    .A1(net266),
    .S(net533),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2168_ (.A0(\wbPeripheralBusInterface.currentAddress[6] ),
    .A1(net267),
    .S(net535),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2169_ (.A0(\wbPeripheralBusInterface.currentAddress[7] ),
    .A1(net268),
    .S(net535),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2170_ (.A0(\wbPeripheralBusInterface.currentAddress[8] ),
    .A1(net269),
    .S(net533),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2171_ (.A0(\wbPeripheralBusInterface.currentAddress[9] ),
    .A1(net270),
    .S(net535),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _2172_ (.A0(\wbPeripheralBusInterface.currentAddress[10] ),
    .A1(net249),
    .S(net533),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _2173_ (.A0(\wbPeripheralBusInterface.currentAddress[11] ),
    .A1(net250),
    .S(net534),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _2174_ (.A0(\wbPeripheralBusInterface.currentAddress[12] ),
    .A1(net251),
    .S(net534),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2175_ (.A0(\wbPeripheralBusInterface.currentAddress[13] ),
    .A1(net252),
    .S(net534),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2176_ (.A0(\wbPeripheralBusInterface.currentAddress[14] ),
    .A1(net253),
    .S(net534),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2177_ (.A0(\wbPeripheralBusInterface.currentAddress[15] ),
    .A1(net254),
    .S(net534),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _2178_ (.A0(\wbPeripheralBusInterface.currentAddress[16] ),
    .A1(net255),
    .S(net534),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2179_ (.A0(\wbPeripheralBusInterface.currentAddress[17] ),
    .A1(net256),
    .S(net535),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2180_ (.A0(\wbPeripheralBusInterface.currentAddress[18] ),
    .A1(net257),
    .S(net534),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2181_ (.A0(\wbPeripheralBusInterface.currentAddress[19] ),
    .A1(net258),
    .S(net534),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2182_ (.A0(\wbPeripheralBusInterface.currentAddress[20] ),
    .A1(net259),
    .S(net534),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2183_ (.A0(\wbPeripheralBusInterface.currentAddress[21] ),
    .A1(net260),
    .S(net534),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2184_ (.A0(\wbPeripheralBusInterface.currentAddress[22] ),
    .A1(net261),
    .S(net535),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2185_ (.A0(\wbPeripheralBusInterface.currentAddress[23] ),
    .A1(net262),
    .S(net535),
    .X(_0055_));
 sky130_fd_sc_hd__nor2_1 _2186_ (.A(net611),
    .B(net531),
    .Y(_0056_));
 sky130_fd_sc_hd__o221a_1 _2187_ (.A1(net310),
    .A2(net581),
    .B1(net531),
    .B2(\videoMemory.wbReadReady ),
    .C1(_0867_),
    .X(_0057_));
 sky130_fd_sc_hd__a21boi_1 _2188_ (.A1(net310),
    .A2(_1353_),
    .B1_N(_0867_),
    .Y(_0058_));
 sky130_fd_sc_hd__nor2_1 _2189_ (.A(net614),
    .B(net437),
    .Y(_0060_));
 sky130_fd_sc_hd__nor2_1 _2190_ (.A(net615),
    .B(net440),
    .Y(_0061_));
 sky130_fd_sc_hd__and2_1 _2191_ (.A(\vga.inVerticalVisibleArea ),
    .B(net609),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _2192_ (.A0(net602),
    .A1(net305),
    .S(net533),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _2193_ (.A0(net598),
    .A1(net306),
    .S(net533),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2194_ (.A0(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .A1(net307),
    .S(net533),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2195_ (.A0(\wbPeripheralBusInterface.currentByteSelect[3] ),
    .A1(net308),
    .S(net533),
    .X(_0078_));
 sky130_fd_sc_hd__nand2_1 _2196_ (.A(\vga.raw_verticalPixelStretchCounter[0] ),
    .B(net528),
    .Y(_0869_));
 sky130_fd_sc_hd__or2_1 _2197_ (.A(\vga.raw_verticalPixelStretchCounter[0] ),
    .B(net529),
    .X(_0870_));
 sky130_fd_sc_hd__and3_1 _2198_ (.A(_0345_),
    .B(_0869_),
    .C(_0870_),
    .X(_0079_));
 sky130_fd_sc_hd__xor2_1 _2199_ (.A(\vga.raw_verticalPixelStretchCounter[1] ),
    .B(_0869_),
    .X(_0871_));
 sky130_fd_sc_hd__nor2_1 _2200_ (.A(_0346_),
    .B(_0871_),
    .Y(_0080_));
 sky130_fd_sc_hd__mux2_1 _2201_ (.A0(\vga.raw_verticalPixelStretchCounter[2] ),
    .A1(_0337_),
    .S(net529),
    .X(_0872_));
 sky130_fd_sc_hd__and3_1 _2202_ (.A(net576),
    .B(_0344_),
    .C(_0872_),
    .X(_0081_));
 sky130_fd_sc_hd__nand2_1 _2203_ (.A(net528),
    .B(_0339_),
    .Y(_0873_));
 sky130_fd_sc_hd__o211a_1 _2204_ (.A1(\vga.raw_verticalPixelStretchCounter[3] ),
    .A2(net528),
    .B1(_0345_),
    .C1(_0873_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2205_ (.A0(\vga.raw_subPixelCounter[0] ),
    .A1(\vga.raw_subPixelCounter_buffered[0] ),
    .S(_0283_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2206_ (.A0(\vga.raw_subPixelCounter[1] ),
    .A1(\vga.raw_subPixelCounter_buffered[1] ),
    .S(_0283_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2207_ (.A0(\vga.raw_subPixelCounter[2] ),
    .A1(\vga.raw_subPixelCounter_buffered[2] ),
    .S(_0283_),
    .X(_0085_));
 sky130_fd_sc_hd__a31o_1 _2208_ (.A1(\vga.raw_verticalPixelCounter[5] ),
    .A2(\vga.raw_verticalPixelCounter[6] ),
    .A3(_0362_),
    .B1(\vga.raw_verticalPixelCounter[7] ),
    .X(_0874_));
 sky130_fd_sc_hd__and3_2 _2209_ (.A(\vga.raw_verticalPixelCounter[6] ),
    .B(\vga.raw_verticalPixelCounter[7] ),
    .C(_0363_),
    .X(_0875_));
 sky130_fd_sc_hd__and3b_1 _2210_ (.A_N(_0875_),
    .B(net576),
    .C(_0874_),
    .X(_0093_));
 sky130_fd_sc_hd__a21oi_1 _2211_ (.A1(\vga.raw_verticalPixelCounter[8] ),
    .A2(_0875_),
    .B1(net532),
    .Y(_0876_));
 sky130_fd_sc_hd__o21a_1 _2212_ (.A1(\vga.raw_verticalPixelCounter[8] ),
    .A2(_0875_),
    .B1(_0876_),
    .X(_0094_));
 sky130_fd_sc_hd__a21oi_1 _2213_ (.A1(\vga.raw_verticalPixelCounter[8] ),
    .A2(_0875_),
    .B1(\vga.raw_verticalPixelCounter[9] ),
    .Y(_0877_));
 sky130_fd_sc_hd__a31o_1 _2214_ (.A1(\vga.raw_verticalPixelCounter[8] ),
    .A2(\vga.raw_verticalPixelCounter[9] ),
    .A3(_0875_),
    .B1(net532),
    .X(_0878_));
 sky130_fd_sc_hd__nor2_1 _2215_ (.A(_0877_),
    .B(_0878_),
    .Y(_0095_));
 sky130_fd_sc_hd__nor2_1 _2216_ (.A(_1329_),
    .B(_0299_),
    .Y(_0879_));
 sky130_fd_sc_hd__a211o_1 _2217_ (.A1(_1329_),
    .A2(_0299_),
    .B1(_0287_),
    .C1(_0286_),
    .X(_0880_));
 sky130_fd_sc_hd__nor2_1 _2218_ (.A(_0879_),
    .B(_0880_),
    .Y(_0096_));
 sky130_fd_sc_hd__and2_1 _2219_ (.A(\vga.raw_subPixelCounter[1] ),
    .B(_0879_),
    .X(_0881_));
 sky130_fd_sc_hd__o21ai_1 _2220_ (.A1(\vga.raw_subPixelCounter[1] ),
    .A2(_0879_),
    .B1(_0285_),
    .Y(_0882_));
 sky130_fd_sc_hd__nor2_1 _2221_ (.A(_0881_),
    .B(_0882_),
    .Y(_0097_));
 sky130_fd_sc_hd__o21ai_1 _2222_ (.A1(\vga.raw_subPixelCounter[2] ),
    .A2(_0881_),
    .B1(_0306_),
    .Y(_0883_));
 sky130_fd_sc_hd__a21oi_1 _2223_ (.A1(\vga.raw_subPixelCounter[2] ),
    .A2(_0881_),
    .B1(_0883_),
    .Y(_0098_));
 sky130_fd_sc_hd__and2_1 _2224_ (.A(\vga.hsync ),
    .B(net603),
    .X(_0108_));
 sky130_fd_sc_hd__and2_1 _2225_ (.A(\vga.vsync ),
    .B(net604),
    .X(_0109_));
 sky130_fd_sc_hd__nand2_2 _2226_ (.A(_0285_),
    .B(_0299_),
    .Y(_0884_));
 sky130_fd_sc_hd__nor2_1 _2227_ (.A(\vga.raw_horizontalPixelStretchCounter[0] ),
    .B(_0884_),
    .Y(_0110_));
 sky130_fd_sc_hd__nor2_1 _2228_ (.A(_0291_),
    .B(_0884_),
    .Y(_0111_));
 sky130_fd_sc_hd__and4_1 _2229_ (.A(_0285_),
    .B(_0288_),
    .C(_0295_),
    .D(_0299_),
    .X(_0112_));
 sky130_fd_sc_hd__nor2_1 _2230_ (.A(_0289_),
    .B(_0884_),
    .Y(_0113_));
 sky130_fd_sc_hd__and4_1 _2231_ (.A(net212),
    .B(net493),
    .C(net501),
    .D(net491),
    .X(_0885_));
 sky130_fd_sc_hd__and2_1 _2232_ (.A(net189),
    .B(net481),
    .X(_0886_));
 sky130_fd_sc_hd__o22a_1 _2233_ (.A1(net497),
    .A2(net505),
    .B1(_0474_),
    .B2(net88),
    .X(_0887_));
 sky130_fd_sc_hd__o32a_1 _2234_ (.A1(_0885_),
    .A2(_0886_),
    .A3(_0887_),
    .B1(net477),
    .B2(net65),
    .X(_0888_));
 sky130_fd_sc_hd__or2_1 _2235_ (.A(net591),
    .B(\vga.currentPixelData[0] ),
    .X(_0889_));
 sky130_fd_sc_hd__o211a_1 _2236_ (.A1(net587),
    .A2(_0888_),
    .B1(_0889_),
    .C1(net539),
    .X(_0114_));
 sky130_fd_sc_hd__and4_1 _2237_ (.A(net213),
    .B(net493),
    .C(net501),
    .D(net491),
    .X(_0890_));
 sky130_fd_sc_hd__and2_1 _2238_ (.A(net200),
    .B(net481),
    .X(_0891_));
 sky130_fd_sc_hd__o22a_2 _2239_ (.A1(net497),
    .A2(net505),
    .B1(net483),
    .B2(net89),
    .X(_0892_));
 sky130_fd_sc_hd__o32a_1 _2240_ (.A1(_0890_),
    .A2(_0891_),
    .A3(_0892_),
    .B1(net477),
    .B2(net76),
    .X(_0893_));
 sky130_fd_sc_hd__or2_1 _2241_ (.A(net591),
    .B(\vga.currentPixelData[1] ),
    .X(_0894_));
 sky130_fd_sc_hd__o211a_1 _2242_ (.A1(net587),
    .A2(_0893_),
    .B1(_0894_),
    .C1(net539),
    .X(_0115_));
 sky130_fd_sc_hd__and4_1 _2243_ (.A(net214),
    .B(net493),
    .C(net501),
    .D(net492),
    .X(_0895_));
 sky130_fd_sc_hd__and2_1 _2244_ (.A(net211),
    .B(net481),
    .X(_0896_));
 sky130_fd_sc_hd__o22a_1 _2245_ (.A1(net497),
    .A2(net505),
    .B1(_0474_),
    .B2(net90),
    .X(_0897_));
 sky130_fd_sc_hd__o32a_1 _2246_ (.A1(_0895_),
    .A2(_0896_),
    .A3(_0897_),
    .B1(net477),
    .B2(net87),
    .X(_0898_));
 sky130_fd_sc_hd__or2_1 _2247_ (.A(net591),
    .B(\vga.currentPixelData[2] ),
    .X(_0899_));
 sky130_fd_sc_hd__o211a_1 _2248_ (.A1(net587),
    .A2(_0898_),
    .B1(_0899_),
    .C1(net539),
    .X(_0116_));
 sky130_fd_sc_hd__and4_1 _2249_ (.A(net215),
    .B(net496),
    .C(net504),
    .D(net491),
    .X(_0900_));
 sky130_fd_sc_hd__and2_1 _2250_ (.A(net220),
    .B(net481),
    .X(_0901_));
 sky130_fd_sc_hd__o22a_2 _2251_ (.A1(net497),
    .A2(net505),
    .B1(net483),
    .B2(net91),
    .X(_0902_));
 sky130_fd_sc_hd__o32a_1 _2252_ (.A1(_0900_),
    .A2(_0901_),
    .A3(_0902_),
    .B1(net477),
    .B2(net96),
    .X(_0903_));
 sky130_fd_sc_hd__or2_1 _2253_ (.A(net591),
    .B(\vga.currentPixelData[3] ),
    .X(_0904_));
 sky130_fd_sc_hd__o211a_1 _2254_ (.A1(net587),
    .A2(_0903_),
    .B1(_0904_),
    .C1(net539),
    .X(_0117_));
 sky130_fd_sc_hd__and4_1 _2255_ (.A(net216),
    .B(net493),
    .C(net501),
    .D(net492),
    .X(_0905_));
 sky130_fd_sc_hd__and2_1 _2256_ (.A(net231),
    .B(net481),
    .X(_0906_));
 sky130_fd_sc_hd__o22a_1 _2257_ (.A1(net497),
    .A2(net505),
    .B1(net484),
    .B2(net92),
    .X(_0907_));
 sky130_fd_sc_hd__o32a_1 _2258_ (.A1(_0905_),
    .A2(_0906_),
    .A3(_0907_),
    .B1(net477),
    .B2(net107),
    .X(_0908_));
 sky130_fd_sc_hd__or2_1 _2259_ (.A(net591),
    .B(\vga.currentPixelData[4] ),
    .X(_0909_));
 sky130_fd_sc_hd__o211a_1 _2260_ (.A1(net587),
    .A2(_0908_),
    .B1(_0909_),
    .C1(net539),
    .X(_0118_));
 sky130_fd_sc_hd__and4_1 _2261_ (.A(net217),
    .B(net493),
    .C(net501),
    .D(net492),
    .X(_0910_));
 sky130_fd_sc_hd__and2_1 _2262_ (.A(net242),
    .B(net481),
    .X(_0911_));
 sky130_fd_sc_hd__o22a_2 _2263_ (.A1(net497),
    .A2(net505),
    .B1(net483),
    .B2(net93),
    .X(_0912_));
 sky130_fd_sc_hd__o32a_1 _2264_ (.A1(_0910_),
    .A2(_0911_),
    .A3(_0912_),
    .B1(net477),
    .B2(net118),
    .X(_0913_));
 sky130_fd_sc_hd__or2_1 _2265_ (.A(net591),
    .B(\vga.currentPixelData[5] ),
    .X(_0914_));
 sky130_fd_sc_hd__o211a_1 _2266_ (.A1(net587),
    .A2(_0913_),
    .B1(_0914_),
    .C1(net539),
    .X(_0119_));
 sky130_fd_sc_hd__and4_1 _2267_ (.A(net218),
    .B(net493),
    .C(net501),
    .D(net492),
    .X(_0915_));
 sky130_fd_sc_hd__and2_1 _2268_ (.A(net245),
    .B(net481),
    .X(_0916_));
 sky130_fd_sc_hd__o22a_1 _2269_ (.A1(net497),
    .A2(net505),
    .B1(net483),
    .B2(net94),
    .X(_0917_));
 sky130_fd_sc_hd__o32a_1 _2270_ (.A1(_0915_),
    .A2(_0916_),
    .A3(_0917_),
    .B1(net480),
    .B2(net121),
    .X(_0918_));
 sky130_fd_sc_hd__or2_1 _2271_ (.A(net591),
    .B(\vga.currentPixelData[6] ),
    .X(_0919_));
 sky130_fd_sc_hd__o211a_1 _2272_ (.A1(net587),
    .A2(_0918_),
    .B1(_0919_),
    .C1(net539),
    .X(_0120_));
 sky130_fd_sc_hd__and4_1 _2273_ (.A(net219),
    .B(net493),
    .C(net501),
    .D(net492),
    .X(_0920_));
 sky130_fd_sc_hd__and2_1 _2274_ (.A(net246),
    .B(net481),
    .X(_0921_));
 sky130_fd_sc_hd__o22a_1 _2275_ (.A1(net497),
    .A2(net505),
    .B1(net484),
    .B2(net95),
    .X(_0922_));
 sky130_fd_sc_hd__o32a_1 _2276_ (.A1(_0920_),
    .A2(_0921_),
    .A3(_0922_),
    .B1(net480),
    .B2(net122),
    .X(_0923_));
 sky130_fd_sc_hd__or2_1 _2277_ (.A(net591),
    .B(\vga.currentPixelData[7] ),
    .X(_0924_));
 sky130_fd_sc_hd__o211a_1 _2278_ (.A1(net587),
    .A2(_0923_),
    .B1(_0924_),
    .C1(net539),
    .X(_0121_));
 sky130_fd_sc_hd__and4_1 _2279_ (.A(net221),
    .B(net495),
    .C(net503),
    .D(net491),
    .X(_0925_));
 sky130_fd_sc_hd__and2_1 _2280_ (.A(net247),
    .B(net481),
    .X(_0926_));
 sky130_fd_sc_hd__o22a_1 _2281_ (.A1(net498),
    .A2(net506),
    .B1(net484),
    .B2(net97),
    .X(_0927_));
 sky130_fd_sc_hd__o32a_1 _2282_ (.A1(_0925_),
    .A2(_0926_),
    .A3(_0927_),
    .B1(net477),
    .B2(net123),
    .X(_0928_));
 sky130_fd_sc_hd__or2_1 _2283_ (.A(net594),
    .B(\vga.currentPixelData[8] ),
    .X(_0929_));
 sky130_fd_sc_hd__o211a_1 _2284_ (.A1(net588),
    .A2(_0928_),
    .B1(_0929_),
    .C1(net540),
    .X(_0122_));
 sky130_fd_sc_hd__and4_1 _2285_ (.A(net222),
    .B(net493),
    .C(net501),
    .D(net491),
    .X(_0930_));
 sky130_fd_sc_hd__and2_1 _2286_ (.A(net248),
    .B(net482),
    .X(_0931_));
 sky130_fd_sc_hd__o22a_1 _2287_ (.A1(net498),
    .A2(net506),
    .B1(net483),
    .B2(net98),
    .X(_0932_));
 sky130_fd_sc_hd__o32a_1 _2288_ (.A1(_0930_),
    .A2(_0931_),
    .A3(_0932_),
    .B1(net477),
    .B2(net124),
    .X(_0933_));
 sky130_fd_sc_hd__or2_1 _2289_ (.A(net594),
    .B(\vga.currentPixelData[9] ),
    .X(_0934_));
 sky130_fd_sc_hd__o211a_1 _2290_ (.A1(net588),
    .A2(_0933_),
    .B1(_0934_),
    .C1(net540),
    .X(_0123_));
 sky130_fd_sc_hd__and4_1 _2291_ (.A(net223),
    .B(net495),
    .C(net503),
    .D(net491),
    .X(_0935_));
 sky130_fd_sc_hd__and2_1 _2292_ (.A(net190),
    .B(net487),
    .X(_0936_));
 sky130_fd_sc_hd__o22a_1 _2293_ (.A1(net498),
    .A2(net506),
    .B1(net484),
    .B2(net99),
    .X(_0937_));
 sky130_fd_sc_hd__o32a_1 _2294_ (.A1(_0935_),
    .A2(_0936_),
    .A3(_0937_),
    .B1(net479),
    .B2(net66),
    .X(_0938_));
 sky130_fd_sc_hd__or2_1 _2295_ (.A(net593),
    .B(\vga.currentPixelData[10] ),
    .X(_0939_));
 sky130_fd_sc_hd__o211a_1 _2296_ (.A1(net590),
    .A2(_0938_),
    .B1(_0939_),
    .C1(net540),
    .X(_0124_));
 sky130_fd_sc_hd__and4_1 _2297_ (.A(net224),
    .B(net495),
    .C(net503),
    .D(net489),
    .X(_0940_));
 sky130_fd_sc_hd__and2_1 _2298_ (.A(net191),
    .B(net487),
    .X(_0941_));
 sky130_fd_sc_hd__o22a_1 _2299_ (.A1(net498),
    .A2(net506),
    .B1(net483),
    .B2(net100),
    .X(_0942_));
 sky130_fd_sc_hd__o32a_1 _2300_ (.A1(_0940_),
    .A2(_0941_),
    .A3(_0942_),
    .B1(net479),
    .B2(net67),
    .X(_0943_));
 sky130_fd_sc_hd__or2_1 _2301_ (.A(net592),
    .B(\vga.currentPixelData[11] ),
    .X(_0944_));
 sky130_fd_sc_hd__o211a_1 _2302_ (.A1(net589),
    .A2(_0943_),
    .B1(_0944_),
    .C1(net541),
    .X(_0125_));
 sky130_fd_sc_hd__and4_1 _2303_ (.A(net225),
    .B(net495),
    .C(net503),
    .D(net490),
    .X(_0945_));
 sky130_fd_sc_hd__and2_1 _2304_ (.A(net192),
    .B(net481),
    .X(_0946_));
 sky130_fd_sc_hd__o22a_1 _2305_ (.A1(net498),
    .A2(net506),
    .B1(net484),
    .B2(net101),
    .X(_0947_));
 sky130_fd_sc_hd__o32a_1 _2306_ (.A1(_0945_),
    .A2(_0946_),
    .A3(_0947_),
    .B1(net480),
    .B2(net68),
    .X(_0948_));
 sky130_fd_sc_hd__or2_1 _2307_ (.A(net591),
    .B(\vga.currentPixelData[12] ),
    .X(_0949_));
 sky130_fd_sc_hd__o211a_1 _2308_ (.A1(net587),
    .A2(_0948_),
    .B1(_0949_),
    .C1(net539),
    .X(_0126_));
 sky130_fd_sc_hd__and4_1 _2309_ (.A(net226),
    .B(net495),
    .C(net503),
    .D(net489),
    .X(_0950_));
 sky130_fd_sc_hd__and2_1 _2310_ (.A(net193),
    .B(net482),
    .X(_0951_));
 sky130_fd_sc_hd__o22a_1 _2311_ (.A1(net498),
    .A2(net506),
    .B1(net483),
    .B2(net102),
    .X(_0952_));
 sky130_fd_sc_hd__o32a_1 _2312_ (.A1(_0950_),
    .A2(_0951_),
    .A3(_0952_),
    .B1(net480),
    .B2(net69),
    .X(_0953_));
 sky130_fd_sc_hd__or2_1 _2313_ (.A(net591),
    .B(\vga.currentPixelData[13] ),
    .X(_0954_));
 sky130_fd_sc_hd__o211a_1 _2314_ (.A1(net587),
    .A2(_0953_),
    .B1(_0954_),
    .C1(net540),
    .X(_0127_));
 sky130_fd_sc_hd__and4_1 _2315_ (.A(net227),
    .B(net495),
    .C(net503),
    .D(net490),
    .X(_0955_));
 sky130_fd_sc_hd__and2_1 _2316_ (.A(net194),
    .B(net482),
    .X(_0956_));
 sky130_fd_sc_hd__o22a_1 _2317_ (.A1(net497),
    .A2(net505),
    .B1(net483),
    .B2(net103),
    .X(_0957_));
 sky130_fd_sc_hd__o32a_1 _2318_ (.A1(_0955_),
    .A2(_0956_),
    .A3(_0957_),
    .B1(net479),
    .B2(net70),
    .X(_0958_));
 sky130_fd_sc_hd__or2_1 _2319_ (.A(net594),
    .B(\vga.currentPixelData[14] ),
    .X(_0959_));
 sky130_fd_sc_hd__o211a_1 _2320_ (.A1(net588),
    .A2(_0958_),
    .B1(_0959_),
    .C1(net540),
    .X(_0128_));
 sky130_fd_sc_hd__and4_1 _2321_ (.A(net228),
    .B(net495),
    .C(net503),
    .D(net489),
    .X(_0960_));
 sky130_fd_sc_hd__and2_1 _2322_ (.A(net195),
    .B(net482),
    .X(_0961_));
 sky130_fd_sc_hd__o22a_1 _2323_ (.A1(net499),
    .A2(net507),
    .B1(net483),
    .B2(net104),
    .X(_0962_));
 sky130_fd_sc_hd__o32a_1 _2324_ (.A1(_0960_),
    .A2(_0961_),
    .A3(_0962_),
    .B1(net477),
    .B2(net71),
    .X(_0963_));
 sky130_fd_sc_hd__or2_1 _2325_ (.A(net594),
    .B(\vga.currentPixelData[15] ),
    .X(_0964_));
 sky130_fd_sc_hd__o211a_1 _2326_ (.A1(net588),
    .A2(_0963_),
    .B1(_0964_),
    .C1(net540),
    .X(_0129_));
 sky130_fd_sc_hd__and4_1 _2327_ (.A(net229),
    .B(net495),
    .C(net503),
    .D(net491),
    .X(_0965_));
 sky130_fd_sc_hd__and2_1 _2328_ (.A(net196),
    .B(net482),
    .X(_0966_));
 sky130_fd_sc_hd__o22a_1 _2329_ (.A1(net497),
    .A2(net505),
    .B1(net483),
    .B2(net105),
    .X(_0967_));
 sky130_fd_sc_hd__o32a_1 _2330_ (.A1(_0965_),
    .A2(_0966_),
    .A3(_0967_),
    .B1(net479),
    .B2(net72),
    .X(_0968_));
 sky130_fd_sc_hd__or2_1 _2331_ (.A(net593),
    .B(\vga.currentPixelData[16] ),
    .X(_0969_));
 sky130_fd_sc_hd__o211a_1 _2332_ (.A1(net588),
    .A2(_0968_),
    .B1(_0969_),
    .C1(net540),
    .X(_0130_));
 sky130_fd_sc_hd__and4_1 _2333_ (.A(net230),
    .B(net494),
    .C(net502),
    .D(net489),
    .X(_0970_));
 sky130_fd_sc_hd__and2_1 _2334_ (.A(net197),
    .B(net482),
    .X(_0971_));
 sky130_fd_sc_hd__o22a_1 _2335_ (.A1(net499),
    .A2(net507),
    .B1(net485),
    .B2(net106),
    .X(_0972_));
 sky130_fd_sc_hd__o32a_1 _2336_ (.A1(_0970_),
    .A2(_0971_),
    .A3(_0972_),
    .B1(net479),
    .B2(net73),
    .X(_0973_));
 sky130_fd_sc_hd__or2_1 _2337_ (.A(net592),
    .B(\vga.currentPixelData[17] ),
    .X(_0974_));
 sky130_fd_sc_hd__o211a_1 _2338_ (.A1(net589),
    .A2(_0973_),
    .B1(_0974_),
    .C1(net541),
    .X(_0131_));
 sky130_fd_sc_hd__and4_1 _2339_ (.A(net232),
    .B(net496),
    .C(net504),
    .D(net490),
    .X(_0975_));
 sky130_fd_sc_hd__and2_2 _2340_ (.A(net198),
    .B(net482),
    .X(_0976_));
 sky130_fd_sc_hd__o22a_1 _2341_ (.A1(net499),
    .A2(net507),
    .B1(net485),
    .B2(net108),
    .X(_0977_));
 sky130_fd_sc_hd__o32a_1 _2342_ (.A1(_0975_),
    .A2(_0976_),
    .A3(_0977_),
    .B1(net478),
    .B2(net74),
    .X(_0978_));
 sky130_fd_sc_hd__or2_1 _2343_ (.A(net592),
    .B(\vga.currentPixelData[18] ),
    .X(_0979_));
 sky130_fd_sc_hd__o211a_1 _2344_ (.A1(net589),
    .A2(_0978_),
    .B1(_0979_),
    .C1(net541),
    .X(_0132_));
 sky130_fd_sc_hd__and4_1 _2345_ (.A(net233),
    .B(net496),
    .C(net504),
    .D(net490),
    .X(_0980_));
 sky130_fd_sc_hd__and2_1 _2346_ (.A(net199),
    .B(net487),
    .X(_0981_));
 sky130_fd_sc_hd__o22a_1 _2347_ (.A1(net499),
    .A2(net507),
    .B1(net485),
    .B2(net109),
    .X(_0982_));
 sky130_fd_sc_hd__o32a_1 _2348_ (.A1(_0980_),
    .A2(_0981_),
    .A3(_0982_),
    .B1(net478),
    .B2(net75),
    .X(_0983_));
 sky130_fd_sc_hd__or2_1 _2349_ (.A(net593),
    .B(\vga.currentPixelData[19] ),
    .X(_0984_));
 sky130_fd_sc_hd__o211a_1 _2350_ (.A1(net590),
    .A2(_0983_),
    .B1(_0984_),
    .C1(net542),
    .X(_0133_));
 sky130_fd_sc_hd__and4_1 _2351_ (.A(net234),
    .B(net494),
    .C(net502),
    .D(net489),
    .X(_0985_));
 sky130_fd_sc_hd__and2_1 _2352_ (.A(net201),
    .B(net487),
    .X(_0986_));
 sky130_fd_sc_hd__o22a_1 _2353_ (.A1(net499),
    .A2(net507),
    .B1(net485),
    .B2(net110),
    .X(_0987_));
 sky130_fd_sc_hd__o32a_1 _2354_ (.A1(_0985_),
    .A2(_0986_),
    .A3(_0987_),
    .B1(net478),
    .B2(net77),
    .X(_0988_));
 sky130_fd_sc_hd__or2_1 _2355_ (.A(net592),
    .B(\vga.currentPixelData[20] ),
    .X(_0989_));
 sky130_fd_sc_hd__o211a_1 _2356_ (.A1(net589),
    .A2(_0988_),
    .B1(_0989_),
    .C1(net541),
    .X(_0134_));
 sky130_fd_sc_hd__and4_1 _2357_ (.A(net235),
    .B(net494),
    .C(net502),
    .D(net490),
    .X(_0990_));
 sky130_fd_sc_hd__and2_1 _2358_ (.A(net202),
    .B(net487),
    .X(_0991_));
 sky130_fd_sc_hd__o22a_1 _2359_ (.A1(net499),
    .A2(net507),
    .B1(net485),
    .B2(net111),
    .X(_0992_));
 sky130_fd_sc_hd__o32a_2 _2360_ (.A1(_0990_),
    .A2(_0991_),
    .A3(_0992_),
    .B1(net478),
    .B2(net78),
    .X(_0993_));
 sky130_fd_sc_hd__or2_1 _2361_ (.A(net592),
    .B(\vga.currentPixelData[21] ),
    .X(_0994_));
 sky130_fd_sc_hd__o211a_1 _2362_ (.A1(net589),
    .A2(_0993_),
    .B1(_0994_),
    .C1(net541),
    .X(_0135_));
 sky130_fd_sc_hd__and4_1 _2363_ (.A(net236),
    .B(net495),
    .C(net503),
    .D(net489),
    .X(_0995_));
 sky130_fd_sc_hd__and2_1 _2364_ (.A(net203),
    .B(net487),
    .X(_0996_));
 sky130_fd_sc_hd__o22a_1 _2365_ (.A1(net500),
    .A2(net508),
    .B1(net486),
    .B2(net112),
    .X(_0997_));
 sky130_fd_sc_hd__o32a_1 _2366_ (.A1(_0995_),
    .A2(_0996_),
    .A3(_0997_),
    .B1(net478),
    .B2(net79),
    .X(_0998_));
 sky130_fd_sc_hd__or2_1 _2367_ (.A(net592),
    .B(\vga.currentPixelData[22] ),
    .X(_0999_));
 sky130_fd_sc_hd__o211a_1 _2368_ (.A1(net589),
    .A2(_0998_),
    .B1(_0999_),
    .C1(net541),
    .X(_0136_));
 sky130_fd_sc_hd__and4_1 _2369_ (.A(net237),
    .B(net494),
    .C(net502),
    .D(net490),
    .X(_1000_));
 sky130_fd_sc_hd__and2_1 _2370_ (.A(net204),
    .B(net487),
    .X(_1001_));
 sky130_fd_sc_hd__o22a_1 _2371_ (.A1(net500),
    .A2(net508),
    .B1(net485),
    .B2(net113),
    .X(_1002_));
 sky130_fd_sc_hd__o32a_1 _2372_ (.A1(_1000_),
    .A2(_1001_),
    .A3(_1002_),
    .B1(net478),
    .B2(net80),
    .X(_1003_));
 sky130_fd_sc_hd__or2_1 _2373_ (.A(net592),
    .B(\vga.currentPixelData[23] ),
    .X(_1004_));
 sky130_fd_sc_hd__o211a_1 _2374_ (.A1(net590),
    .A2(_1003_),
    .B1(_1004_),
    .C1(net542),
    .X(_0137_));
 sky130_fd_sc_hd__and4_1 _2375_ (.A(net238),
    .B(net494),
    .C(net502),
    .D(net489),
    .X(_1005_));
 sky130_fd_sc_hd__and2_1 _2376_ (.A(net205),
    .B(net487),
    .X(_1006_));
 sky130_fd_sc_hd__o22a_1 _2377_ (.A1(net500),
    .A2(net508),
    .B1(net485),
    .B2(net114),
    .X(_1007_));
 sky130_fd_sc_hd__o32a_1 _2378_ (.A1(_1005_),
    .A2(_1006_),
    .A3(_1007_),
    .B1(net478),
    .B2(net81),
    .X(_1008_));
 sky130_fd_sc_hd__or2_1 _2379_ (.A(net592),
    .B(\vga.currentPixelData[24] ),
    .X(_1009_));
 sky130_fd_sc_hd__o211a_1 _2380_ (.A1(net589),
    .A2(_1008_),
    .B1(_1009_),
    .C1(net541),
    .X(_0138_));
 sky130_fd_sc_hd__and4_1 _2381_ (.A(net239),
    .B(net494),
    .C(net502),
    .D(net490),
    .X(_1010_));
 sky130_fd_sc_hd__and2_1 _2382_ (.A(net206),
    .B(net487),
    .X(_1011_));
 sky130_fd_sc_hd__o22a_1 _2383_ (.A1(net500),
    .A2(net508),
    .B1(net485),
    .B2(net115),
    .X(_1012_));
 sky130_fd_sc_hd__o32a_1 _2384_ (.A1(_1010_),
    .A2(_1011_),
    .A3(_1012_),
    .B1(net478),
    .B2(net82),
    .X(_1013_));
 sky130_fd_sc_hd__or2_1 _2385_ (.A(net592),
    .B(\vga.currentPixelData[25] ),
    .X(_1014_));
 sky130_fd_sc_hd__o211a_1 _2386_ (.A1(net589),
    .A2(_1013_),
    .B1(_1014_),
    .C1(net542),
    .X(_0139_));
 sky130_fd_sc_hd__and4_1 _2387_ (.A(net240),
    .B(net494),
    .C(net502),
    .D(net489),
    .X(_1015_));
 sky130_fd_sc_hd__and2_1 _2388_ (.A(net207),
    .B(net487),
    .X(_1016_));
 sky130_fd_sc_hd__o22a_1 _2389_ (.A1(net499),
    .A2(net507),
    .B1(net485),
    .B2(net116),
    .X(_1017_));
 sky130_fd_sc_hd__o32a_1 _2390_ (.A1(_1015_),
    .A2(_1016_),
    .A3(_1017_),
    .B1(net478),
    .B2(net83),
    .X(_1018_));
 sky130_fd_sc_hd__or2_1 _2391_ (.A(net593),
    .B(\vga.currentPixelData[26] ),
    .X(_1019_));
 sky130_fd_sc_hd__o211a_1 _2392_ (.A1(net589),
    .A2(_1018_),
    .B1(_1019_),
    .C1(net542),
    .X(_0140_));
 sky130_fd_sc_hd__and4_1 _2393_ (.A(net241),
    .B(net494),
    .C(net502),
    .D(net489),
    .X(_1020_));
 sky130_fd_sc_hd__and2_1 _2394_ (.A(net208),
    .B(net488),
    .X(_1021_));
 sky130_fd_sc_hd__o22a_1 _2395_ (.A1(net499),
    .A2(net507),
    .B1(net485),
    .B2(net117),
    .X(_1022_));
 sky130_fd_sc_hd__o32a_1 _2396_ (.A1(_1020_),
    .A2(_1021_),
    .A3(_1022_),
    .B1(net479),
    .B2(net84),
    .X(_1023_));
 sky130_fd_sc_hd__or2_1 _2397_ (.A(net593),
    .B(\vga.currentPixelData[27] ),
    .X(_1024_));
 sky130_fd_sc_hd__o211a_1 _2398_ (.A1(net590),
    .A2(_1023_),
    .B1(_1024_),
    .C1(net541),
    .X(_0141_));
 sky130_fd_sc_hd__and4_1 _2399_ (.A(net243),
    .B(net494),
    .C(net502),
    .D(net489),
    .X(_1025_));
 sky130_fd_sc_hd__and2_1 _2400_ (.A(net209),
    .B(net488),
    .X(_1026_));
 sky130_fd_sc_hd__o22a_1 _2401_ (.A1(net499),
    .A2(net507),
    .B1(net486),
    .B2(net119),
    .X(_1027_));
 sky130_fd_sc_hd__o32a_1 _2402_ (.A1(_1025_),
    .A2(_1026_),
    .A3(_1027_),
    .B1(net478),
    .B2(net85),
    .X(_1028_));
 sky130_fd_sc_hd__or2_1 _2403_ (.A(net593),
    .B(\vga.currentPixelData[28] ),
    .X(_1029_));
 sky130_fd_sc_hd__o211a_1 _2404_ (.A1(net590),
    .A2(_1028_),
    .B1(_1029_),
    .C1(net541),
    .X(_0142_));
 sky130_fd_sc_hd__and4_1 _2405_ (.A(net244),
    .B(net494),
    .C(net502),
    .D(net490),
    .X(_1030_));
 sky130_fd_sc_hd__and2_1 _2406_ (.A(net210),
    .B(net488),
    .X(_1031_));
 sky130_fd_sc_hd__o22a_1 _2407_ (.A1(net499),
    .A2(net507),
    .B1(net486),
    .B2(net120),
    .X(_1032_));
 sky130_fd_sc_hd__o32a_1 _2408_ (.A1(_1030_),
    .A2(_1031_),
    .A3(_1032_),
    .B1(net479),
    .B2(net86),
    .X(_1033_));
 sky130_fd_sc_hd__or2_1 _2409_ (.A(\vga.currentPixelData[29] ),
    .B(net592),
    .X(_1034_));
 sky130_fd_sc_hd__o211a_1 _2410_ (.A1(net589),
    .A2(_1033_),
    .B1(_1034_),
    .C1(net541),
    .X(_0143_));
 sky130_fd_sc_hd__xnor2_1 _2411_ (.A(\vga.horizontalWholeLineCompare[8] ),
    .B(\vga.horizontalCounter[8] ),
    .Y(_1035_));
 sky130_fd_sc_hd__xnor2_1 _2412_ (.A(\vga.horizontalWholeLineCompare[3] ),
    .B(\vga.horizontalCounter[3] ),
    .Y(_1036_));
 sky130_fd_sc_hd__xnor2_1 _2413_ (.A(\vga.horizontalWholeLineCompare[9] ),
    .B(\vga.horizontalCounter[9] ),
    .Y(_1037_));
 sky130_fd_sc_hd__or2_1 _2414_ (.A(\vga.horizontalWholeLineCompare[1] ),
    .B(\vga.horizontalCounter[1] ),
    .X(_1038_));
 sky130_fd_sc_hd__nand2_1 _2415_ (.A(\vga.horizontalWholeLineCompare[1] ),
    .B(\vga.horizontalCounter[1] ),
    .Y(_1039_));
 sky130_fd_sc_hd__a22o_1 _2416_ (.A1(\vga.horizontalWholeLineCompare[0] ),
    .A2(_1332_),
    .B1(\vga.horizontalCounter[5] ),
    .B2(_1305_),
    .X(_1040_));
 sky130_fd_sc_hd__a221o_1 _2417_ (.A1(_1306_),
    .A2(\vga.horizontalCounter[6] ),
    .B1(_1339_),
    .B2(\vga.horizontalWholeLineCompare[7] ),
    .C1(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__o221a_1 _2418_ (.A1(\vga.horizontalWholeLineCompare[2] ),
    .A2(_1334_),
    .B1(\vga.horizontalCounter[5] ),
    .B2(_1305_),
    .C1(_1037_),
    .X(_1042_));
 sky130_fd_sc_hd__o22a_1 _2419_ (.A1(\vga.horizontalWholeLineCompare[4] ),
    .A2(_1336_),
    .B1(_1339_),
    .B2(\vga.horizontalWholeLineCompare[7] ),
    .X(_1043_));
 sky130_fd_sc_hd__a22o_1 _2420_ (.A1(\vga.horizontalWholeLineCompare[2] ),
    .A2(_1334_),
    .B1(_1336_),
    .B2(\vga.horizontalWholeLineCompare[4] ),
    .X(_1044_));
 sky130_fd_sc_hd__a22o_1 _2421_ (.A1(\vga.horizontalWholeLineCompare[6] ),
    .A2(_1338_),
    .B1(_1342_),
    .B2(\vga.horizontalWholeLineCompare[10] ),
    .X(_1045_));
 sky130_fd_sc_hd__a21oi_1 _2422_ (.A1(_1038_),
    .A2(_1039_),
    .B1(_1041_),
    .Y(_1046_));
 sky130_fd_sc_hd__o221a_1 _2423_ (.A1(\vga.horizontalWholeLineCompare[0] ),
    .A2(_1332_),
    .B1(_1342_),
    .B2(\vga.horizontalWholeLineCompare[10] ),
    .C1(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__and4b_1 _2424_ (.A_N(_1044_),
    .B(_1035_),
    .C(_1042_),
    .D(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__and4b_4 _2425_ (.A_N(_1045_),
    .B(_1036_),
    .C(_1043_),
    .D(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__o22a_1 _2426_ (.A1(\vga.verticalWholeLineCompare[7] ),
    .A2(_1320_),
    .B1(_1323_),
    .B2(\vga.verticalWholeLineCompare[4] ),
    .X(_1050_));
 sky130_fd_sc_hd__o221a_1 _2427_ (.A1(\vga.verticalWholeLineCompare[9] ),
    .A2(_1318_),
    .B1(\vga.verticalCounter[5] ),
    .B2(_1294_),
    .C1(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__xnor2_1 _2428_ (.A(\vga.verticalWholeLineCompare[3] ),
    .B(\vga.verticalCounter[3] ),
    .Y(_1052_));
 sky130_fd_sc_hd__o221a_1 _2429_ (.A1(_1292_),
    .A2(\vga.verticalCounter[1] ),
    .B1(_1327_),
    .B2(\vga.verticalWholeLineCompare[0] ),
    .C1(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__xnor2_1 _2430_ (.A(\vga.verticalWholeLineCompare[8] ),
    .B(\vga.verticalCounter[8] ),
    .Y(_1054_));
 sky130_fd_sc_hd__o221a_1 _2431_ (.A1(_1295_),
    .A2(\vga.verticalCounter[6] ),
    .B1(_1326_),
    .B2(\vga.verticalWholeLineCompare[1] ),
    .C1(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__o2bb2a_1 _2432_ (.A1_N(\vga.verticalWholeLineCompare[2] ),
    .A2_N(_1325_),
    .B1(_1322_),
    .B2(\vga.verticalWholeLineCompare[5] ),
    .X(_1056_));
 sky130_fd_sc_hd__o221a_1 _2433_ (.A1(_1296_),
    .A2(\vga.verticalCounter[7] ),
    .B1(_1325_),
    .B2(\vga.verticalWholeLineCompare[2] ),
    .C1(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__o2bb2a_1 _2434_ (.A1_N(\vga.verticalWholeLineCompare[9] ),
    .A2_N(_1318_),
    .B1(_1321_),
    .B2(\vga.verticalWholeLineCompare[6] ),
    .X(_1058_));
 sky130_fd_sc_hd__o221a_1 _2435_ (.A1(_1293_),
    .A2(\vga.verticalCounter[4] ),
    .B1(\vga.verticalCounter[0] ),
    .B2(_1291_),
    .C1(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__and3_1 _2436_ (.A(_1055_),
    .B(_1057_),
    .C(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__and4_4 _2437_ (.A(_1049_),
    .B(_1051_),
    .C(_1053_),
    .D(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__nor2_8 _2438_ (.A(_0283_),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__inv_2 _2439_ (.A(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__xor2_1 _2440_ (.A(\vga.verticalVisibleAreaCompare[0] ),
    .B(\vga.verticalCounter[0] ),
    .X(_1064_));
 sky130_fd_sc_hd__or2_1 _2441_ (.A(\vga.verticalVisibleAreaCompare[9] ),
    .B(\vga.verticalCounter[9] ),
    .X(_1065_));
 sky130_fd_sc_hd__nand2_1 _2442_ (.A(\vga.verticalVisibleAreaCompare[9] ),
    .B(\vga.verticalCounter[9] ),
    .Y(_1066_));
 sky130_fd_sc_hd__a221o_1 _2443_ (.A1(\vga.verticalVisibleAreaCompare[2] ),
    .A2(_1325_),
    .B1(_1065_),
    .B2(_1066_),
    .C1(_0283_),
    .X(_1067_));
 sky130_fd_sc_hd__xor2_1 _2444_ (.A(\vga.verticalVisibleAreaCompare[3] ),
    .B(\vga.verticalCounter[3] ),
    .X(_1068_));
 sky130_fd_sc_hd__a221o_1 _2445_ (.A1(_1303_),
    .A2(\vga.verticalCounter[5] ),
    .B1(_1326_),
    .B2(\vga.verticalVisibleAreaCompare[1] ),
    .C1(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__a22o_1 _2446_ (.A1(\vga.verticalVisibleAreaCompare[6] ),
    .A2(_1321_),
    .B1(_1322_),
    .B2(\vga.verticalVisibleAreaCompare[5] ),
    .X(_1070_));
 sky130_fd_sc_hd__a221o_1 _2447_ (.A1(\vga.verticalVisibleAreaCompare[8] ),
    .A2(_1319_),
    .B1(_1323_),
    .B2(\vga.verticalVisibleAreaCompare[4] ),
    .C1(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__o22a_1 _2448_ (.A1(\vga.verticalVisibleAreaCompare[7] ),
    .A2(_1320_),
    .B1(_1326_),
    .B2(\vga.verticalVisibleAreaCompare[1] ),
    .X(_1072_));
 sky130_fd_sc_hd__o2bb2a_1 _2449_ (.A1_N(\vga.verticalVisibleAreaCompare[7] ),
    .A2_N(_1320_),
    .B1(_1323_),
    .B2(\vga.verticalVisibleAreaCompare[4] ),
    .X(_1073_));
 sky130_fd_sc_hd__o221a_1 _2450_ (.A1(\vga.verticalVisibleAreaCompare[8] ),
    .A2(_1319_),
    .B1(_1321_),
    .B2(\vga.verticalVisibleAreaCompare[6] ),
    .C1(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__o211a_1 _2451_ (.A1(\vga.verticalVisibleAreaCompare[2] ),
    .A2(_1325_),
    .B1(_1072_),
    .C1(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__or3b_1 _2452_ (.A(_1069_),
    .B(_1071_),
    .C_N(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__or4b_4 _2453_ (.A(_1064_),
    .B(_1067_),
    .C(_1076_),
    .D_N(_1049_),
    .X(_1077_));
 sky130_fd_sc_hd__o21a_1 _2454_ (.A1(\vga.inVerticalVisibleArea ),
    .A2(_1063_),
    .B1(_1077_),
    .X(_0144_));
 sky130_fd_sc_hd__and2_1 _2455_ (.A(\vga.verticalCounter[0] ),
    .B(_1049_),
    .X(_1078_));
 sky130_fd_sc_hd__o21ai_1 _2456_ (.A1(\vga.verticalCounter[0] ),
    .A2(_1049_),
    .B1(_1062_),
    .Y(_1079_));
 sky130_fd_sc_hd__nor2_1 _2457_ (.A(_1078_),
    .B(_1079_),
    .Y(_0145_));
 sky130_fd_sc_hd__and3_1 _2458_ (.A(\vga.verticalCounter[1] ),
    .B(\vga.verticalCounter[0] ),
    .C(_1049_),
    .X(_1080_));
 sky130_fd_sc_hd__inv_2 _2459_ (.A(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__o211a_1 _2460_ (.A1(\vga.verticalCounter[1] ),
    .A2(_1078_),
    .B1(_1081_),
    .C1(_1062_),
    .X(_0146_));
 sky130_fd_sc_hd__nor2_2 _2461_ (.A(_1325_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__inv_2 _2462_ (.A(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__o211a_1 _2463_ (.A1(\vga.verticalCounter[2] ),
    .A2(_1080_),
    .B1(_1083_),
    .C1(_1062_),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_1 _2464_ (.A(_1324_),
    .B(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__o21ai_1 _2465_ (.A1(\vga.verticalCounter[3] ),
    .A2(_1082_),
    .B1(_1062_),
    .Y(_1085_));
 sky130_fd_sc_hd__nor2_1 _2466_ (.A(_1084_),
    .B(_1085_),
    .Y(_0148_));
 sky130_fd_sc_hd__or2_1 _2467_ (.A(\vga.verticalCounter[4] ),
    .B(_1084_),
    .X(_1086_));
 sky130_fd_sc_hd__and3_1 _2468_ (.A(\vga.verticalCounter[4] ),
    .B(\vga.verticalCounter[3] ),
    .C(_1082_),
    .X(_1087_));
 sky130_fd_sc_hd__and3b_1 _2469_ (.A_N(_1087_),
    .B(_1062_),
    .C(_1086_),
    .X(_0149_));
 sky130_fd_sc_hd__or2_1 _2470_ (.A(\vga.verticalCounter[5] ),
    .B(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__and2_1 _2471_ (.A(\vga.verticalCounter[5] ),
    .B(_1087_),
    .X(_1089_));
 sky130_fd_sc_hd__and3b_1 _2472_ (.A_N(_1089_),
    .B(_1062_),
    .C(_1088_),
    .X(_0150_));
 sky130_fd_sc_hd__and3_1 _2473_ (.A(\vga.verticalCounter[6] ),
    .B(\vga.verticalCounter[5] ),
    .C(_1087_),
    .X(_1090_));
 sky130_fd_sc_hd__o21ai_1 _2474_ (.A1(\vga.verticalCounter[6] ),
    .A2(_1089_),
    .B1(_1062_),
    .Y(_1091_));
 sky130_fd_sc_hd__nor2_1 _2475_ (.A(_1090_),
    .B(_1091_),
    .Y(_0151_));
 sky130_fd_sc_hd__nand2_1 _2476_ (.A(\vga.verticalCounter[7] ),
    .B(_1090_),
    .Y(_1092_));
 sky130_fd_sc_hd__o211a_1 _2477_ (.A1(\vga.verticalCounter[7] ),
    .A2(_1090_),
    .B1(_1092_),
    .C1(_1062_),
    .X(_0152_));
 sky130_fd_sc_hd__nand2_1 _2478_ (.A(_1319_),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__nor2_1 _2479_ (.A(_1319_),
    .B(_1092_),
    .Y(_1094_));
 sky130_fd_sc_hd__and3b_1 _2480_ (.A_N(_1094_),
    .B(_1062_),
    .C(_1093_),
    .X(_0153_));
 sky130_fd_sc_hd__a21oi_1 _2481_ (.A1(\vga.verticalCounter[9] ),
    .A2(_1094_),
    .B1(_1063_),
    .Y(_1095_));
 sky130_fd_sc_hd__o21a_1 _2482_ (.A1(\vga.verticalCounter[9] ),
    .A2(_1094_),
    .B1(_1095_),
    .X(_0154_));
 sky130_fd_sc_hd__xnor2_1 _2483_ (.A(\vga.verticalSyncPulseCompare[9] ),
    .B(\vga.verticalCounter[9] ),
    .Y(_1096_));
 sky130_fd_sc_hd__xor2_1 _2484_ (.A(\vga.verticalSyncPulseCompare[0] ),
    .B(\vga.verticalCounter[0] ),
    .X(_1097_));
 sky130_fd_sc_hd__xor2_1 _2485_ (.A(\vga.verticalSyncPulseCompare[4] ),
    .B(\vga.verticalCounter[4] ),
    .X(_1098_));
 sky130_fd_sc_hd__a221o_1 _2486_ (.A1(_1300_),
    .A2(\vga.verticalCounter[6] ),
    .B1(\vga.verticalCounter[3] ),
    .B2(_1299_),
    .C1(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__a22o_1 _2487_ (.A1(\vga.verticalSyncPulseCompare[2] ),
    .A2(_1325_),
    .B1(\vga.verticalCounter[1] ),
    .B2(_1297_),
    .X(_1100_));
 sky130_fd_sc_hd__a221o_1 _2488_ (.A1(\vga.verticalSyncPulseCompare[7] ),
    .A2(_1320_),
    .B1(_1322_),
    .B2(\vga.verticalSyncPulseCompare[5] ),
    .C1(_1097_),
    .X(_1101_));
 sky130_fd_sc_hd__a221o_1 _2489_ (.A1(\vga.verticalSyncPulseCompare[6] ),
    .A2(_1321_),
    .B1(_1324_),
    .B2(\vga.verticalSyncPulseCompare[3] ),
    .C1(_1100_),
    .X(_1102_));
 sky130_fd_sc_hd__o22a_1 _2490_ (.A1(\vga.verticalSyncPulseCompare[8] ),
    .A2(_1319_),
    .B1(\vga.verticalCounter[1] ),
    .B2(_1297_),
    .X(_1103_));
 sky130_fd_sc_hd__o2bb2a_1 _2491_ (.A1_N(\vga.verticalSyncPulseCompare[8] ),
    .A2_N(_1319_),
    .B1(_1325_),
    .B2(\vga.verticalSyncPulseCompare[2] ),
    .X(_1104_));
 sky130_fd_sc_hd__o221a_1 _2492_ (.A1(\vga.verticalSyncPulseCompare[7] ),
    .A2(_1320_),
    .B1(_1322_),
    .B2(\vga.verticalSyncPulseCompare[5] ),
    .C1(_1096_),
    .X(_1105_));
 sky130_fd_sc_hd__and4_1 _2493_ (.A(_1049_),
    .B(_1103_),
    .C(_1104_),
    .D(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__or4b_4 _2494_ (.A(_1099_),
    .B(_1101_),
    .C(_1102_),
    .D_N(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__xor2_1 _2495_ (.A(\vga.verticalFrontPorchCompare[6] ),
    .B(\vga.verticalCounter[6] ),
    .X(_1108_));
 sky130_fd_sc_hd__nand2_1 _2496_ (.A(\vga.verticalFrontPorchCompare[7] ),
    .B(\vga.verticalCounter[7] ),
    .Y(_1109_));
 sky130_fd_sc_hd__or2_1 _2497_ (.A(\vga.verticalFrontPorchCompare[7] ),
    .B(\vga.verticalCounter[7] ),
    .X(_1110_));
 sky130_fd_sc_hd__a221o_1 _2498_ (.A1(\vga.verticalFrontPorchCompare[9] ),
    .A2(_1318_),
    .B1(_1109_),
    .B2(_1110_),
    .C1(_0283_),
    .X(_1111_));
 sky130_fd_sc_hd__a22o_1 _2499_ (.A1(\vga.verticalFrontPorchCompare[4] ),
    .A2(_1323_),
    .B1(_1325_),
    .B2(\vga.verticalFrontPorchCompare[2] ),
    .X(_1112_));
 sky130_fd_sc_hd__a221o_1 _2500_ (.A1(\vga.verticalFrontPorchCompare[8] ),
    .A2(_1319_),
    .B1(\vga.verticalCounter[0] ),
    .B2(_1301_),
    .C1(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__a2bb2o_1 _2501_ (.A1_N(\vga.verticalFrontPorchCompare[9] ),
    .A2_N(_1318_),
    .B1(_1322_),
    .B2(\vga.verticalFrontPorchCompare[5] ),
    .X(_1114_));
 sky130_fd_sc_hd__a221o_1 _2502_ (.A1(_1302_),
    .A2(\vga.verticalCounter[2] ),
    .B1(_1326_),
    .B2(\vga.verticalFrontPorchCompare[1] ),
    .C1(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__o2bb2a_1 _2503_ (.A1_N(\vga.verticalFrontPorchCompare[3] ),
    .A2_N(_1324_),
    .B1(_1326_),
    .B2(\vga.verticalFrontPorchCompare[1] ),
    .X(_1116_));
 sky130_fd_sc_hd__o22a_1 _2504_ (.A1(\vga.verticalFrontPorchCompare[3] ),
    .A2(_1324_),
    .B1(\vga.verticalCounter[0] ),
    .B2(_1301_),
    .X(_1117_));
 sky130_fd_sc_hd__o221a_1 _2505_ (.A1(\vga.verticalFrontPorchCompare[8] ),
    .A2(_1319_),
    .B1(_1322_),
    .B2(\vga.verticalFrontPorchCompare[5] ),
    .C1(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__o211a_1 _2506_ (.A1(\vga.verticalFrontPorchCompare[4] ),
    .A2(_1323_),
    .B1(_1116_),
    .C1(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__or3b_1 _2507_ (.A(_1113_),
    .B(_1115_),
    .C_N(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__or4b_2 _2508_ (.A(_1108_),
    .B(_1111_),
    .C(_1120_),
    .D_N(_1049_),
    .X(_1121_));
 sky130_fd_sc_hd__a21boi_2 _2509_ (.A1(_0061_),
    .A2(_1107_),
    .B1_N(_1121_),
    .Y(_0155_));
 sky130_fd_sc_hd__nor2_8 _2510_ (.A(_0283_),
    .B(_1049_),
    .Y(_1122_));
 sky130_fd_sc_hd__clkinv_4 _2511_ (.A(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__o2bb2a_1 _2512_ (.A1_N(net543),
    .A2_N(net529),
    .B1(_1123_),
    .B2(\vga.inHorizontalVisibleArea ),
    .X(_0156_));
 sky130_fd_sc_hd__xnor2_1 _2513_ (.A(\vga.horizontalSyncPulseCompare[2] ),
    .B(\vga.horizontalCounter[2] ),
    .Y(_1124_));
 sky130_fd_sc_hd__xnor2_1 _2514_ (.A(\vga.horizontalSyncPulseCompare[8] ),
    .B(\vga.horizontalCounter[8] ),
    .Y(_1125_));
 sky130_fd_sc_hd__o221a_1 _2515_ (.A1(_1308_),
    .A2(\vga.horizontalCounter[0] ),
    .B1(_1339_),
    .B2(\vga.horizontalSyncPulseCompare[7] ),
    .C1(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__o221a_1 _2516_ (.A1(_1309_),
    .A2(\vga.horizontalCounter[3] ),
    .B1(_1336_),
    .B2(\vga.horizontalSyncPulseCompare[4] ),
    .C1(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__o2bb2a_1 _2517_ (.A1_N(\vga.horizontalSyncPulseCompare[7] ),
    .A2_N(_1339_),
    .B1(_1333_),
    .B2(\vga.horizontalSyncPulseCompare[1] ),
    .X(_1128_));
 sky130_fd_sc_hd__o221a_1 _2518_ (.A1(\vga.horizontalSyncPulseCompare[3] ),
    .A2(_1335_),
    .B1(_1341_),
    .B2(\vga.horizontalSyncPulseCompare[9] ),
    .C1(_1124_),
    .X(_1129_));
 sky130_fd_sc_hd__o2bb2a_1 _2519_ (.A1_N(\vga.horizontalSyncPulseCompare[1] ),
    .A2_N(_1333_),
    .B1(_1342_),
    .B2(\vga.horizontalSyncPulseCompare[10] ),
    .X(_1130_));
 sky130_fd_sc_hd__o221a_1 _2520_ (.A1(\vga.horizontalSyncPulseCompare[5] ),
    .A2(_1337_),
    .B1(_1338_),
    .B2(\vga.horizontalSyncPulseCompare[6] ),
    .C1(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__a22o_1 _2521_ (.A1(\vga.horizontalSyncPulseCompare[4] ),
    .A2(_1336_),
    .B1(_1337_),
    .B2(\vga.horizontalSyncPulseCompare[5] ),
    .X(_1132_));
 sky130_fd_sc_hd__a221oi_1 _2522_ (.A1(\vga.horizontalSyncPulseCompare[9] ),
    .A2(_1341_),
    .B1(_1342_),
    .B2(\vga.horizontalSyncPulseCompare[10] ),
    .C1(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__o221a_1 _2523_ (.A1(\vga.horizontalSyncPulseCompare[0] ),
    .A2(_1332_),
    .B1(\vga.horizontalCounter[6] ),
    .B2(_1310_),
    .C1(_1128_),
    .X(_1134_));
 sky130_fd_sc_hd__and3_1 _2524_ (.A(_1131_),
    .B(_1133_),
    .C(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__xor2_1 _2525_ (.A(\vga.horizontalFrontPorchCompare[1] ),
    .B(\vga.horizontalCounter[1] ),
    .X(_1136_));
 sky130_fd_sc_hd__nor2_1 _2526_ (.A(\vga.horizontalFrontPorchCompare[8] ),
    .B(_1340_),
    .Y(_1137_));
 sky130_fd_sc_hd__o22a_1 _2527_ (.A1(_1312_),
    .A2(\vga.horizontalCounter[2] ),
    .B1(_1335_),
    .B2(\vga.horizontalFrontPorchCompare[3] ),
    .X(_1138_));
 sky130_fd_sc_hd__nor2_1 _2528_ (.A(\vga.horizontalFrontPorchCompare[7] ),
    .B(_1339_),
    .Y(_1139_));
 sky130_fd_sc_hd__nor2_1 _2529_ (.A(\vga.horizontalFrontPorchCompare[0] ),
    .B(_1332_),
    .Y(_1140_));
 sky130_fd_sc_hd__o22a_1 _2530_ (.A1(\vga.horizontalFrontPorchCompare[5] ),
    .A2(_1337_),
    .B1(_1342_),
    .B2(\vga.horizontalFrontPorchCompare[10] ),
    .X(_1141_));
 sky130_fd_sc_hd__o21ai_1 _2531_ (.A1(\vga.horizontalFrontPorchCompare[9] ),
    .A2(_1341_),
    .B1(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__a221o_1 _2532_ (.A1(_1313_),
    .A2(\vga.horizontalCounter[4] ),
    .B1(_1341_),
    .B2(\vga.horizontalFrontPorchCompare[9] ),
    .C1(_1137_),
    .X(_1143_));
 sky130_fd_sc_hd__a221o_1 _2533_ (.A1(\vga.horizontalFrontPorchCompare[4] ),
    .A2(_1336_),
    .B1(\vga.horizontalCounter[6] ),
    .B2(_1314_),
    .C1(_1136_),
    .X(_1144_));
 sky130_fd_sc_hd__a22o_1 _2534_ (.A1(_1312_),
    .A2(\vga.horizontalCounter[2] ),
    .B1(_1337_),
    .B2(\vga.horizontalFrontPorchCompare[5] ),
    .X(_1145_));
 sky130_fd_sc_hd__a221o_1 _2535_ (.A1(\vga.horizontalFrontPorchCompare[7] ),
    .A2(_1339_),
    .B1(_1342_),
    .B2(\vga.horizontalFrontPorchCompare[10] ),
    .C1(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__a221o_1 _2536_ (.A1(\vga.horizontalFrontPorchCompare[3] ),
    .A2(_1335_),
    .B1(_1340_),
    .B2(\vga.horizontalFrontPorchCompare[8] ),
    .C1(_1139_),
    .X(_1147_));
 sky130_fd_sc_hd__a221o_1 _2537_ (.A1(\vga.horizontalFrontPorchCompare[0] ),
    .A2(_1332_),
    .B1(_1338_),
    .B2(\vga.horizontalFrontPorchCompare[6] ),
    .C1(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__or4_1 _2538_ (.A(_1143_),
    .B(_1144_),
    .C(_1146_),
    .D(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__or4b_2 _2539_ (.A(_1140_),
    .B(_1142_),
    .C(_1149_),
    .D_N(_1138_),
    .X(_1150_));
 sky130_fd_sc_hd__a31o_1 _2540_ (.A1(_1127_),
    .A2(_1129_),
    .A3(_1135_),
    .B1(\vga.hsync ),
    .X(_1151_));
 sky130_fd_sc_hd__a21o_1 _2541_ (.A1(_1150_),
    .A2(_1151_),
    .B1(_0283_),
    .X(_0158_));
 sky130_fd_sc_hd__nor2_1 _2542_ (.A(\vga.horizontalCounter[0] ),
    .B(_1123_),
    .Y(_0159_));
 sky130_fd_sc_hd__or2_1 _2543_ (.A(\vga.horizontalCounter[0] ),
    .B(\vga.horizontalCounter[1] ),
    .X(_1152_));
 sky130_fd_sc_hd__nand2_2 _2544_ (.A(\vga.horizontalCounter[0] ),
    .B(\vga.horizontalCounter[1] ),
    .Y(_1153_));
 sky130_fd_sc_hd__and3_1 _2545_ (.A(_1122_),
    .B(_1152_),
    .C(_1153_),
    .X(_0160_));
 sky130_fd_sc_hd__nor2_4 _2546_ (.A(_1334_),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__nand2_1 _2547_ (.A(_1334_),
    .B(_1153_),
    .Y(_1155_));
 sky130_fd_sc_hd__and3b_1 _2548_ (.A_N(_1154_),
    .B(_1155_),
    .C(_1122_),
    .X(_0161_));
 sky130_fd_sc_hd__and2_1 _2549_ (.A(\vga.horizontalCounter[3] ),
    .B(_1154_),
    .X(_1156_));
 sky130_fd_sc_hd__o21ai_1 _2550_ (.A1(\vga.horizontalCounter[3] ),
    .A2(_1154_),
    .B1(_1122_),
    .Y(_1157_));
 sky130_fd_sc_hd__nor2_1 _2551_ (.A(_1156_),
    .B(_1157_),
    .Y(_0162_));
 sky130_fd_sc_hd__and3_2 _2552_ (.A(\vga.horizontalCounter[3] ),
    .B(\vga.horizontalCounter[4] ),
    .C(_1154_),
    .X(_1158_));
 sky130_fd_sc_hd__o21ai_1 _2553_ (.A1(\vga.horizontalCounter[4] ),
    .A2(_1156_),
    .B1(_1122_),
    .Y(_1159_));
 sky130_fd_sc_hd__nor2_1 _2554_ (.A(_1158_),
    .B(_1159_),
    .Y(_0163_));
 sky130_fd_sc_hd__and2_1 _2555_ (.A(\vga.horizontalCounter[5] ),
    .B(_1158_),
    .X(_1160_));
 sky130_fd_sc_hd__o21ai_1 _2556_ (.A1(\vga.horizontalCounter[5] ),
    .A2(_1158_),
    .B1(_1122_),
    .Y(_1161_));
 sky130_fd_sc_hd__nor2_1 _2557_ (.A(_1160_),
    .B(_1161_),
    .Y(_0164_));
 sky130_fd_sc_hd__or2_1 _2558_ (.A(\vga.horizontalCounter[6] ),
    .B(_1160_),
    .X(_1162_));
 sky130_fd_sc_hd__and3_1 _2559_ (.A(\vga.horizontalCounter[5] ),
    .B(\vga.horizontalCounter[6] ),
    .C(_1158_),
    .X(_1163_));
 sky130_fd_sc_hd__and3b_1 _2560_ (.A_N(_1163_),
    .B(_1122_),
    .C(_1162_),
    .X(_0165_));
 sky130_fd_sc_hd__nand2_1 _2561_ (.A(\vga.horizontalCounter[7] ),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__o211a_1 _2562_ (.A1(\vga.horizontalCounter[7] ),
    .A2(_1163_),
    .B1(_1164_),
    .C1(_1122_),
    .X(_0166_));
 sky130_fd_sc_hd__nor2_1 _2563_ (.A(_1340_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__a211oi_1 _2564_ (.A1(_1340_),
    .A2(_1164_),
    .B1(_1165_),
    .C1(_1123_),
    .Y(_0167_));
 sky130_fd_sc_hd__nand2_1 _2565_ (.A(\vga.horizontalCounter[9] ),
    .B(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__o211a_1 _2566_ (.A1(\vga.horizontalCounter[9] ),
    .A2(_1165_),
    .B1(_1166_),
    .C1(_1122_),
    .X(_0168_));
 sky130_fd_sc_hd__nand2_1 _2567_ (.A(_1342_),
    .B(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__o211a_1 _2568_ (.A1(_1342_),
    .A2(_1166_),
    .B1(_1167_),
    .C1(_1122_),
    .X(_0169_));
 sky130_fd_sc_hd__nand3_4 _2569_ (.A(net598),
    .B(net584),
    .C(_0527_),
    .Y(_1168_));
 sky130_fd_sc_hd__and4_4 _2570_ (.A(net583),
    .B(_1355_),
    .C(_0267_),
    .D(_0567_),
    .X(_1169_));
 sky130_fd_sc_hd__mux2_1 _2571_ (.A0(net275),
    .A1(\vga.configuration[12] ),
    .S(_1168_),
    .X(_1170_));
 sky130_fd_sc_hd__and2_1 _2572_ (.A(net604),
    .B(_1170_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(net274),
    .A1(\vga.configuration[11] ),
    .S(_1168_),
    .X(_1171_));
 sky130_fd_sc_hd__and2_1 _2574_ (.A(net603),
    .B(_1171_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _2575_ (.A0(net273),
    .A1(\vga.configuration[10] ),
    .S(_1168_),
    .X(_1172_));
 sky130_fd_sc_hd__and2_1 _2576_ (.A(net605),
    .B(_1172_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2577_ (.A0(net303),
    .A1(\vga.configuration[9] ),
    .S(_1168_),
    .X(_1173_));
 sky130_fd_sc_hd__and2_1 _2578_ (.A(net604),
    .B(_1173_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2579_ (.A0(net302),
    .A1(\vga.configuration[8] ),
    .S(_1168_),
    .X(_1174_));
 sky130_fd_sc_hd__and2_1 _2580_ (.A(net604),
    .B(_1174_),
    .X(_0174_));
 sky130_fd_sc_hd__and2_1 _2581_ (.A(net601),
    .B(_1169_),
    .X(_1175_));
 sky130_fd_sc_hd__nand2_4 _2582_ (.A(net601),
    .B(_1169_),
    .Y(_1176_));
 sky130_fd_sc_hd__and3_1 _2583_ (.A(net602),
    .B(net301),
    .C(_1169_),
    .X(_1177_));
 sky130_fd_sc_hd__a211o_1 _2584_ (.A1(\vga.configuration[7] ),
    .A2(_1176_),
    .B1(_1177_),
    .C1(net613),
    .X(_0175_));
 sky130_fd_sc_hd__or2_1 _2585_ (.A(\vga.configuration[6] ),
    .B(_1175_),
    .X(_1178_));
 sky130_fd_sc_hd__o211a_1 _2586_ (.A1(net300),
    .A2(_1176_),
    .B1(_1178_),
    .C1(net606),
    .X(_0176_));
 sky130_fd_sc_hd__and3_1 _2587_ (.A(net602),
    .B(net299),
    .C(_1169_),
    .X(_1179_));
 sky130_fd_sc_hd__a211o_1 _2588_ (.A1(\vga.configuration[5] ),
    .A2(_1176_),
    .B1(_1179_),
    .C1(net613),
    .X(_0177_));
 sky130_fd_sc_hd__or2_1 _2589_ (.A(\vga.configuration[4] ),
    .B(_1175_),
    .X(_1180_));
 sky130_fd_sc_hd__o211a_1 _2590_ (.A1(net298),
    .A2(_1176_),
    .B1(_1180_),
    .C1(net606),
    .X(_0178_));
 sky130_fd_sc_hd__and3_1 _2591_ (.A(net601),
    .B(net297),
    .C(_1169_),
    .X(_1181_));
 sky130_fd_sc_hd__a211o_1 _2592_ (.A1(\vga.configuration[3] ),
    .A2(_1176_),
    .B1(_1181_),
    .C1(net613),
    .X(_0179_));
 sky130_fd_sc_hd__or2_1 _2593_ (.A(\vga.configuration[2] ),
    .B(_1175_),
    .X(_1182_));
 sky130_fd_sc_hd__o211a_1 _2594_ (.A1(net294),
    .A2(_1176_),
    .B1(_1182_),
    .C1(net605),
    .X(_0180_));
 sky130_fd_sc_hd__and3_1 _2595_ (.A(net601),
    .B(net283),
    .C(_1169_),
    .X(_1183_));
 sky130_fd_sc_hd__a211o_1 _2596_ (.A1(\vga.configuration[1] ),
    .A2(_1176_),
    .B1(_1183_),
    .C1(net613),
    .X(_0181_));
 sky130_fd_sc_hd__or2_1 _2597_ (.A(\vga.configuration[0] ),
    .B(_1175_),
    .X(_1184_));
 sky130_fd_sc_hd__o211a_1 _2598_ (.A1(net272),
    .A2(_1176_),
    .B1(_1184_),
    .C1(net606),
    .X(_0182_));
 sky130_fd_sc_hd__and3_2 _2599_ (.A(net598),
    .B(net584),
    .C(_0536_),
    .X(_1185_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(\vga.horizontalVisibleAreaCompare[10] ),
    .A1(net273),
    .S(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__and2_1 _2601_ (.A(net605),
    .B(_1186_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(_1317_),
    .A1(_1344_),
    .S(_1185_),
    .X(_1187_));
 sky130_fd_sc_hd__nand2_1 _2603_ (.A(net605),
    .B(_1187_),
    .Y(_0184_));
 sky130_fd_sc_hd__mux2_1 _2604_ (.A0(_1316_),
    .A1(_1343_),
    .S(_1185_),
    .X(_1188_));
 sky130_fd_sc_hd__nand2_1 _2605_ (.A(net605),
    .B(_1188_),
    .Y(_0185_));
 sky130_fd_sc_hd__and3_4 _2606_ (.A(net602),
    .B(net584),
    .C(_0536_),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(\vga.horizontalVisibleAreaCompare[7] ),
    .A1(net301),
    .S(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__and2_1 _2608_ (.A(net603),
    .B(_1190_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(\vga.horizontalVisibleAreaCompare[6] ),
    .A1(net300),
    .S(_1189_),
    .X(_1191_));
 sky130_fd_sc_hd__and2_1 _2610_ (.A(net603),
    .B(_1191_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(\vga.horizontalVisibleAreaCompare[5] ),
    .A1(net299),
    .S(_1189_),
    .X(_1192_));
 sky130_fd_sc_hd__and2_1 _2612_ (.A(net603),
    .B(_1192_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(\vga.horizontalVisibleAreaCompare[4] ),
    .A1(net298),
    .S(_1189_),
    .X(_1193_));
 sky130_fd_sc_hd__or2_1 _2614_ (.A(net611),
    .B(_1193_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(\vga.horizontalVisibleAreaCompare[3] ),
    .A1(net297),
    .S(_1189_),
    .X(_1194_));
 sky130_fd_sc_hd__or2_1 _2616_ (.A(net610),
    .B(_1194_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(\vga.horizontalVisibleAreaCompare[2] ),
    .A1(net294),
    .S(_1189_),
    .X(_1195_));
 sky130_fd_sc_hd__or2_1 _2618_ (.A(net610),
    .B(_1195_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _2619_ (.A0(\vga.horizontalVisibleAreaCompare[1] ),
    .A1(net283),
    .S(_1189_),
    .X(_1196_));
 sky130_fd_sc_hd__or2_1 _2620_ (.A(net610),
    .B(_1196_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2621_ (.A0(\vga.horizontalVisibleAreaCompare[0] ),
    .A1(net272),
    .S(_1189_),
    .X(_1197_));
 sky130_fd_sc_hd__or2_1 _2622_ (.A(net610),
    .B(_1197_),
    .X(_0193_));
 sky130_fd_sc_hd__and3_2 _2623_ (.A(net598),
    .B(net584),
    .C(_0542_),
    .X(_1198_));
 sky130_fd_sc_hd__mux2_1 _2624_ (.A0(\vga.horizontalFrontPorchCompare[10] ),
    .A1(net273),
    .S(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__and2_1 _2625_ (.A(net603),
    .B(_1199_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2626_ (.A0(\vga.horizontalFrontPorchCompare[9] ),
    .A1(net303),
    .S(_1198_),
    .X(_1200_));
 sky130_fd_sc_hd__or2_1 _2627_ (.A(net612),
    .B(_1200_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _2628_ (.A0(\vga.horizontalFrontPorchCompare[8] ),
    .A1(net302),
    .S(_1198_),
    .X(_1201_));
 sky130_fd_sc_hd__or2_1 _2629_ (.A(net613),
    .B(_1201_),
    .X(_0196_));
 sky130_fd_sc_hd__and3_4 _2630_ (.A(net602),
    .B(net584),
    .C(_0542_),
    .X(_1202_));
 sky130_fd_sc_hd__mux2_1 _2631_ (.A0(\vga.horizontalFrontPorchCompare[7] ),
    .A1(net301),
    .S(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__and2_1 _2632_ (.A(net603),
    .B(_1203_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _2633_ (.A0(\vga.horizontalFrontPorchCompare[6] ),
    .A1(net300),
    .S(_1202_),
    .X(_1204_));
 sky130_fd_sc_hd__or2_1 _2634_ (.A(net611),
    .B(_1204_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2635_ (.A0(\vga.horizontalFrontPorchCompare[5] ),
    .A1(net299),
    .S(_1202_),
    .X(_1205_));
 sky130_fd_sc_hd__and2_1 _2636_ (.A(net603),
    .B(_1205_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _2637_ (.A0(\vga.horizontalFrontPorchCompare[4] ),
    .A1(net298),
    .S(_1202_),
    .X(_1206_));
 sky130_fd_sc_hd__and2_1 _2638_ (.A(net604),
    .B(_1206_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2639_ (.A0(\vga.horizontalFrontPorchCompare[3] ),
    .A1(net297),
    .S(_1202_),
    .X(_1207_));
 sky130_fd_sc_hd__and2_1 _2640_ (.A(net603),
    .B(_1207_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2641_ (.A0(\vga.horizontalFrontPorchCompare[2] ),
    .A1(net294),
    .S(_1202_),
    .X(_1208_));
 sky130_fd_sc_hd__or2_1 _2642_ (.A(net611),
    .B(_1208_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2643_ (.A0(\vga.horizontalFrontPorchCompare[1] ),
    .A1(net283),
    .S(_1202_),
    .X(_1209_));
 sky130_fd_sc_hd__or2_1 _2644_ (.A(net610),
    .B(_1209_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(\vga.horizontalFrontPorchCompare[0] ),
    .A1(net272),
    .S(_1202_),
    .X(_1210_));
 sky130_fd_sc_hd__or2_1 _2646_ (.A(net611),
    .B(_1210_),
    .X(_0204_));
 sky130_fd_sc_hd__and3_2 _2647_ (.A(net597),
    .B(net583),
    .C(_0546_),
    .X(_1211_));
 sky130_fd_sc_hd__mux2_1 _2648_ (.A0(\vga.horizontalSyncPulseCompare[10] ),
    .A1(net273),
    .S(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__and2_1 _2649_ (.A(net605),
    .B(_1212_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2650_ (.A0(_1311_),
    .A1(_1344_),
    .S(_1211_),
    .X(_1213_));
 sky130_fd_sc_hd__nand2_1 _2651_ (.A(net605),
    .B(_1213_),
    .Y(_0206_));
 sky130_fd_sc_hd__mux2_1 _2652_ (.A0(\vga.horizontalSyncPulseCompare[8] ),
    .A1(net302),
    .S(_1211_),
    .X(_1214_));
 sky130_fd_sc_hd__or2_1 _2653_ (.A(net613),
    .B(_1214_),
    .X(_0207_));
 sky130_fd_sc_hd__and3_4 _2654_ (.A(net601),
    .B(net583),
    .C(_0546_),
    .X(_1215_));
 sky130_fd_sc_hd__mux2_1 _2655_ (.A0(\vga.horizontalSyncPulseCompare[7] ),
    .A1(net301),
    .S(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__or2_1 _2656_ (.A(net614),
    .B(_1216_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _2657_ (.A0(\vga.horizontalSyncPulseCompare[6] ),
    .A1(net300),
    .S(_1215_),
    .X(_1217_));
 sky130_fd_sc_hd__or2_1 _2658_ (.A(net614),
    .B(_1217_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(\vga.horizontalSyncPulseCompare[5] ),
    .A1(net299),
    .S(_1215_),
    .X(_1218_));
 sky130_fd_sc_hd__and2_1 _2660_ (.A(net608),
    .B(_1218_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(\vga.horizontalSyncPulseCompare[4] ),
    .A1(net298),
    .S(_1215_),
    .X(_1219_));
 sky130_fd_sc_hd__and2_1 _2662_ (.A(net605),
    .B(_1219_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(\vga.horizontalSyncPulseCompare[3] ),
    .A1(net297),
    .S(_1215_),
    .X(_1220_));
 sky130_fd_sc_hd__and2_1 _2664_ (.A(net605),
    .B(_1220_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(\vga.horizontalSyncPulseCompare[2] ),
    .A1(net294),
    .S(_1215_),
    .X(_1221_));
 sky130_fd_sc_hd__or2_1 _2666_ (.A(net613),
    .B(_1221_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _2667_ (.A0(\vga.horizontalSyncPulseCompare[1] ),
    .A1(net283),
    .S(_1215_),
    .X(_1222_));
 sky130_fd_sc_hd__or2_1 _2668_ (.A(net613),
    .B(_1222_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2669_ (.A0(\vga.horizontalSyncPulseCompare[0] ),
    .A1(net272),
    .S(_1215_),
    .X(_1223_));
 sky130_fd_sc_hd__or2_1 _2670_ (.A(net618),
    .B(_1223_),
    .X(_0215_));
 sky130_fd_sc_hd__and3_4 _2671_ (.A(net583),
    .B(_0539_),
    .C(_0571_),
    .X(_1224_));
 sky130_fd_sc_hd__and2_2 _2672_ (.A(net596),
    .B(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__and2b_1 _2673_ (.A_N(_1225_),
    .B(\vga.horizontalWholeLineCompare[10] ),
    .X(_1226_));
 sky130_fd_sc_hd__a211o_1 _2674_ (.A1(net273),
    .A2(_1225_),
    .B1(_1226_),
    .C1(net614),
    .X(_0216_));
 sky130_fd_sc_hd__a21oi_1 _2675_ (.A1(_1344_),
    .A2(_1225_),
    .B1(net614),
    .Y(_1227_));
 sky130_fd_sc_hd__o21a_1 _2676_ (.A1(\vga.horizontalWholeLineCompare[9] ),
    .A2(_1225_),
    .B1(_1227_),
    .X(_0217_));
 sky130_fd_sc_hd__a21oi_1 _2677_ (.A1(_1343_),
    .A2(_1225_),
    .B1(net614),
    .Y(_1228_));
 sky130_fd_sc_hd__o21a_1 _2678_ (.A1(\vga.horizontalWholeLineCompare[8] ),
    .A2(_1225_),
    .B1(_1228_),
    .X(_0218_));
 sky130_fd_sc_hd__nand2_1 _2679_ (.A(net599),
    .B(_1224_),
    .Y(_1229_));
 sky130_fd_sc_hd__nor2_1 _2680_ (.A(net301),
    .B(net512),
    .Y(_1230_));
 sky130_fd_sc_hd__a211oi_1 _2681_ (.A1(_1307_),
    .A2(net512),
    .B1(_1230_),
    .C1(net614),
    .Y(_0219_));
 sky130_fd_sc_hd__nand2_1 _2682_ (.A(_1306_),
    .B(net512),
    .Y(_1231_));
 sky130_fd_sc_hd__o211a_1 _2683_ (.A1(net300),
    .A2(net512),
    .B1(_1231_),
    .C1(net608),
    .X(_0220_));
 sky130_fd_sc_hd__nand2_1 _2684_ (.A(_1305_),
    .B(net512),
    .Y(_1232_));
 sky130_fd_sc_hd__o211a_1 _2685_ (.A1(net299),
    .A2(net512),
    .B1(_1232_),
    .C1(net608),
    .X(_0221_));
 sky130_fd_sc_hd__and3_1 _2686_ (.A(net599),
    .B(net298),
    .C(_1224_),
    .X(_1233_));
 sky130_fd_sc_hd__a211o_1 _2687_ (.A1(\vga.horizontalWholeLineCompare[4] ),
    .A2(net512),
    .B1(_1233_),
    .C1(net616),
    .X(_0222_));
 sky130_fd_sc_hd__and3_1 _2688_ (.A(net599),
    .B(net297),
    .C(_1224_),
    .X(_1234_));
 sky130_fd_sc_hd__a211o_1 _2689_ (.A1(\vga.horizontalWholeLineCompare[3] ),
    .A2(net512),
    .B1(_1234_),
    .C1(net616),
    .X(_0223_));
 sky130_fd_sc_hd__and3_1 _2690_ (.A(net599),
    .B(net294),
    .C(_1224_),
    .X(_1235_));
 sky130_fd_sc_hd__a211o_1 _2691_ (.A1(\vga.horizontalWholeLineCompare[2] ),
    .A2(net512),
    .B1(_1235_),
    .C1(net614),
    .X(_0224_));
 sky130_fd_sc_hd__and3_1 _2692_ (.A(net599),
    .B(net283),
    .C(_1224_),
    .X(_1236_));
 sky130_fd_sc_hd__a211o_1 _2693_ (.A1(\vga.horizontalWholeLineCompare[1] ),
    .A2(net512),
    .B1(_1236_),
    .C1(net614),
    .X(_0225_));
 sky130_fd_sc_hd__and3_1 _2694_ (.A(net599),
    .B(net272),
    .C(_1224_),
    .X(_1237_));
 sky130_fd_sc_hd__a211o_1 _2695_ (.A1(\vga.horizontalWholeLineCompare[0] ),
    .A2(_1229_),
    .B1(_1237_),
    .C1(net616),
    .X(_0226_));
 sky130_fd_sc_hd__nor2_4 _2696_ (.A(_1352_),
    .B(_0577_),
    .Y(_1238_));
 sky130_fd_sc_hd__nand2_1 _2697_ (.A(net596),
    .B(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__mux2_1 _2698_ (.A0(net303),
    .A1(\vga.verticalVisibleAreaCompare[9] ),
    .S(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__or2_1 _2699_ (.A(net615),
    .B(_1240_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _2700_ (.A0(_1343_),
    .A1(_1304_),
    .S(_1239_),
    .X(_1241_));
 sky130_fd_sc_hd__nor2_1 _2701_ (.A(net614),
    .B(_1241_),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_8 _2702_ (.A(net599),
    .B(_1238_),
    .Y(_1242_));
 sky130_fd_sc_hd__mux2_1 _2703_ (.A0(net301),
    .A1(\vga.verticalVisibleAreaCompare[7] ),
    .S(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__and2_1 _2704_ (.A(net607),
    .B(_1243_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _2705_ (.A0(net300),
    .A1(\vga.verticalVisibleAreaCompare[6] ),
    .S(_1242_),
    .X(_1244_));
 sky130_fd_sc_hd__or2_1 _2706_ (.A(net616),
    .B(_1244_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _2707_ (.A0(net299),
    .A1(\vga.verticalVisibleAreaCompare[5] ),
    .S(_1242_),
    .X(_1245_));
 sky130_fd_sc_hd__and2_1 _2708_ (.A(net607),
    .B(_1245_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(net298),
    .A1(\vga.verticalVisibleAreaCompare[4] ),
    .S(_1242_),
    .X(_1246_));
 sky130_fd_sc_hd__or2_1 _2710_ (.A(net616),
    .B(_1246_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _2711_ (.A0(net297),
    .A1(\vga.verticalVisibleAreaCompare[3] ),
    .S(_1242_),
    .X(_1247_));
 sky130_fd_sc_hd__and2_1 _2712_ (.A(net607),
    .B(_1247_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2713_ (.A0(net294),
    .A1(\vga.verticalVisibleAreaCompare[2] ),
    .S(_1242_),
    .X(_1248_));
 sky130_fd_sc_hd__or2_1 _2714_ (.A(net616),
    .B(_1248_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2715_ (.A0(net283),
    .A1(\vga.verticalVisibleAreaCompare[1] ),
    .S(_1242_),
    .X(_1249_));
 sky130_fd_sc_hd__or2_1 _2716_ (.A(net616),
    .B(_1249_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _2717_ (.A0(net272),
    .A1(\vga.verticalVisibleAreaCompare[0] ),
    .S(_1242_),
    .X(_1250_));
 sky130_fd_sc_hd__or2_1 _2718_ (.A(net616),
    .B(_1250_),
    .X(_0236_));
 sky130_fd_sc_hd__nor2_8 _2719_ (.A(_1352_),
    .B(_0556_),
    .Y(_1251_));
 sky130_fd_sc_hd__nand2_1 _2720_ (.A(net597),
    .B(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__a31o_1 _2721_ (.A1(net597),
    .A2(net303),
    .A3(_1251_),
    .B1(net615),
    .X(_1253_));
 sky130_fd_sc_hd__a21o_1 _2722_ (.A1(\vga.verticalFrontPorchCompare[9] ),
    .A2(_1252_),
    .B1(_1253_),
    .X(_0237_));
 sky130_fd_sc_hd__a21o_1 _2723_ (.A1(net597),
    .A2(_1251_),
    .B1(\vga.verticalFrontPorchCompare[8] ),
    .X(_1254_));
 sky130_fd_sc_hd__o211a_1 _2724_ (.A1(net302),
    .A2(_1252_),
    .B1(_1254_),
    .C1(net608),
    .X(_0238_));
 sky130_fd_sc_hd__nand2_8 _2725_ (.A(net599),
    .B(_1251_),
    .Y(_1255_));
 sky130_fd_sc_hd__mux2_1 _2726_ (.A0(net301),
    .A1(\vga.verticalFrontPorchCompare[7] ),
    .S(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__and2_1 _2727_ (.A(net607),
    .B(_1256_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _2728_ (.A0(net300),
    .A1(\vga.verticalFrontPorchCompare[6] ),
    .S(_1255_),
    .X(_1257_));
 sky130_fd_sc_hd__or2_1 _2729_ (.A(net616),
    .B(_1257_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2730_ (.A0(net299),
    .A1(\vga.verticalFrontPorchCompare[5] ),
    .S(_1255_),
    .X(_1258_));
 sky130_fd_sc_hd__and2_1 _2731_ (.A(net607),
    .B(_1258_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(net298),
    .A1(\vga.verticalFrontPorchCompare[4] ),
    .S(_1255_),
    .X(_1259_));
 sky130_fd_sc_hd__or2_1 _2733_ (.A(net617),
    .B(_1259_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(net297),
    .A1(\vga.verticalFrontPorchCompare[3] ),
    .S(_1255_),
    .X(_1260_));
 sky130_fd_sc_hd__or2_1 _2735_ (.A(net617),
    .B(_1260_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _2736_ (.A0(net294),
    .A1(\vga.verticalFrontPorchCompare[2] ),
    .S(_1255_),
    .X(_1261_));
 sky130_fd_sc_hd__and2_1 _2737_ (.A(net607),
    .B(_1261_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(net283),
    .A1(\vga.verticalFrontPorchCompare[1] ),
    .S(_1255_),
    .X(_1262_));
 sky130_fd_sc_hd__and2_1 _2739_ (.A(net607),
    .B(_1262_),
    .X(_0245_));
 sky130_fd_sc_hd__a21oi_1 _2740_ (.A1(_1301_),
    .A2(_1255_),
    .B1(net616),
    .Y(_1263_));
 sky130_fd_sc_hd__o21a_1 _2741_ (.A1(net272),
    .A2(_1255_),
    .B1(_1263_),
    .X(_0246_));
 sky130_fd_sc_hd__and3_1 _2742_ (.A(net597),
    .B(net583),
    .C(_0570_),
    .X(_1264_));
 sky130_fd_sc_hd__and2b_1 _2743_ (.A_N(_1264_),
    .B(\vga.verticalSyncPulseCompare[9] ),
    .X(_1265_));
 sky130_fd_sc_hd__a211o_1 _2744_ (.A1(net303),
    .A2(_1264_),
    .B1(_1265_),
    .C1(net615),
    .X(_0247_));
 sky130_fd_sc_hd__a21oi_1 _2745_ (.A1(_1343_),
    .A2(_1264_),
    .B1(net615),
    .Y(_1266_));
 sky130_fd_sc_hd__o21a_1 _2746_ (.A1(\vga.verticalSyncPulseCompare[8] ),
    .A2(_1264_),
    .B1(_1266_),
    .X(_0248_));
 sky130_fd_sc_hd__and3_4 _2747_ (.A(net600),
    .B(net583),
    .C(_0570_),
    .X(_1267_));
 sky130_fd_sc_hd__nand3_4 _2748_ (.A(net600),
    .B(net583),
    .C(_0570_),
    .Y(_1268_));
 sky130_fd_sc_hd__or2_1 _2749_ (.A(\vga.verticalSyncPulseCompare[7] ),
    .B(_1267_),
    .X(_1269_));
 sky130_fd_sc_hd__o211a_1 _2750_ (.A1(net301),
    .A2(_1268_),
    .B1(_1269_),
    .C1(net609),
    .X(_0249_));
 sky130_fd_sc_hd__nor2_1 _2751_ (.A(_1300_),
    .B(_1267_),
    .Y(_1270_));
 sky130_fd_sc_hd__a211o_1 _2752_ (.A1(net300),
    .A2(_1267_),
    .B1(_1270_),
    .C1(net617),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _2753_ (.A(\vga.verticalSyncPulseCompare[5] ),
    .B(_1267_),
    .X(_1271_));
 sky130_fd_sc_hd__o211a_1 _2754_ (.A1(net299),
    .A2(_1268_),
    .B1(_1271_),
    .C1(net607),
    .X(_0251_));
 sky130_fd_sc_hd__a21o_1 _2755_ (.A1(\vga.verticalSyncPulseCompare[4] ),
    .A2(_1268_),
    .B1(net617),
    .X(_1272_));
 sky130_fd_sc_hd__a21o_1 _2756_ (.A1(net298),
    .A2(_1267_),
    .B1(_1272_),
    .X(_0252_));
 sky130_fd_sc_hd__nor2_1 _2757_ (.A(_1299_),
    .B(_1267_),
    .Y(_1273_));
 sky130_fd_sc_hd__a211o_1 _2758_ (.A1(net297),
    .A2(_1267_),
    .B1(_1273_),
    .C1(net617),
    .X(_0253_));
 sky130_fd_sc_hd__nor2_1 _2759_ (.A(_1298_),
    .B(_1267_),
    .Y(_1274_));
 sky130_fd_sc_hd__a211o_1 _2760_ (.A1(net294),
    .A2(_1267_),
    .B1(_1274_),
    .C1(net617),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_1 _2761_ (.A(_1297_),
    .B(_1268_),
    .Y(_1275_));
 sky130_fd_sc_hd__o211a_1 _2762_ (.A1(net283),
    .A2(_1268_),
    .B1(_1275_),
    .C1(net607),
    .X(_0255_));
 sky130_fd_sc_hd__or2_1 _2763_ (.A(\vga.verticalSyncPulseCompare[0] ),
    .B(_1267_),
    .X(_1276_));
 sky130_fd_sc_hd__o211a_1 _2764_ (.A1(net272),
    .A2(_1268_),
    .B1(_1276_),
    .C1(net607),
    .X(_0256_));
 sky130_fd_sc_hd__and3_2 _2765_ (.A(net583),
    .B(_0569_),
    .C(_0571_),
    .X(_1277_));
 sky130_fd_sc_hd__nand2_1 _2766_ (.A(net596),
    .B(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__nor2_1 _2767_ (.A(_1344_),
    .B(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__a211o_1 _2768_ (.A1(\vga.verticalWholeLineCompare[9] ),
    .A2(_1278_),
    .B1(_1279_),
    .C1(net615),
    .X(_0257_));
 sky130_fd_sc_hd__a21o_1 _2769_ (.A1(net596),
    .A2(_1277_),
    .B1(\vga.verticalWholeLineCompare[8] ),
    .X(_1280_));
 sky130_fd_sc_hd__o211a_1 _2770_ (.A1(net302),
    .A2(_1278_),
    .B1(_1280_),
    .C1(net608),
    .X(_0258_));
 sky130_fd_sc_hd__and2_2 _2771_ (.A(net600),
    .B(_1277_),
    .X(_1281_));
 sky130_fd_sc_hd__nand2_2 _2772_ (.A(net600),
    .B(_1277_),
    .Y(_1282_));
 sky130_fd_sc_hd__nand2_1 _2773_ (.A(_1296_),
    .B(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__o211a_1 _2774_ (.A1(net301),
    .A2(_1282_),
    .B1(_1283_),
    .C1(net608),
    .X(_0259_));
 sky130_fd_sc_hd__nor2_1 _2775_ (.A(_1295_),
    .B(net511),
    .Y(_1284_));
 sky130_fd_sc_hd__a211o_1 _2776_ (.A1(net300),
    .A2(net511),
    .B1(_1284_),
    .C1(net617),
    .X(_0260_));
 sky130_fd_sc_hd__nor2_1 _2777_ (.A(_1294_),
    .B(net511),
    .Y(_1285_));
 sky130_fd_sc_hd__a211o_1 _2778_ (.A1(net299),
    .A2(_1281_),
    .B1(_1285_),
    .C1(net617),
    .X(_0261_));
 sky130_fd_sc_hd__nor2_1 _2779_ (.A(_1293_),
    .B(net511),
    .Y(_1286_));
 sky130_fd_sc_hd__a211o_1 _2780_ (.A1(net298),
    .A2(net511),
    .B1(_1286_),
    .C1(net617),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _2781_ (.A(\vga.verticalWholeLineCompare[3] ),
    .B(net511),
    .X(_1287_));
 sky130_fd_sc_hd__o211a_1 _2782_ (.A1(net297),
    .A2(_1282_),
    .B1(_1287_),
    .C1(net608),
    .X(_0263_));
 sky130_fd_sc_hd__or2_1 _2783_ (.A(\vga.verticalWholeLineCompare[2] ),
    .B(net511),
    .X(_1288_));
 sky130_fd_sc_hd__o211a_1 _2784_ (.A1(net294),
    .A2(_1282_),
    .B1(_1288_),
    .C1(net608),
    .X(_0264_));
 sky130_fd_sc_hd__nor2_1 _2785_ (.A(_1292_),
    .B(net511),
    .Y(_1289_));
 sky130_fd_sc_hd__a211o_1 _2786_ (.A1(net283),
    .A2(_1281_),
    .B1(_1289_),
    .C1(net615),
    .X(_0265_));
 sky130_fd_sc_hd__nor2_1 _2787_ (.A(_1291_),
    .B(net511),
    .Y(_1290_));
 sky130_fd_sc_hd__a211o_1 _2788_ (.A1(net272),
    .A2(net511),
    .B1(_1290_),
    .C1(net615),
    .X(_0266_));
 sky130_fd_sc_hd__dfxtp_1 _2789_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_0000_),
    .Q(net444));
 sky130_fd_sc_hd__dfxtp_1 _2790_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_0001_),
    .Q(net455));
 sky130_fd_sc_hd__dfxtp_1 _2791_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_0002_),
    .Q(net466));
 sky130_fd_sc_hd__dfxtp_1 _2792_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_0003_),
    .Q(net469));
 sky130_fd_sc_hd__dfxtp_1 _2793_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_0004_),
    .Q(net470));
 sky130_fd_sc_hd__dfxtp_1 _2794_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_0005_),
    .Q(net471));
 sky130_fd_sc_hd__dfxtp_1 _2795_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_0006_),
    .Q(net472));
 sky130_fd_sc_hd__dfxtp_1 _2796_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0007_),
    .Q(net473));
 sky130_fd_sc_hd__dfxtp_1 _2797_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_0008_),
    .Q(net474));
 sky130_fd_sc_hd__dfxtp_1 _2798_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_0009_),
    .Q(net475));
 sky130_fd_sc_hd__dfxtp_1 _2799_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0010_),
    .Q(net445));
 sky130_fd_sc_hd__dfxtp_2 _2800_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_0011_),
    .Q(net446));
 sky130_fd_sc_hd__dfxtp_1 _2801_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_0012_),
    .Q(net447));
 sky130_fd_sc_hd__dfxtp_1 _2802_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0013_),
    .Q(net448));
 sky130_fd_sc_hd__dfxtp_1 _2803_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0014_),
    .Q(net449));
 sky130_fd_sc_hd__dfxtp_1 _2804_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0015_),
    .Q(net450));
 sky130_fd_sc_hd__dfxtp_1 _2805_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0016_),
    .Q(net451));
 sky130_fd_sc_hd__dfxtp_1 _2806_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0017_),
    .Q(net452));
 sky130_fd_sc_hd__dfxtp_1 _2807_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0018_),
    .Q(net453));
 sky130_fd_sc_hd__dfxtp_4 _2808_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0019_),
    .Q(net454));
 sky130_fd_sc_hd__dfxtp_4 _2809_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0020_),
    .Q(net456));
 sky130_fd_sc_hd__dfxtp_2 _2810_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0021_),
    .Q(net457));
 sky130_fd_sc_hd__dfxtp_1 _2811_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0022_),
    .Q(net458));
 sky130_fd_sc_hd__dfxtp_4 _2812_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0023_),
    .Q(net459));
 sky130_fd_sc_hd__dfxtp_4 _2813_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0024_),
    .Q(net460));
 sky130_fd_sc_hd__dfxtp_2 _2814_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_0025_),
    .Q(net461));
 sky130_fd_sc_hd__dfxtp_2 _2815_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0026_),
    .Q(net462));
 sky130_fd_sc_hd__dfxtp_2 _2816_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0027_),
    .Q(net463));
 sky130_fd_sc_hd__dfxtp_2 _2817_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_0028_),
    .Q(net464));
 sky130_fd_sc_hd__dfxtp_2 _2818_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0029_),
    .Q(net465));
 sky130_fd_sc_hd__dfxtp_2 _2819_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0030_),
    .Q(net467));
 sky130_fd_sc_hd__dfxtp_2 _2820_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0031_),
    .Q(net468));
 sky130_fd_sc_hd__dfxtp_1 _2821_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_0032_),
    .Q(net443));
 sky130_fd_sc_hd__dfxtp_1 _2822_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_0033_),
    .Q(net476));
 sky130_fd_sc_hd__dfxtp_4 _2823_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0034_),
    .Q(\wbPeripheralBusInterface.currentAddress[2] ));
 sky130_fd_sc_hd__dfxtp_4 _2824_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0035_),
    .Q(\wbPeripheralBusInterface.currentAddress[3] ));
 sky130_fd_sc_hd__dfxtp_4 _2825_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_0036_),
    .Q(\wbPeripheralBusInterface.currentAddress[4] ));
 sky130_fd_sc_hd__dfxtp_4 _2826_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0037_),
    .Q(\wbPeripheralBusInterface.currentAddress[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2827_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0038_),
    .Q(\wbPeripheralBusInterface.currentAddress[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2828_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0039_),
    .Q(\wbPeripheralBusInterface.currentAddress[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2829_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0040_),
    .Q(\wbPeripheralBusInterface.currentAddress[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2830_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0041_),
    .Q(\wbPeripheralBusInterface.currentAddress[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2831_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0042_),
    .Q(\wbPeripheralBusInterface.currentAddress[10] ));
 sky130_fd_sc_hd__dfxtp_4 _2832_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0043_),
    .Q(\wbPeripheralBusInterface.currentAddress[11] ));
 sky130_fd_sc_hd__dfxtp_4 _2833_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0044_),
    .Q(\wbPeripheralBusInterface.currentAddress[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2834_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0045_),
    .Q(\wbPeripheralBusInterface.currentAddress[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2835_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0046_),
    .Q(\wbPeripheralBusInterface.currentAddress[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2836_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0047_),
    .Q(\wbPeripheralBusInterface.currentAddress[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2837_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0048_),
    .Q(\wbPeripheralBusInterface.currentAddress[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2838_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0049_),
    .Q(\wbPeripheralBusInterface.currentAddress[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2839_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0050_),
    .Q(\wbPeripheralBusInterface.currentAddress[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2840_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0051_),
    .Q(\wbPeripheralBusInterface.currentAddress[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2841_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0052_),
    .Q(\wbPeripheralBusInterface.currentAddress[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2842_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0053_),
    .Q(\wbPeripheralBusInterface.currentAddress[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2843_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0054_),
    .Q(\wbPeripheralBusInterface.currentAddress[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2844_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0055_),
    .Q(\wbPeripheralBusInterface.currentAddress[23] ));
 sky130_fd_sc_hd__dfxtp_4 _2845_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_0056_),
    .Q(\videoMemory.wbReadReady ));
 sky130_fd_sc_hd__dfxtp_4 _2846_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0057_),
    .Q(\wbPeripheralBusInterface.state[0] ));
 sky130_fd_sc_hd__dfxtp_4 _2847_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_0058_),
    .Q(\wbPeripheralBusInterface.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2848_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net543),
    .Q(\vga.stateRegister.baseReadData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2849_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0060_),
    .Q(\vga.stateRegister.baseReadData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2850_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0061_),
    .Q(\vga.stateRegister.baseReadData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2851_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0062_),
    .Q(\vga.stateRegister.baseReadData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2852_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0063_),
    .Q(\vga.stateRegister.baseReadData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2853_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_0064_),
    .Q(\vga.raw_directPixelCounterVertical[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2854_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_0065_),
    .Q(\vga.raw_directPixelCounterVertical[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2855_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_0066_),
    .Q(\vga.raw_directPixelCounterVertical[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2856_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0067_),
    .Q(\vga.raw_directPixelCounterVertical[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2857_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0068_),
    .Q(\vga.raw_directPixelCounterVertical[4] ));
 sky130_fd_sc_hd__dfxtp_4 _2858_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0069_),
    .Q(\vga.raw_directPixelCounterVertical[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2859_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0070_),
    .Q(\vga.raw_directPixelCounterVertical[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2860_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0071_),
    .Q(\vga.raw_directPixelCounterVertical[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2861_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0072_),
    .Q(\vga.raw_directPixelCounterVertical[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2862_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0073_),
    .Q(\vga.raw_directPixelCounterVertical[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2863_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0074_),
    .Q(\vga.raw_directPixelCounterVertical[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2864_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0075_),
    .Q(\wbPeripheralBusInterface.currentByteSelect[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2865_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0076_),
    .Q(\wbPeripheralBusInterface.currentByteSelect[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2866_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_0077_),
    .Q(\wbPeripheralBusInterface.currentByteSelect[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2867_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_0078_),
    .Q(\wbPeripheralBusInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2868_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_0079_),
    .Q(\vga.raw_verticalPixelStretchCounter[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2869_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_0080_),
    .Q(\vga.raw_verticalPixelStretchCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2870_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_0081_),
    .Q(\vga.raw_verticalPixelStretchCounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2871_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_0082_),
    .Q(\vga.raw_verticalPixelStretchCounter[3] ));
 sky130_fd_sc_hd__dfxtp_4 _2872_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0083_),
    .Q(\vga.raw_subPixelCounter_buffered[0] ));
 sky130_fd_sc_hd__dfxtp_4 _2873_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0084_),
    .Q(\vga.raw_subPixelCounter_buffered[1] ));
 sky130_fd_sc_hd__dfxtp_4 _2874_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0085_),
    .Q(\vga.raw_subPixelCounter_buffered[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2875_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_0086_),
    .Q(\vga.raw_verticalPixelCounter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2876_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_0087_),
    .Q(\vga.raw_verticalPixelCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2877_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0088_),
    .Q(\vga.raw_verticalPixelCounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2878_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0089_),
    .Q(\vga.raw_verticalPixelCounter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2879_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0090_),
    .Q(\vga.raw_verticalPixelCounter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2880_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0091_),
    .Q(\vga.raw_verticalPixelCounter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2881_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0092_),
    .Q(\vga.raw_verticalPixelCounter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2882_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0093_),
    .Q(\vga.raw_verticalPixelCounter[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2883_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0094_),
    .Q(\vga.raw_verticalPixelCounter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2884_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0095_),
    .Q(\vga.raw_verticalPixelCounter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2885_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0096_),
    .Q(\vga.raw_subPixelCounter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2886_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0097_),
    .Q(\vga.raw_subPixelCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2887_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0098_),
    .Q(\vga.raw_subPixelCounter[2] ));
 sky130_fd_sc_hd__dfxtp_4 _2888_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0099_),
    .Q(\vga.raw_horizontalPixelCounter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _2889_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_0100_),
    .Q(\vga.raw_horizontalPixelCounter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2890_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_0101_),
    .Q(\vga.raw_horizontalPixelCounter[2] ));
 sky130_fd_sc_hd__dfxtp_4 _2891_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0102_),
    .Q(\vga.raw_horizontalPixelCounter[3] ));
 sky130_fd_sc_hd__dfxtp_4 _2892_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0103_),
    .Q(\vga.raw_horizontalPixelCounter[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2893_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0104_),
    .Q(\vga.raw_horizontalPixelCounter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2894_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0105_),
    .Q(\vga.raw_horizontalPixelCounter[6] ));
 sky130_fd_sc_hd__dfxtp_4 _2895_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0106_),
    .Q(\vga.raw_horizontalPixelCounter[7] ));
 sky130_fd_sc_hd__dfxtp_4 _2896_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0107_),
    .Q(\vga.raw_horizontalPixelCounter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2897_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_0108_),
    .Q(\vga.lastHSync ));
 sky130_fd_sc_hd__dfxtp_1 _2898_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_0109_),
    .Q(\vga.lastVSync ));
 sky130_fd_sc_hd__dfxtp_4 _2899_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0110_),
    .Q(\vga.raw_horizontalPixelStretchCounter[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2900_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0111_),
    .Q(\vga.raw_horizontalPixelStretchCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2901_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0112_),
    .Q(\vga.raw_horizontalPixelStretchCounter[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2902_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0113_),
    .Q(\vga.raw_horizontalPixelStretchCounter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2903_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0114_),
    .Q(\vga.currentPixelData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2904_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0115_),
    .Q(\vga.currentPixelData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2905_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0116_),
    .Q(\vga.currentPixelData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2906_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0117_),
    .Q(\vga.currentPixelData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2907_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0118_),
    .Q(\vga.currentPixelData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2908_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0119_),
    .Q(\vga.currentPixelData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2909_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0120_),
    .Q(\vga.currentPixelData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2910_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0121_),
    .Q(\vga.currentPixelData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2911_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0122_),
    .Q(\vga.currentPixelData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2912_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0123_),
    .Q(\vga.currentPixelData[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2913_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0124_),
    .Q(\vga.currentPixelData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2914_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0125_),
    .Q(\vga.currentPixelData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2915_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0126_),
    .Q(\vga.currentPixelData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2916_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0127_),
    .Q(\vga.currentPixelData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2917_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0128_),
    .Q(\vga.currentPixelData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2918_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0129_),
    .Q(\vga.currentPixelData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2919_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0130_),
    .Q(\vga.currentPixelData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2920_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0131_),
    .Q(\vga.currentPixelData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2921_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0132_),
    .Q(\vga.currentPixelData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2922_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0133_),
    .Q(\vga.currentPixelData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2923_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0134_),
    .Q(\vga.currentPixelData[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2924_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0135_),
    .Q(\vga.currentPixelData[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2925_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0136_),
    .Q(\vga.currentPixelData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2926_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0137_),
    .Q(\vga.currentPixelData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2927_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0138_),
    .Q(\vga.currentPixelData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2928_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0139_),
    .Q(\vga.currentPixelData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2929_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0140_),
    .Q(\vga.currentPixelData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2930_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0141_),
    .Q(\vga.currentPixelData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2931_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0142_),
    .Q(\vga.currentPixelData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2932_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0143_),
    .Q(\vga.currentPixelData[29] ));
 sky130_fd_sc_hd__dfxtp_4 _2933_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0144_),
    .Q(\vga.inVerticalVisibleArea ));
 sky130_fd_sc_hd__dfxtp_4 _2934_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0145_),
    .Q(\vga.verticalCounter[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2935_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0146_),
    .Q(\vga.verticalCounter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2936_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0147_),
    .Q(\vga.verticalCounter[2] ));
 sky130_fd_sc_hd__dfxtp_4 _2937_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0148_),
    .Q(\vga.verticalCounter[3] ));
 sky130_fd_sc_hd__dfxtp_4 _2938_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0149_),
    .Q(\vga.verticalCounter[4] ));
 sky130_fd_sc_hd__dfxtp_4 _2939_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0150_),
    .Q(\vga.verticalCounter[5] ));
 sky130_fd_sc_hd__dfxtp_4 _2940_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0151_),
    .Q(\vga.verticalCounter[6] ));
 sky130_fd_sc_hd__dfxtp_4 _2941_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0152_),
    .Q(\vga.verticalCounter[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2942_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0153_),
    .Q(\vga.verticalCounter[8] ));
 sky130_fd_sc_hd__dfxtp_4 _2943_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0154_),
    .Q(\vga.verticalCounter[9] ));
 sky130_fd_sc_hd__dfxtp_2 _2944_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0155_),
    .Q(\vga.vsync ));
 sky130_fd_sc_hd__dfxtp_1 _2945_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0156_),
    .Q(\vga.inHorizontalVisibleArea ));
 sky130_fd_sc_hd__dfxtp_1 _2946_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0157_),
    .Q(\vga.loadPixelData ));
 sky130_fd_sc_hd__dfxtp_4 _2947_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0158_),
    .Q(\vga.hsync ));
 sky130_fd_sc_hd__dfxtp_4 _2948_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0159_),
    .Q(\vga.horizontalCounter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _2949_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0160_),
    .Q(\vga.horizontalCounter[1] ));
 sky130_fd_sc_hd__dfxtp_4 _2950_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0161_),
    .Q(\vga.horizontalCounter[2] ));
 sky130_fd_sc_hd__dfxtp_4 _2951_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0162_),
    .Q(\vga.horizontalCounter[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2952_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0163_),
    .Q(\vga.horizontalCounter[4] ));
 sky130_fd_sc_hd__dfxtp_4 _2953_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0164_),
    .Q(\vga.horizontalCounter[5] ));
 sky130_fd_sc_hd__dfxtp_4 _2954_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0165_),
    .Q(\vga.horizontalCounter[6] ));
 sky130_fd_sc_hd__dfxtp_2 _2955_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0166_),
    .Q(\vga.horizontalCounter[7] ));
 sky130_fd_sc_hd__dfxtp_4 _2956_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0167_),
    .Q(\vga.horizontalCounter[8] ));
 sky130_fd_sc_hd__dfxtp_2 _2957_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0168_),
    .Q(\vga.horizontalCounter[9] ));
 sky130_fd_sc_hd__dfxtp_2 _2958_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0169_),
    .Q(\vga.horizontalCounter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2959_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_0170_),
    .Q(\vga.configuration[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2960_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_0171_),
    .Q(\vga.configuration[11] ));
 sky130_fd_sc_hd__dfxtp_4 _2961_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_0172_),
    .Q(\vga.configuration[10] ));
 sky130_fd_sc_hd__dfxtp_2 _2962_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_0173_),
    .Q(\vga.configuration[9] ));
 sky130_fd_sc_hd__dfxtp_4 _2963_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_0174_),
    .Q(\vga.configuration[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2964_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_0175_),
    .Q(\vga.configuration[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2965_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0176_),
    .Q(\vga.configuration[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2966_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0177_),
    .Q(\vga.configuration[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2967_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0178_),
    .Q(\vga.configuration[4] ));
 sky130_fd_sc_hd__dfxtp_4 _2968_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0179_),
    .Q(\vga.configuration[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2969_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0180_),
    .Q(\vga.configuration[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2970_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0181_),
    .Q(\vga.configuration[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2971_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0182_),
    .Q(\vga.configuration[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2972_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0183_),
    .Q(\vga.horizontalVisibleAreaCompare[10] ));
 sky130_fd_sc_hd__dfxtp_2 _2973_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0184_),
    .Q(\vga.horizontalVisibleAreaCompare[9] ));
 sky130_fd_sc_hd__dfxtp_2 _2974_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0185_),
    .Q(\vga.horizontalVisibleAreaCompare[8] ));
 sky130_fd_sc_hd__dfxtp_4 _2975_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_0186_),
    .Q(\vga.horizontalVisibleAreaCompare[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2976_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_0187_),
    .Q(\vga.horizontalVisibleAreaCompare[6] ));
 sky130_fd_sc_hd__dfxtp_2 _2977_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_0188_),
    .Q(\vga.horizontalVisibleAreaCompare[5] ));
 sky130_fd_sc_hd__dfxtp_2 _2978_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_0189_),
    .Q(\vga.horizontalVisibleAreaCompare[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2979_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0190_),
    .Q(\vga.horizontalVisibleAreaCompare[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2980_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_0191_),
    .Q(\vga.horizontalVisibleAreaCompare[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2981_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0192_),
    .Q(\vga.horizontalVisibleAreaCompare[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2982_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_0193_),
    .Q(\vga.horizontalVisibleAreaCompare[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2983_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0194_),
    .Q(\vga.horizontalFrontPorchCompare[10] ));
 sky130_fd_sc_hd__dfxtp_2 _2984_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_0195_),
    .Q(\vga.horizontalFrontPorchCompare[9] ));
 sky130_fd_sc_hd__dfxtp_2 _2985_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_0196_),
    .Q(\vga.horizontalFrontPorchCompare[8] ));
 sky130_fd_sc_hd__dfxtp_2 _2986_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0197_),
    .Q(\vga.horizontalFrontPorchCompare[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2987_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0198_),
    .Q(\vga.horizontalFrontPorchCompare[6] ));
 sky130_fd_sc_hd__dfxtp_2 _2988_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0199_),
    .Q(\vga.horizontalFrontPorchCompare[5] ));
 sky130_fd_sc_hd__dfxtp_2 _2989_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0200_),
    .Q(\vga.horizontalFrontPorchCompare[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2990_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0201_),
    .Q(\vga.horizontalFrontPorchCompare[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2991_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0202_),
    .Q(\vga.horizontalFrontPorchCompare[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2992_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0203_),
    .Q(\vga.horizontalFrontPorchCompare[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2993_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0204_),
    .Q(\vga.horizontalFrontPorchCompare[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2994_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0205_),
    .Q(\vga.horizontalSyncPulseCompare[10] ));
 sky130_fd_sc_hd__dfxtp_2 _2995_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0206_),
    .Q(\vga.horizontalSyncPulseCompare[9] ));
 sky130_fd_sc_hd__dfxtp_2 _2996_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0207_),
    .Q(\vga.horizontalSyncPulseCompare[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2997_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0208_),
    .Q(\vga.horizontalSyncPulseCompare[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2998_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0209_),
    .Q(\vga.horizontalSyncPulseCompare[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2999_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0210_),
    .Q(\vga.horizontalSyncPulseCompare[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3000_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0211_),
    .Q(\vga.horizontalSyncPulseCompare[4] ));
 sky130_fd_sc_hd__dfxtp_2 _3001_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0212_),
    .Q(\vga.horizontalSyncPulseCompare[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3002_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0213_),
    .Q(\vga.horizontalSyncPulseCompare[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3003_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0214_),
    .Q(\vga.horizontalSyncPulseCompare[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3004_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0215_),
    .Q(\vga.horizontalSyncPulseCompare[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3005_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0216_),
    .Q(\vga.horizontalWholeLineCompare[10] ));
 sky130_fd_sc_hd__dfxtp_2 _3006_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0217_),
    .Q(\vga.horizontalWholeLineCompare[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3007_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0218_),
    .Q(\vga.horizontalWholeLineCompare[8] ));
 sky130_fd_sc_hd__dfxtp_2 _3008_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0219_),
    .Q(\vga.horizontalWholeLineCompare[7] ));
 sky130_fd_sc_hd__dfxtp_2 _3009_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0220_),
    .Q(\vga.horizontalWholeLineCompare[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3010_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0221_),
    .Q(\vga.horizontalWholeLineCompare[5] ));
 sky130_fd_sc_hd__dfxtp_2 _3011_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0222_),
    .Q(\vga.horizontalWholeLineCompare[4] ));
 sky130_fd_sc_hd__dfxtp_2 _3012_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0223_),
    .Q(\vga.horizontalWholeLineCompare[3] ));
 sky130_fd_sc_hd__dfxtp_2 _3013_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0224_),
    .Q(\vga.horizontalWholeLineCompare[2] ));
 sky130_fd_sc_hd__dfxtp_2 _3014_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0225_),
    .Q(\vga.horizontalWholeLineCompare[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3015_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0226_),
    .Q(\vga.horizontalWholeLineCompare[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3016_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0227_),
    .Q(\vga.verticalVisibleAreaCompare[9] ));
 sky130_fd_sc_hd__dfxtp_2 _3017_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0228_),
    .Q(\vga.verticalVisibleAreaCompare[8] ));
 sky130_fd_sc_hd__dfxtp_2 _3018_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0229_),
    .Q(\vga.verticalVisibleAreaCompare[7] ));
 sky130_fd_sc_hd__dfxtp_2 _3019_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0230_),
    .Q(\vga.verticalVisibleAreaCompare[6] ));
 sky130_fd_sc_hd__dfxtp_2 _3020_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0231_),
    .Q(\vga.verticalVisibleAreaCompare[5] ));
 sky130_fd_sc_hd__dfxtp_2 _3021_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0232_),
    .Q(\vga.verticalVisibleAreaCompare[4] ));
 sky130_fd_sc_hd__dfxtp_2 _3022_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0233_),
    .Q(\vga.verticalVisibleAreaCompare[3] ));
 sky130_fd_sc_hd__dfxtp_2 _3023_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0234_),
    .Q(\vga.verticalVisibleAreaCompare[2] ));
 sky130_fd_sc_hd__dfxtp_2 _3024_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0235_),
    .Q(\vga.verticalVisibleAreaCompare[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3025_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0236_),
    .Q(\vga.verticalVisibleAreaCompare[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3026_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0237_),
    .Q(\vga.verticalFrontPorchCompare[9] ));
 sky130_fd_sc_hd__dfxtp_2 _3027_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0238_),
    .Q(\vga.verticalFrontPorchCompare[8] ));
 sky130_fd_sc_hd__dfxtp_2 _3028_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0239_),
    .Q(\vga.verticalFrontPorchCompare[7] ));
 sky130_fd_sc_hd__dfxtp_2 _3029_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0240_),
    .Q(\vga.verticalFrontPorchCompare[6] ));
 sky130_fd_sc_hd__dfxtp_2 _3030_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0241_),
    .Q(\vga.verticalFrontPorchCompare[5] ));
 sky130_fd_sc_hd__dfxtp_2 _3031_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0242_),
    .Q(\vga.verticalFrontPorchCompare[4] ));
 sky130_fd_sc_hd__dfxtp_2 _3032_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0243_),
    .Q(\vga.verticalFrontPorchCompare[3] ));
 sky130_fd_sc_hd__dfxtp_2 _3033_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0244_),
    .Q(\vga.verticalFrontPorchCompare[2] ));
 sky130_fd_sc_hd__dfxtp_2 _3034_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0245_),
    .Q(\vga.verticalFrontPorchCompare[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3035_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0246_),
    .Q(\vga.verticalFrontPorchCompare[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3036_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0247_),
    .Q(\vga.verticalSyncPulseCompare[9] ));
 sky130_fd_sc_hd__dfxtp_2 _3037_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0248_),
    .Q(\vga.verticalSyncPulseCompare[8] ));
 sky130_fd_sc_hd__dfxtp_2 _3038_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0249_),
    .Q(\vga.verticalSyncPulseCompare[7] ));
 sky130_fd_sc_hd__dfxtp_2 _3039_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0250_),
    .Q(\vga.verticalSyncPulseCompare[6] ));
 sky130_fd_sc_hd__dfxtp_2 _3040_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0251_),
    .Q(\vga.verticalSyncPulseCompare[5] ));
 sky130_fd_sc_hd__dfxtp_2 _3041_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0252_),
    .Q(\vga.verticalSyncPulseCompare[4] ));
 sky130_fd_sc_hd__dfxtp_2 _3042_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0253_),
    .Q(\vga.verticalSyncPulseCompare[3] ));
 sky130_fd_sc_hd__dfxtp_2 _3043_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0254_),
    .Q(\vga.verticalSyncPulseCompare[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3044_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0255_),
    .Q(\vga.verticalSyncPulseCompare[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3045_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0256_),
    .Q(\vga.verticalSyncPulseCompare[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3046_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0257_),
    .Q(\vga.verticalWholeLineCompare[9] ));
 sky130_fd_sc_hd__dfxtp_2 _3047_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0258_),
    .Q(\vga.verticalWholeLineCompare[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3048_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0259_),
    .Q(\vga.verticalWholeLineCompare[7] ));
 sky130_fd_sc_hd__dfxtp_2 _3049_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0260_),
    .Q(\vga.verticalWholeLineCompare[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3050_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0261_),
    .Q(\vga.verticalWholeLineCompare[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3051_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0262_),
    .Q(\vga.verticalWholeLineCompare[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3052_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0263_),
    .Q(\vga.verticalWholeLineCompare[3] ));
 sky130_fd_sc_hd__dfxtp_2 _3053_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0264_),
    .Q(\vga.verticalWholeLineCompare[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3054_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0265_),
    .Q(\vga.verticalWholeLineCompare[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3055_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0266_),
    .Q(\vga.verticalWholeLineCompare[0] ));
 sky130_fd_sc_hd__buf_2 _3057_ (.A(clknet_leaf_4_wb_clk_i),
    .X(net329));
 sky130_fd_sc_hd__buf_2 _3058_ (.A(clknet_leaf_69_wb_clk_i),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 _3059_ (.A(net311),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 _3060_ (.A(net312),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 _3061_ (.A(net313),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 _3062_ (.A(net314),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_2 _3063_ (.A(net315),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_2 _3064_ (.A(net316),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 _3065_ (.A(net317),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_2 _3066_ (.A(net318),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_2 _3067_ (.A(net319),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_2 _3068_ (.A(net320),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_2 _3069_ (.A(net321),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_2 _3070_ (.A(net322),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_2 _3071_ (.A(net323),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_2 _3072_ (.A(net324),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_2 _3073_ (.A(net325),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 _3074_ (.A(net326),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_2 _3075_ (.A(net327),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 _3076_ (.A(net328),
    .X(net389));
 sky130_fd_sc_hd__buf_2 _3077_ (.A(clknet_leaf_39_wb_clk_i),
    .X(net390));
 sky130_fd_sc_hd__buf_2 _3078_ (.A(clknet_leaf_43_wb_clk_i),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_2 _3079_ (.A(net335),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_2 _3080_ (.A(net346),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 _3081_ (.A(net357),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_2 _3082_ (.A(net360),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_2 _3083_ (.A(net361),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_2 _3084_ (.A(net362),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 _3085_ (.A(net363),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_2 _3086_ (.A(net364),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_2 _3087_ (.A(net365),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_2 _3088_ (.A(net366),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_2 _3089_ (.A(net336),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 _3090_ (.A(net337),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_2 _3091_ (.A(net338),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_2 _3092_ (.A(net339),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_2 _3093_ (.A(net340),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_2 _3094_ (.A(net341),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_2 _3095_ (.A(net342),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_2 _3096_ (.A(net343),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 _3097_ (.A(net344),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_2 _3098_ (.A(net345),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_2 _3099_ (.A(net347),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_2 _3100_ (.A(net348),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_2 _3101_ (.A(net349),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_2 _3102_ (.A(net350),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_2 _3103_ (.A(net351),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_2 _3104_ (.A(net352),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_2 _3105_ (.A(net353),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_2 _3106_ (.A(net354),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_2 _3107_ (.A(net355),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_2 _3108_ (.A(net356),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_2 _3109_ (.A(net358),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_2 _3110_ (.A(net359),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_2 _3111_ (.A(net367),
    .X(net428));
 sky130_fd_sc_hd__buf_2 _3112_ (.A(net566),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_4 _3113_ (.A(net573),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 _3114_ (.A(net370),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_2 _3115_ (.A(net371),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_51_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_52_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_53_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_54_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_55_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_56_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_57_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_58_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_59_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_60_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_61_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_62_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_63_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_64_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_65_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_66_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_67_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_68_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_69_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__buf_4 fanout477 (.A(net480),
    .X(net477));
 sky130_fd_sc_hd__buf_4 fanout478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__buf_4 fanout479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__buf_2 fanout480 (.A(_0475_),
    .X(net480));
 sky130_fd_sc_hd__buf_2 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_2 fanout482 (.A(_0474_),
    .X(net482));
 sky130_fd_sc_hd__buf_4 fanout483 (.A(net486),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_2 fanout484 (.A(net486),
    .X(net484));
 sky130_fd_sc_hd__buf_4 fanout485 (.A(net486),
    .X(net485));
 sky130_fd_sc_hd__buf_2 fanout486 (.A(net488),
    .X(net486));
 sky130_fd_sc_hd__buf_2 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_2 fanout488 (.A(_0474_),
    .X(net488));
 sky130_fd_sc_hd__buf_2 fanout489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_4 fanout490 (.A(net491),
    .X(net490));
 sky130_fd_sc_hd__buf_2 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__buf_4 fanout492 (.A(_0473_),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_4 fanout493 (.A(net496),
    .X(net493));
 sky130_fd_sc_hd__buf_2 fanout494 (.A(net495),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_4 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__buf_2 fanout496 (.A(_0466_),
    .X(net496));
 sky130_fd_sc_hd__buf_4 fanout497 (.A(net500),
    .X(net497));
 sky130_fd_sc_hd__buf_2 fanout498 (.A(net500),
    .X(net498));
 sky130_fd_sc_hd__buf_4 fanout499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_4 fanout500 (.A(_0465_),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_4 fanout501 (.A(net504),
    .X(net501));
 sky130_fd_sc_hd__buf_2 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_4 fanout503 (.A(net504),
    .X(net503));
 sky130_fd_sc_hd__buf_2 fanout504 (.A(_0468_),
    .X(net504));
 sky130_fd_sc_hd__buf_4 fanout505 (.A(net508),
    .X(net505));
 sky130_fd_sc_hd__buf_2 fanout506 (.A(net508),
    .X(net506));
 sky130_fd_sc_hd__buf_4 fanout507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_4 fanout508 (.A(_0467_),
    .X(net508));
 sky130_fd_sc_hd__buf_6 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_6 fanout510 (.A(_0785_),
    .X(net510));
 sky130_fd_sc_hd__buf_4 fanout511 (.A(_1281_),
    .X(net511));
 sky130_fd_sc_hd__buf_4 fanout512 (.A(_1229_),
    .X(net512));
 sky130_fd_sc_hd__buf_4 fanout513 (.A(_0589_),
    .X(net513));
 sky130_fd_sc_hd__buf_4 fanout514 (.A(_0564_),
    .X(net514));
 sky130_fd_sc_hd__buf_4 fanout515 (.A(_0563_),
    .X(net515));
 sky130_fd_sc_hd__buf_4 fanout516 (.A(_0558_),
    .X(net516));
 sky130_fd_sc_hd__buf_4 fanout517 (.A(_0548_),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_8 fanout518 (.A(_0547_),
    .X(net518));
 sky130_fd_sc_hd__buf_4 fanout519 (.A(_0544_),
    .X(net519));
 sky130_fd_sc_hd__buf_4 fanout520 (.A(_0538_),
    .X(net520));
 sky130_fd_sc_hd__buf_4 fanout521 (.A(_0529_),
    .X(net521));
 sky130_fd_sc_hd__buf_6 fanout522 (.A(net524),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_4 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_6 fanout524 (.A(net525),
    .X(net524));
 sky130_fd_sc_hd__buf_8 fanout525 (.A(_0521_),
    .X(net525));
 sky130_fd_sc_hd__buf_6 fanout526 (.A(_0520_),
    .X(net526));
 sky130_fd_sc_hd__buf_6 fanout527 (.A(_0520_),
    .X(net527));
 sky130_fd_sc_hd__buf_6 fanout528 (.A(net529),
    .X(net528));
 sky130_fd_sc_hd__buf_4 fanout529 (.A(_0330_),
    .X(net529));
 sky130_fd_sc_hd__buf_8 fanout530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__buf_12 fanout531 (.A(_0277_),
    .X(net531));
 sky130_fd_sc_hd__buf_6 fanout532 (.A(_0313_),
    .X(net532));
 sky130_fd_sc_hd__buf_6 fanout533 (.A(net535),
    .X(net533));
 sky130_fd_sc_hd__buf_6 fanout534 (.A(net535),
    .X(net534));
 sky130_fd_sc_hd__buf_6 fanout535 (.A(_0868_),
    .X(net535));
 sky130_fd_sc_hd__buf_4 fanout536 (.A(net538),
    .X(net536));
 sky130_fd_sc_hd__buf_2 fanout537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_16 fanout538 (.A(_0791_),
    .X(net538));
 sky130_fd_sc_hd__buf_4 fanout539 (.A(net540),
    .X(net539));
 sky130_fd_sc_hd__buf_4 fanout540 (.A(net543),
    .X(net540));
 sky130_fd_sc_hd__buf_4 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__buf_2 fanout542 (.A(net543),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_8 fanout543 (.A(_0059_),
    .X(net543));
 sky130_fd_sc_hd__buf_6 fanout544 (.A(_0282_),
    .X(net544));
 sky130_fd_sc_hd__buf_6 fanout545 (.A(net547),
    .X(net545));
 sky130_fd_sc_hd__buf_4 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_4 fanout547 (.A(_0282_),
    .X(net547));
 sky130_fd_sc_hd__buf_4 fanout548 (.A(net552),
    .X(net548));
 sky130_fd_sc_hd__buf_6 fanout549 (.A(net551),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_4 fanout550 (.A(net551),
    .X(net550));
 sky130_fd_sc_hd__buf_2 fanout551 (.A(net552),
    .X(net551));
 sky130_fd_sc_hd__buf_2 fanout552 (.A(_0281_),
    .X(net552));
 sky130_fd_sc_hd__buf_4 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__buf_4 fanout554 (.A(_0280_),
    .X(net554));
 sky130_fd_sc_hd__buf_4 fanout555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__buf_4 fanout556 (.A(_0280_),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_4 fanout557 (.A(net558),
    .X(net557));
 sky130_fd_sc_hd__buf_6 fanout558 (.A(net559),
    .X(net558));
 sky130_fd_sc_hd__buf_4 fanout559 (.A(net560),
    .X(net559));
 sky130_fd_sc_hd__buf_4 fanout560 (.A(_0274_),
    .X(net560));
 sky130_fd_sc_hd__buf_4 fanout561 (.A(net564),
    .X(net561));
 sky130_fd_sc_hd__buf_6 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__buf_6 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__buf_8 fanout564 (.A(_0273_),
    .X(net564));
 sky130_fd_sc_hd__buf_4 fanout565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__buf_2 fanout566 (.A(net572),
    .X(net566));
 sky130_fd_sc_hd__buf_4 fanout567 (.A(net572),
    .X(net567));
 sky130_fd_sc_hd__buf_4 fanout568 (.A(net572),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_4 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_4 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_4 fanout571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__buf_4 fanout572 (.A(net368),
    .X(net572));
 sky130_fd_sc_hd__buf_6 fanout573 (.A(net369),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_2 fanout574 (.A(net369),
    .X(net574));
 sky130_fd_sc_hd__buf_6 fanout575 (.A(_0463_),
    .X(net575));
 sky130_fd_sc_hd__buf_6 fanout576 (.A(_0312_),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_16 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__buf_12 fanout578 (.A(_0276_),
    .X(net578));
 sky130_fd_sc_hd__buf_4 fanout579 (.A(_0275_),
    .X(net579));
 sky130_fd_sc_hd__buf_12 fanout580 (.A(_1354_),
    .X(net580));
 sky130_fd_sc_hd__buf_6 fanout581 (.A(_1354_),
    .X(net581));
 sky130_fd_sc_hd__buf_4 fanout582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__buf_6 fanout583 (.A(net584),
    .X(net583));
 sky130_fd_sc_hd__buf_6 fanout584 (.A(_1351_),
    .X(net584));
 sky130_fd_sc_hd__buf_4 fanout585 (.A(_1351_),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_4 fanout586 (.A(_1351_),
    .X(net586));
 sky130_fd_sc_hd__buf_4 fanout587 (.A(_1328_),
    .X(net587));
 sky130_fd_sc_hd__buf_2 fanout588 (.A(_1328_),
    .X(net588));
 sky130_fd_sc_hd__buf_4 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_4 fanout590 (.A(_1328_),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_4 fanout591 (.A(net594),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_4 fanout592 (.A(net593),
    .X(net592));
 sky130_fd_sc_hd__buf_4 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_4 fanout594 (.A(\vga.loadPixelData ),
    .X(net594));
 sky130_fd_sc_hd__buf_6 fanout595 (.A(\vga.raw_horizontalPixelCounter[0] ),
    .X(net595));
 sky130_fd_sc_hd__buf_4 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__buf_4 fanout597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__buf_4 fanout598 (.A(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_16 fanout599 (.A(net601),
    .X(net599));
 sky130_fd_sc_hd__buf_4 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__buf_8 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_6 fanout602 (.A(\wbPeripheralBusInterface.currentByteSelect[0] ),
    .X(net602));
 sky130_fd_sc_hd__buf_4 fanout603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_4 fanout604 (.A(net609),
    .X(net604));
 sky130_fd_sc_hd__buf_6 fanout605 (.A(net609),
    .X(net605));
 sky130_fd_sc_hd__buf_6 fanout606 (.A(net609),
    .X(net606));
 sky130_fd_sc_hd__buf_4 fanout607 (.A(net609),
    .X(net607));
 sky130_fd_sc_hd__buf_6 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__buf_12 fanout609 (.A(_1331_),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_8 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__buf_4 fanout611 (.A(net613),
    .X(net611));
 sky130_fd_sc_hd__buf_4 fanout612 (.A(net613),
    .X(net612));
 sky130_fd_sc_hd__buf_8 fanout613 (.A(net618),
    .X(net613));
 sky130_fd_sc_hd__buf_6 fanout614 (.A(net618),
    .X(net614));
 sky130_fd_sc_hd__buf_4 fanout615 (.A(net618),
    .X(net615));
 sky130_fd_sc_hd__buf_4 fanout616 (.A(net618),
    .X(net616));
 sky130_fd_sc_hd__buf_4 fanout617 (.A(net618),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_16 fanout618 (.A(net304),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(sram0_dout0[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(sram0_dout0[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input100 (.A(sram0_dout1[43]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 input101 (.A(sram0_dout1[44]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 input102 (.A(sram0_dout1[45]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(sram0_dout1[46]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 input104 (.A(sram0_dout1[47]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 input105 (.A(sram0_dout1[48]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 input106 (.A(sram0_dout1[49]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 input107 (.A(sram0_dout1[4]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 input108 (.A(sram0_dout1[50]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 input109 (.A(sram0_dout1[51]),
    .X(net109));
 sky130_fd_sc_hd__buf_2 input11 (.A(sram0_dout0[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input110 (.A(sram0_dout1[52]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 input111 (.A(sram0_dout1[53]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 input112 (.A(sram0_dout1[54]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 input113 (.A(sram0_dout1[55]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 input114 (.A(sram0_dout1[56]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 input115 (.A(sram0_dout1[57]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 input116 (.A(sram0_dout1[58]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 input117 (.A(sram0_dout1[59]),
    .X(net117));
 sky130_fd_sc_hd__buf_4 input118 (.A(sram0_dout1[5]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 input119 (.A(sram0_dout1[60]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(sram0_dout0[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input120 (.A(sram0_dout1[61]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 input121 (.A(sram0_dout1[6]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 input122 (.A(sram0_dout1[7]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 input123 (.A(sram0_dout1[8]),
    .X(net123));
 sky130_fd_sc_hd__buf_4 input124 (.A(sram0_dout1[9]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(sram1_dout0[0]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(sram1_dout0[10]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(sram1_dout0[11]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(sram1_dout0[12]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(sram1_dout0[13]),
    .X(net129));
 sky130_fd_sc_hd__buf_2 input13 (.A(sram0_dout0[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(sram1_dout0[14]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(sram1_dout0[15]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(sram1_dout0[16]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(sram1_dout0[17]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input134 (.A(sram1_dout0[18]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(sram1_dout0[19]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(sram1_dout0[1]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 input137 (.A(sram1_dout0[20]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 input138 (.A(sram1_dout0[21]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 input139 (.A(sram1_dout0[22]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(sram0_dout0[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input140 (.A(sram1_dout0[23]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 input141 (.A(sram1_dout0[24]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(sram1_dout0[25]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(sram1_dout0[26]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 input144 (.A(sram1_dout0[27]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(sram1_dout0[28]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 input146 (.A(sram1_dout0[29]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(sram1_dout0[2]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 input148 (.A(sram1_dout0[30]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 input149 (.A(sram1_dout0[31]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(sram0_dout0[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input150 (.A(sram1_dout0[32]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 input151 (.A(sram1_dout0[33]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 input152 (.A(sram1_dout0[34]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 input153 (.A(sram1_dout0[35]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 input154 (.A(sram1_dout0[36]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 input155 (.A(sram1_dout0[37]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 input156 (.A(sram1_dout0[38]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 input157 (.A(sram1_dout0[39]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 input158 (.A(sram1_dout0[3]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 input159 (.A(sram1_dout0[40]),
    .X(net159));
 sky130_fd_sc_hd__buf_2 input16 (.A(sram0_dout0[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input160 (.A(sram1_dout0[41]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 input161 (.A(sram1_dout0[42]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 input162 (.A(sram1_dout0[43]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 input163 (.A(sram1_dout0[44]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 input164 (.A(sram1_dout0[45]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 input165 (.A(sram1_dout0[46]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 input166 (.A(sram1_dout0[47]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 input167 (.A(sram1_dout0[48]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 input168 (.A(sram1_dout0[49]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 input169 (.A(sram1_dout0[4]),
    .X(net169));
 sky130_fd_sc_hd__buf_2 input17 (.A(sram0_dout0[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input170 (.A(sram1_dout0[50]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 input171 (.A(sram1_dout0[51]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(sram1_dout0[52]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 input173 (.A(sram1_dout0[53]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 input174 (.A(sram1_dout0[54]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 input175 (.A(sram1_dout0[55]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 input176 (.A(sram1_dout0[56]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 input177 (.A(sram1_dout0[57]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 input178 (.A(sram1_dout0[58]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 input179 (.A(sram1_dout0[59]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(sram0_dout0[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(sram1_dout0[5]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 input181 (.A(sram1_dout0[60]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 input182 (.A(sram1_dout0[61]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 input183 (.A(sram1_dout0[62]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 input184 (.A(sram1_dout0[63]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 input185 (.A(sram1_dout0[6]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(sram1_dout0[7]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 input187 (.A(sram1_dout0[8]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 input188 (.A(sram1_dout0[9]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 input189 (.A(sram1_dout1[0]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(sram0_dout0[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(sram1_dout1[10]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 input191 (.A(sram1_dout1[11]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 input192 (.A(sram1_dout1[12]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_2 input193 (.A(sram1_dout1[13]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 input194 (.A(sram1_dout1[14]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input195 (.A(sram1_dout1[15]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 input196 (.A(sram1_dout1[16]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 input197 (.A(sram1_dout1[17]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(sram1_dout1[18]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 input199 (.A(sram1_dout1[19]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(sram0_dout0[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(sram0_dout0[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input200 (.A(sram1_dout1[1]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 input201 (.A(sram1_dout1[20]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 input202 (.A(sram1_dout1[21]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 input203 (.A(sram1_dout1[22]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 input204 (.A(sram1_dout1[23]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 input205 (.A(sram1_dout1[24]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 input206 (.A(sram1_dout1[25]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 input207 (.A(sram1_dout1[26]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 input208 (.A(sram1_dout1[27]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 input209 (.A(sram1_dout1[28]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(sram0_dout0[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input210 (.A(sram1_dout1[29]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 input211 (.A(sram1_dout1[2]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 input212 (.A(sram1_dout1[32]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(sram1_dout1[33]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 input214 (.A(sram1_dout1[34]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 input215 (.A(sram1_dout1[35]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 input216 (.A(sram1_dout1[36]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 input217 (.A(sram1_dout1[37]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 input218 (.A(sram1_dout1[38]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 input219 (.A(sram1_dout1[39]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(sram0_dout0[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input220 (.A(sram1_dout1[3]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_2 input221 (.A(sram1_dout1[40]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 input222 (.A(sram1_dout1[41]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 input223 (.A(sram1_dout1[42]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 input224 (.A(sram1_dout1[43]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 input225 (.A(sram1_dout1[44]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 input226 (.A(sram1_dout1[45]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 input227 (.A(sram1_dout1[46]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 input228 (.A(sram1_dout1[47]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 input229 (.A(sram1_dout1[48]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(sram0_dout0[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input230 (.A(sram1_dout1[49]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 input231 (.A(sram1_dout1[4]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 input232 (.A(sram1_dout1[50]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 input233 (.A(sram1_dout1[51]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 input234 (.A(sram1_dout1[52]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 input235 (.A(sram1_dout1[53]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 input236 (.A(sram1_dout1[54]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 input237 (.A(sram1_dout1[55]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 input238 (.A(sram1_dout1[56]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 input239 (.A(sram1_dout1[57]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(sram0_dout0[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input240 (.A(sram1_dout1[58]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 input241 (.A(sram1_dout1[59]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 input242 (.A(sram1_dout1[5]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 input243 (.A(sram1_dout1[60]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 input244 (.A(sram1_dout1[61]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 input245 (.A(sram1_dout1[6]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 input246 (.A(sram1_dout1[7]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 input247 (.A(sram1_dout1[8]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 input248 (.A(sram1_dout1[9]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 input249 (.A(wb_adr_i[10]),
    .X(net249));
 sky130_fd_sc_hd__buf_2 input25 (.A(sram0_dout0[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input250 (.A(wb_adr_i[11]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 input251 (.A(wb_adr_i[12]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_2 input252 (.A(wb_adr_i[13]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 input253 (.A(wb_adr_i[14]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 input254 (.A(wb_adr_i[15]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 input255 (.A(wb_adr_i[16]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_2 input256 (.A(wb_adr_i[17]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 input257 (.A(wb_adr_i[18]),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 input258 (.A(wb_adr_i[19]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 input259 (.A(wb_adr_i[20]),
    .X(net259));
 sky130_fd_sc_hd__buf_4 input26 (.A(sram0_dout0[32]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input260 (.A(wb_adr_i[21]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_2 input261 (.A(wb_adr_i[22]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 input262 (.A(wb_adr_i[23]),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 input263 (.A(wb_adr_i[2]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 input264 (.A(wb_adr_i[3]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 input265 (.A(wb_adr_i[4]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_2 input266 (.A(wb_adr_i[5]),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 input267 (.A(wb_adr_i[6]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 input268 (.A(wb_adr_i[7]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 input269 (.A(wb_adr_i[8]),
    .X(net269));
 sky130_fd_sc_hd__buf_4 input27 (.A(sram0_dout0[33]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input270 (.A(wb_adr_i[9]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 input271 (.A(wb_cyc_i),
    .X(net271));
 sky130_fd_sc_hd__buf_12 input272 (.A(wb_data_i[0]),
    .X(net272));
 sky130_fd_sc_hd__buf_6 input273 (.A(wb_data_i[10]),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 input274 (.A(wb_data_i[11]),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 input275 (.A(wb_data_i[12]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 input276 (.A(wb_data_i[13]),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_4 input277 (.A(wb_data_i[14]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 input278 (.A(wb_data_i[15]),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 input279 (.A(wb_data_i[16]),
    .X(net279));
 sky130_fd_sc_hd__buf_4 input28 (.A(sram0_dout0[34]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input280 (.A(wb_data_i[17]),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_4 input281 (.A(wb_data_i[18]),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_4 input282 (.A(wb_data_i[19]),
    .X(net282));
 sky130_fd_sc_hd__buf_12 input283 (.A(wb_data_i[1]),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_4 input284 (.A(wb_data_i[20]),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 input285 (.A(wb_data_i[21]),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_4 input286 (.A(wb_data_i[22]),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 input287 (.A(wb_data_i[23]),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 input288 (.A(wb_data_i[24]),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_4 input289 (.A(wb_data_i[25]),
    .X(net289));
 sky130_fd_sc_hd__buf_4 input29 (.A(sram0_dout0[35]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input290 (.A(wb_data_i[26]),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 input291 (.A(wb_data_i[27]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 input292 (.A(wb_data_i[28]),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 input293 (.A(wb_data_i[29]),
    .X(net293));
 sky130_fd_sc_hd__buf_12 input294 (.A(wb_data_i[2]),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 input295 (.A(wb_data_i[30]),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 input296 (.A(wb_data_i[31]),
    .X(net296));
 sky130_fd_sc_hd__buf_12 input297 (.A(wb_data_i[3]),
    .X(net297));
 sky130_fd_sc_hd__buf_12 input298 (.A(wb_data_i[4]),
    .X(net298));
 sky130_fd_sc_hd__buf_12 input299 (.A(wb_data_i[5]),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(sram0_dout0[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input30 (.A(sram0_dout0[36]),
    .X(net30));
 sky130_fd_sc_hd__buf_12 input300 (.A(wb_data_i[6]),
    .X(net300));
 sky130_fd_sc_hd__buf_12 input301 (.A(wb_data_i[7]),
    .X(net301));
 sky130_fd_sc_hd__buf_8 input302 (.A(wb_data_i[8]),
    .X(net302));
 sky130_fd_sc_hd__buf_8 input303 (.A(wb_data_i[9]),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_2 input304 (.A(wb_rst_i),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 input305 (.A(wb_sel_i[0]),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_2 input306 (.A(wb_sel_i[1]),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 input307 (.A(wb_sel_i[2]),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 input308 (.A(wb_sel_i[3]),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 input309 (.A(wb_stb_i),
    .X(net309));
 sky130_fd_sc_hd__buf_4 input31 (.A(sram0_dout0[37]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input310 (.A(wb_we_i),
    .X(net310));
 sky130_fd_sc_hd__buf_4 input32 (.A(sram0_dout0[38]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(sram0_dout0[39]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(sram0_dout0[3]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(sram0_dout0[40]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(sram0_dout0[41]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(sram0_dout0[42]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(sram0_dout0[43]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(sram0_dout0[44]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(sram0_dout0[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(sram0_dout0[45]),
    .X(net40));
 sky130_fd_sc_hd__buf_4 input41 (.A(sram0_dout0[46]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(sram0_dout0[47]),
    .X(net42));
 sky130_fd_sc_hd__buf_4 input43 (.A(sram0_dout0[48]),
    .X(net43));
 sky130_fd_sc_hd__buf_4 input44 (.A(sram0_dout0[49]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(sram0_dout0[4]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(sram0_dout0[50]),
    .X(net46));
 sky130_fd_sc_hd__buf_4 input47 (.A(sram0_dout0[51]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(sram0_dout0[52]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(sram0_dout0[53]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(sram0_dout0[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(sram0_dout0[54]),
    .X(net50));
 sky130_fd_sc_hd__buf_4 input51 (.A(sram0_dout0[55]),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(sram0_dout0[56]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(sram0_dout0[57]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(sram0_dout0[58]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(sram0_dout0[59]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(sram0_dout0[5]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(sram0_dout0[60]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(sram0_dout0[61]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(sram0_dout0[62]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(sram0_dout0[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input60 (.A(sram0_dout0[63]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(sram0_dout0[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(sram0_dout0[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(sram0_dout0[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(sram0_dout0[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 input65 (.A(sram0_dout1[0]),
    .X(net65));
 sky130_fd_sc_hd__buf_4 input66 (.A(sram0_dout1[10]),
    .X(net66));
 sky130_fd_sc_hd__buf_4 input67 (.A(sram0_dout1[11]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 input68 (.A(sram0_dout1[12]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(sram0_dout1[13]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(sram0_dout0[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input70 (.A(sram0_dout1[14]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 input71 (.A(sram0_dout1[15]),
    .X(net71));
 sky130_fd_sc_hd__buf_4 input72 (.A(sram0_dout1[16]),
    .X(net72));
 sky130_fd_sc_hd__buf_4 input73 (.A(sram0_dout1[17]),
    .X(net73));
 sky130_fd_sc_hd__buf_4 input74 (.A(sram0_dout1[18]),
    .X(net74));
 sky130_fd_sc_hd__buf_4 input75 (.A(sram0_dout1[19]),
    .X(net75));
 sky130_fd_sc_hd__buf_4 input76 (.A(sram0_dout1[1]),
    .X(net76));
 sky130_fd_sc_hd__buf_4 input77 (.A(sram0_dout1[20]),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input78 (.A(sram0_dout1[21]),
    .X(net78));
 sky130_fd_sc_hd__buf_4 input79 (.A(sram0_dout1[22]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input8 (.A(sram0_dout0[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input80 (.A(sram0_dout1[23]),
    .X(net80));
 sky130_fd_sc_hd__buf_4 input81 (.A(sram0_dout1[24]),
    .X(net81));
 sky130_fd_sc_hd__buf_4 input82 (.A(sram0_dout1[25]),
    .X(net82));
 sky130_fd_sc_hd__buf_4 input83 (.A(sram0_dout1[26]),
    .X(net83));
 sky130_fd_sc_hd__buf_4 input84 (.A(sram0_dout1[27]),
    .X(net84));
 sky130_fd_sc_hd__buf_4 input85 (.A(sram0_dout1[28]),
    .X(net85));
 sky130_fd_sc_hd__buf_4 input86 (.A(sram0_dout1[29]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(sram0_dout1[2]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 input88 (.A(sram0_dout1[32]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 input89 (.A(sram0_dout1[33]),
    .X(net89));
 sky130_fd_sc_hd__buf_2 input9 (.A(sram0_dout0[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input90 (.A(sram0_dout1[34]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(sram0_dout1[35]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(sram0_dout1[36]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(sram0_dout1[37]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 input94 (.A(sram0_dout1[38]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 input95 (.A(sram0_dout1[39]),
    .X(net95));
 sky130_fd_sc_hd__buf_4 input96 (.A(sram0_dout1[3]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 input97 (.A(sram0_dout1[40]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 input98 (.A(sram0_dout1[41]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 input99 (.A(sram0_dout1[42]),
    .X(net99));
 sky130_fd_sc_hd__buf_4 output311 (.A(net311),
    .X(sram0_addr0[0]));
 sky130_fd_sc_hd__buf_4 output312 (.A(net312),
    .X(sram0_addr0[1]));
 sky130_fd_sc_hd__buf_4 output313 (.A(net313),
    .X(sram0_addr0[2]));
 sky130_fd_sc_hd__buf_4 output314 (.A(net314),
    .X(sram0_addr0[3]));
 sky130_fd_sc_hd__buf_4 output315 (.A(net315),
    .X(sram0_addr0[4]));
 sky130_fd_sc_hd__buf_4 output316 (.A(net316),
    .X(sram0_addr0[5]));
 sky130_fd_sc_hd__buf_4 output317 (.A(net317),
    .X(sram0_addr0[6]));
 sky130_fd_sc_hd__buf_4 output318 (.A(net318),
    .X(sram0_addr0[7]));
 sky130_fd_sc_hd__buf_4 output319 (.A(net319),
    .X(sram0_addr0[8]));
 sky130_fd_sc_hd__buf_4 output320 (.A(net320),
    .X(sram0_addr1[0]));
 sky130_fd_sc_hd__buf_4 output321 (.A(net321),
    .X(sram0_addr1[1]));
 sky130_fd_sc_hd__buf_4 output322 (.A(net322),
    .X(sram0_addr1[2]));
 sky130_fd_sc_hd__buf_4 output323 (.A(net323),
    .X(sram0_addr1[3]));
 sky130_fd_sc_hd__buf_4 output324 (.A(net324),
    .X(sram0_addr1[4]));
 sky130_fd_sc_hd__buf_4 output325 (.A(net325),
    .X(sram0_addr1[5]));
 sky130_fd_sc_hd__buf_4 output326 (.A(net326),
    .X(sram0_addr1[6]));
 sky130_fd_sc_hd__buf_4 output327 (.A(net327),
    .X(sram0_addr1[7]));
 sky130_fd_sc_hd__buf_4 output328 (.A(net328),
    .X(sram0_addr1[8]));
 sky130_fd_sc_hd__clkbuf_2 output329 (.A(net329),
    .X(sram0_clk0));
 sky130_fd_sc_hd__clkbuf_2 output330 (.A(net330),
    .X(sram0_clk1));
 sky130_fd_sc_hd__buf_4 output331 (.A(net331),
    .X(sram0_csb0[0]));
 sky130_fd_sc_hd__buf_4 output332 (.A(net332),
    .X(sram0_csb0[1]));
 sky130_fd_sc_hd__buf_4 output333 (.A(net333),
    .X(sram0_csb1[0]));
 sky130_fd_sc_hd__buf_4 output334 (.A(net334),
    .X(sram0_csb1[1]));
 sky130_fd_sc_hd__buf_4 output335 (.A(net335),
    .X(sram0_din0[0]));
 sky130_fd_sc_hd__buf_4 output336 (.A(net336),
    .X(sram0_din0[10]));
 sky130_fd_sc_hd__buf_4 output337 (.A(net337),
    .X(sram0_din0[11]));
 sky130_fd_sc_hd__buf_4 output338 (.A(net338),
    .X(sram0_din0[12]));
 sky130_fd_sc_hd__buf_4 output339 (.A(net339),
    .X(sram0_din0[13]));
 sky130_fd_sc_hd__buf_4 output340 (.A(net340),
    .X(sram0_din0[14]));
 sky130_fd_sc_hd__buf_4 output341 (.A(net341),
    .X(sram0_din0[15]));
 sky130_fd_sc_hd__buf_4 output342 (.A(net342),
    .X(sram0_din0[16]));
 sky130_fd_sc_hd__buf_4 output343 (.A(net343),
    .X(sram0_din0[17]));
 sky130_fd_sc_hd__buf_4 output344 (.A(net344),
    .X(sram0_din0[18]));
 sky130_fd_sc_hd__buf_4 output345 (.A(net345),
    .X(sram0_din0[19]));
 sky130_fd_sc_hd__buf_4 output346 (.A(net346),
    .X(sram0_din0[1]));
 sky130_fd_sc_hd__buf_4 output347 (.A(net347),
    .X(sram0_din0[20]));
 sky130_fd_sc_hd__buf_4 output348 (.A(net348),
    .X(sram0_din0[21]));
 sky130_fd_sc_hd__buf_4 output349 (.A(net349),
    .X(sram0_din0[22]));
 sky130_fd_sc_hd__buf_4 output350 (.A(net350),
    .X(sram0_din0[23]));
 sky130_fd_sc_hd__buf_4 output351 (.A(net351),
    .X(sram0_din0[24]));
 sky130_fd_sc_hd__buf_4 output352 (.A(net352),
    .X(sram0_din0[25]));
 sky130_fd_sc_hd__buf_4 output353 (.A(net353),
    .X(sram0_din0[26]));
 sky130_fd_sc_hd__buf_4 output354 (.A(net354),
    .X(sram0_din0[27]));
 sky130_fd_sc_hd__buf_4 output355 (.A(net355),
    .X(sram0_din0[28]));
 sky130_fd_sc_hd__buf_4 output356 (.A(net356),
    .X(sram0_din0[29]));
 sky130_fd_sc_hd__buf_4 output357 (.A(net357),
    .X(sram0_din0[2]));
 sky130_fd_sc_hd__buf_4 output358 (.A(net358),
    .X(sram0_din0[30]));
 sky130_fd_sc_hd__buf_4 output359 (.A(net359),
    .X(sram0_din0[31]));
 sky130_fd_sc_hd__buf_4 output360 (.A(net360),
    .X(sram0_din0[3]));
 sky130_fd_sc_hd__buf_4 output361 (.A(net361),
    .X(sram0_din0[4]));
 sky130_fd_sc_hd__buf_4 output362 (.A(net362),
    .X(sram0_din0[5]));
 sky130_fd_sc_hd__buf_4 output363 (.A(net363),
    .X(sram0_din0[6]));
 sky130_fd_sc_hd__buf_4 output364 (.A(net364),
    .X(sram0_din0[7]));
 sky130_fd_sc_hd__buf_4 output365 (.A(net365),
    .X(sram0_din0[8]));
 sky130_fd_sc_hd__buf_4 output366 (.A(net366),
    .X(sram0_din0[9]));
 sky130_fd_sc_hd__buf_4 output367 (.A(net367),
    .X(sram0_web0));
 sky130_fd_sc_hd__buf_4 output368 (.A(net567),
    .X(sram0_wmask0[0]));
 sky130_fd_sc_hd__buf_4 output369 (.A(net573),
    .X(sram0_wmask0[1]));
 sky130_fd_sc_hd__buf_4 output370 (.A(net370),
    .X(sram0_wmask0[2]));
 sky130_fd_sc_hd__buf_4 output371 (.A(net371),
    .X(sram0_wmask0[3]));
 sky130_fd_sc_hd__buf_4 output372 (.A(net372),
    .X(sram1_addr0[0]));
 sky130_fd_sc_hd__buf_4 output373 (.A(net373),
    .X(sram1_addr0[1]));
 sky130_fd_sc_hd__buf_4 output374 (.A(net374),
    .X(sram1_addr0[2]));
 sky130_fd_sc_hd__buf_4 output375 (.A(net375),
    .X(sram1_addr0[3]));
 sky130_fd_sc_hd__buf_4 output376 (.A(net376),
    .X(sram1_addr0[4]));
 sky130_fd_sc_hd__buf_4 output377 (.A(net377),
    .X(sram1_addr0[5]));
 sky130_fd_sc_hd__buf_4 output378 (.A(net378),
    .X(sram1_addr0[6]));
 sky130_fd_sc_hd__buf_4 output379 (.A(net379),
    .X(sram1_addr0[7]));
 sky130_fd_sc_hd__buf_4 output380 (.A(net380),
    .X(sram1_addr0[8]));
 sky130_fd_sc_hd__buf_4 output381 (.A(net381),
    .X(sram1_addr1[0]));
 sky130_fd_sc_hd__buf_4 output382 (.A(net382),
    .X(sram1_addr1[1]));
 sky130_fd_sc_hd__buf_4 output383 (.A(net383),
    .X(sram1_addr1[2]));
 sky130_fd_sc_hd__buf_4 output384 (.A(net384),
    .X(sram1_addr1[3]));
 sky130_fd_sc_hd__buf_4 output385 (.A(net385),
    .X(sram1_addr1[4]));
 sky130_fd_sc_hd__buf_4 output386 (.A(net386),
    .X(sram1_addr1[5]));
 sky130_fd_sc_hd__buf_4 output387 (.A(net387),
    .X(sram1_addr1[6]));
 sky130_fd_sc_hd__buf_4 output388 (.A(net388),
    .X(sram1_addr1[7]));
 sky130_fd_sc_hd__buf_4 output389 (.A(net389),
    .X(sram1_addr1[8]));
 sky130_fd_sc_hd__clkbuf_2 output390 (.A(net390),
    .X(sram1_clk0));
 sky130_fd_sc_hd__clkbuf_2 output391 (.A(net391),
    .X(sram1_clk1));
 sky130_fd_sc_hd__buf_4 output392 (.A(net392),
    .X(sram1_csb0[0]));
 sky130_fd_sc_hd__buf_4 output393 (.A(net393),
    .X(sram1_csb0[1]));
 sky130_fd_sc_hd__buf_4 output394 (.A(net394),
    .X(sram1_csb1[0]));
 sky130_fd_sc_hd__buf_4 output395 (.A(net395),
    .X(sram1_csb1[1]));
 sky130_fd_sc_hd__buf_4 output396 (.A(net396),
    .X(sram1_din0[0]));
 sky130_fd_sc_hd__buf_4 output397 (.A(net397),
    .X(sram1_din0[10]));
 sky130_fd_sc_hd__buf_4 output398 (.A(net398),
    .X(sram1_din0[11]));
 sky130_fd_sc_hd__buf_4 output399 (.A(net399),
    .X(sram1_din0[12]));
 sky130_fd_sc_hd__buf_4 output400 (.A(net400),
    .X(sram1_din0[13]));
 sky130_fd_sc_hd__buf_4 output401 (.A(net401),
    .X(sram1_din0[14]));
 sky130_fd_sc_hd__buf_4 output402 (.A(net402),
    .X(sram1_din0[15]));
 sky130_fd_sc_hd__buf_4 output403 (.A(net403),
    .X(sram1_din0[16]));
 sky130_fd_sc_hd__buf_4 output404 (.A(net404),
    .X(sram1_din0[17]));
 sky130_fd_sc_hd__buf_4 output405 (.A(net405),
    .X(sram1_din0[18]));
 sky130_fd_sc_hd__buf_4 output406 (.A(net406),
    .X(sram1_din0[19]));
 sky130_fd_sc_hd__buf_4 output407 (.A(net407),
    .X(sram1_din0[1]));
 sky130_fd_sc_hd__buf_4 output408 (.A(net408),
    .X(sram1_din0[20]));
 sky130_fd_sc_hd__buf_4 output409 (.A(net409),
    .X(sram1_din0[21]));
 sky130_fd_sc_hd__buf_4 output410 (.A(net410),
    .X(sram1_din0[22]));
 sky130_fd_sc_hd__buf_4 output411 (.A(net411),
    .X(sram1_din0[23]));
 sky130_fd_sc_hd__buf_4 output412 (.A(net412),
    .X(sram1_din0[24]));
 sky130_fd_sc_hd__buf_4 output413 (.A(net413),
    .X(sram1_din0[25]));
 sky130_fd_sc_hd__buf_4 output414 (.A(net414),
    .X(sram1_din0[26]));
 sky130_fd_sc_hd__buf_4 output415 (.A(net415),
    .X(sram1_din0[27]));
 sky130_fd_sc_hd__buf_4 output416 (.A(net416),
    .X(sram1_din0[28]));
 sky130_fd_sc_hd__buf_4 output417 (.A(net417),
    .X(sram1_din0[29]));
 sky130_fd_sc_hd__buf_4 output418 (.A(net418),
    .X(sram1_din0[2]));
 sky130_fd_sc_hd__buf_4 output419 (.A(net419),
    .X(sram1_din0[30]));
 sky130_fd_sc_hd__buf_4 output420 (.A(net420),
    .X(sram1_din0[31]));
 sky130_fd_sc_hd__buf_4 output421 (.A(net421),
    .X(sram1_din0[3]));
 sky130_fd_sc_hd__buf_4 output422 (.A(net422),
    .X(sram1_din0[4]));
 sky130_fd_sc_hd__buf_4 output423 (.A(net423),
    .X(sram1_din0[5]));
 sky130_fd_sc_hd__buf_4 output424 (.A(net424),
    .X(sram1_din0[6]));
 sky130_fd_sc_hd__buf_4 output425 (.A(net425),
    .X(sram1_din0[7]));
 sky130_fd_sc_hd__buf_4 output426 (.A(net426),
    .X(sram1_din0[8]));
 sky130_fd_sc_hd__buf_4 output427 (.A(net427),
    .X(sram1_din0[9]));
 sky130_fd_sc_hd__buf_4 output428 (.A(net428),
    .X(sram1_web0));
 sky130_fd_sc_hd__buf_4 output429 (.A(net429),
    .X(sram1_wmask0[0]));
 sky130_fd_sc_hd__buf_4 output430 (.A(net430),
    .X(sram1_wmask0[1]));
 sky130_fd_sc_hd__buf_4 output431 (.A(net431),
    .X(sram1_wmask0[2]));
 sky130_fd_sc_hd__buf_4 output432 (.A(net432),
    .X(sram1_wmask0[3]));
 sky130_fd_sc_hd__buf_4 output433 (.A(net433),
    .X(vga_b[0]));
 sky130_fd_sc_hd__buf_4 output434 (.A(net434),
    .X(vga_b[1]));
 sky130_fd_sc_hd__buf_4 output435 (.A(net435),
    .X(vga_g[0]));
 sky130_fd_sc_hd__buf_4 output436 (.A(net436),
    .X(vga_g[1]));
 sky130_fd_sc_hd__buf_4 output437 (.A(net437),
    .X(vga_hsync));
 sky130_fd_sc_hd__buf_4 output438 (.A(net438),
    .X(vga_r[0]));
 sky130_fd_sc_hd__buf_4 output439 (.A(net439),
    .X(vga_r[1]));
 sky130_fd_sc_hd__buf_4 output440 (.A(net440),
    .X(vga_vsync));
 sky130_fd_sc_hd__buf_4 output441 (.A(net441),
    .X(video_irq[0]));
 sky130_fd_sc_hd__buf_4 output442 (.A(net442),
    .X(video_irq[1]));
 sky130_fd_sc_hd__buf_4 output443 (.A(net443),
    .X(wb_ack_o));
 sky130_fd_sc_hd__buf_4 output444 (.A(net444),
    .X(wb_data_o[0]));
 sky130_fd_sc_hd__buf_4 output445 (.A(net445),
    .X(wb_data_o[10]));
 sky130_fd_sc_hd__buf_4 output446 (.A(net446),
    .X(wb_data_o[11]));
 sky130_fd_sc_hd__buf_4 output447 (.A(net447),
    .X(wb_data_o[12]));
 sky130_fd_sc_hd__buf_4 output448 (.A(net448),
    .X(wb_data_o[13]));
 sky130_fd_sc_hd__buf_4 output449 (.A(net449),
    .X(wb_data_o[14]));
 sky130_fd_sc_hd__buf_4 output450 (.A(net450),
    .X(wb_data_o[15]));
 sky130_fd_sc_hd__buf_4 output451 (.A(net451),
    .X(wb_data_o[16]));
 sky130_fd_sc_hd__buf_4 output452 (.A(net452),
    .X(wb_data_o[17]));
 sky130_fd_sc_hd__buf_4 output453 (.A(net453),
    .X(wb_data_o[18]));
 sky130_fd_sc_hd__buf_4 output454 (.A(net454),
    .X(wb_data_o[19]));
 sky130_fd_sc_hd__buf_4 output455 (.A(net455),
    .X(wb_data_o[1]));
 sky130_fd_sc_hd__buf_4 output456 (.A(net456),
    .X(wb_data_o[20]));
 sky130_fd_sc_hd__buf_4 output457 (.A(net457),
    .X(wb_data_o[21]));
 sky130_fd_sc_hd__buf_4 output458 (.A(net458),
    .X(wb_data_o[22]));
 sky130_fd_sc_hd__buf_4 output459 (.A(net459),
    .X(wb_data_o[23]));
 sky130_fd_sc_hd__buf_4 output460 (.A(net460),
    .X(wb_data_o[24]));
 sky130_fd_sc_hd__buf_4 output461 (.A(net461),
    .X(wb_data_o[25]));
 sky130_fd_sc_hd__buf_4 output462 (.A(net462),
    .X(wb_data_o[26]));
 sky130_fd_sc_hd__buf_4 output463 (.A(net463),
    .X(wb_data_o[27]));
 sky130_fd_sc_hd__buf_4 output464 (.A(net464),
    .X(wb_data_o[28]));
 sky130_fd_sc_hd__buf_4 output465 (.A(net465),
    .X(wb_data_o[29]));
 sky130_fd_sc_hd__buf_4 output466 (.A(net466),
    .X(wb_data_o[2]));
 sky130_fd_sc_hd__buf_4 output467 (.A(net467),
    .X(wb_data_o[30]));
 sky130_fd_sc_hd__buf_4 output468 (.A(net468),
    .X(wb_data_o[31]));
 sky130_fd_sc_hd__buf_4 output469 (.A(net469),
    .X(wb_data_o[3]));
 sky130_fd_sc_hd__buf_4 output470 (.A(net470),
    .X(wb_data_o[4]));
 sky130_fd_sc_hd__buf_4 output471 (.A(net471),
    .X(wb_data_o[5]));
 sky130_fd_sc_hd__buf_4 output472 (.A(net472),
    .X(wb_data_o[6]));
 sky130_fd_sc_hd__buf_4 output473 (.A(net473),
    .X(wb_data_o[7]));
 sky130_fd_sc_hd__buf_4 output474 (.A(net474),
    .X(wb_data_o[8]));
 sky130_fd_sc_hd__buf_4 output475 (.A(net475),
    .X(wb_data_o[9]));
 sky130_fd_sc_hd__buf_4 output476 (.A(net476),
    .X(wb_stall_o));
 assign wb_error_o = net619;
endmodule

