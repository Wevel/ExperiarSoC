* NGSPICE file created from PWM.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

.subckt PWM clk peripheralBus_address[0] peripheralBus_address[10] peripheralBus_address[11]
+ peripheralBus_address[12] peripheralBus_address[13] peripheralBus_address[14] peripheralBus_address[15]
+ peripheralBus_address[16] peripheralBus_address[17] peripheralBus_address[18] peripheralBus_address[19]
+ peripheralBus_address[1] peripheralBus_address[20] peripheralBus_address[21] peripheralBus_address[22]
+ peripheralBus_address[23] peripheralBus_address[2] peripheralBus_address[3] peripheralBus_address[4]
+ peripheralBus_address[5] peripheralBus_address[6] peripheralBus_address[7] peripheralBus_address[8]
+ peripheralBus_address[9] peripheralBus_busy peripheralBus_data[0] peripheralBus_data[10]
+ peripheralBus_data[11] peripheralBus_data[12] peripheralBus_data[13] peripheralBus_data[14]
+ peripheralBus_data[15] peripheralBus_data[16] peripheralBus_data[17] peripheralBus_data[18]
+ peripheralBus_data[19] peripheralBus_data[1] peripheralBus_data[20] peripheralBus_data[21]
+ peripheralBus_data[22] peripheralBus_data[23] peripheralBus_data[24] peripheralBus_data[25]
+ peripheralBus_data[26] peripheralBus_data[27] peripheralBus_data[28] peripheralBus_data[29]
+ peripheralBus_data[2] peripheralBus_data[30] peripheralBus_data[31] peripheralBus_data[3]
+ peripheralBus_data[4] peripheralBus_data[5] peripheralBus_data[6] peripheralBus_data[7]
+ peripheralBus_data[8] peripheralBus_data[9] peripheralBus_oe peripheralBus_we pwm_en[0]
+ pwm_en[10] pwm_en[11] pwm_en[12] pwm_en[13] pwm_en[14] pwm_en[15] pwm_en[1] pwm_en[2]
+ pwm_en[3] pwm_en[4] pwm_en[5] pwm_en[6] pwm_en[7] pwm_en[8] pwm_en[9] pwm_out[0]
+ pwm_out[10] pwm_out[11] pwm_out[12] pwm_out[13] pwm_out[14] pwm_out[15] pwm_out[1]
+ pwm_out[2] pwm_out[3] pwm_out[4] pwm_out[5] pwm_out[6] pwm_out[7] pwm_out[8] pwm_out[9]
+ rst vccd1 vssd1
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10669__A1 _10665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ _09671_/A vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06883_ _06883_/A vssd1 vssd1 vccd1 vccd1 _06883_/X sky130_fd_sc_hd__clkbuf_1
X_13206__362 vssd1 vssd1 vccd1 vccd1 _13206__362/HI _13829_/A sky130_fd_sc_hd__conb_1
XFILLER_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08622_ _09397_/C vssd1 vssd1 vccd1 vccd1 _13553_/A sky130_fd_sc_hd__buf_4
XFILLER_55_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08553_ _13584_/A vssd1 vssd1 vccd1 vccd1 _08553_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07504_ _07504_/A _07504_/B _07510_/C vssd1 vssd1 vccd1 vccd1 _07505_/A sky130_fd_sc_hd__or3_1
X_08484_ _08480_/X _08483_/X _08498_/S vssd1 vssd1 vccd1 vccd1 _11705_/C sky130_fd_sc_hd__mux2_1
XFILLER_50_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07435_ _07442_/A _07435_/B vssd1 vssd1 vccd1 vccd1 _07436_/A sky130_fd_sc_hd__or2_1
XFILLER_23_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07366_ _07393_/A vssd1 vssd1 vccd1 vccd1 _07377_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10693__B _11412_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09105_ input27/X vssd1 vssd1 vccd1 vccd1 _11503_/B sky130_fd_sc_hd__inv_6
X_06317_ _06317_/A vssd1 vssd1 vccd1 vccd1 _06317_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07297_ _07297_/A vssd1 vssd1 vccd1 vccd1 _07297_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09036_ _11677_/B _11677_/A _11676_/B _11676_/A _08941_/X _08942_/X vssd1 vssd1 vccd1
+ vccd1 _09036_/X sky130_fd_sc_hd__mux4_2
XFILLER_163_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09938_ _14035_/Z _08695_/X _09953_/S vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10109__B1 _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08948__S1 _08947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ _09869_/A _09869_/B _09869_/C vssd1 vssd1 vccd1 vccd1 _09869_/Y sky130_fd_sc_hd__nor3_1
XFILLER_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11900_ _11900_/A vssd1 vssd1 vccd1 vccd1 _12902_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09722__B _13557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12880_ _12904_/CLK _12880_/D vssd1 vssd1 vccd1 vccd1 _14008_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11831_ _11834_/A _11831_/B vssd1 vssd1 vccd1 vccd1 _11832_/A sky130_fd_sc_hd__and2_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11762_/A vssd1 vssd1 vccd1 vccd1 _12868_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13501_/A _07620_/X vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__ebufn_8
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _13973_/Z _13781_/A _10723_/S vssd1 vssd1 vccd1 vccd1 _10714_/B sky130_fd_sc_hd__mux2_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11695_/B _11695_/C _11569_/X vssd1 vssd1 vccd1 vccd1 _11694_/B sky130_fd_sc_hd__o21ai_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13432_ _13432_/A _07800_/X vssd1 vssd1 vccd1 vccd1 _14104_/Z sky130_fd_sc_hd__ebufn_8
X_10644_ _10385_/X _10638_/X _10643_/X _10550_/X vssd1 vssd1 vccd1 vccd1 _12585_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08354__A _08358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13363_ _13363_/A _08286_/X vssd1 vssd1 vccd1 vccd1 _14067_/Z sky130_fd_sc_hd__ebufn_8
X_10575_ _13716_/A _12572_/Q _10584_/S vssd1 vssd1 vccd1 vccd1 _10576_/B sky130_fd_sc_hd__mux2_1
XFILLER_158_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12314_ _12320_/CLK _12314_/D vssd1 vssd1 vccd1 vccd1 _12314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13149__305 vssd1 vssd1 vccd1 vccd1 _13149__305/HI _13706_/A sky130_fd_sc_hd__conb_1
XFILLER_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09202__A1 _09379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ _12251_/CLK _12245_/D vssd1 vssd1 vccd1 vccd1 _12245_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_repeater127_A _13979_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09185__A _13626_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ _12176_/A _12176_/B _12176_/C _12176_/D vssd1 vssd1 vccd1 vccd1 _12177_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_69_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ _12703_/Q _13944_/A vssd1 vssd1 vccd1 vccd1 _11127_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11058_ _10408_/X _11055_/X _11057_/X _11053_/X vssd1 vssd1 vccd1 vccd1 _12688_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_output56_A _13569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09061__S0 _08941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ _10077_/A vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08248__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07220_ _07220_/A _07231_/B _07228_/C vssd1 vssd1 vccd1 vccd1 _07221_/A sky130_fd_sc_hd__or3_1
Xrepeater60 _14072_/Z vssd1 vssd1 vccd1 vccd1 _13976_/Z sky130_fd_sc_hd__buf_12
Xrepeater71 peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 _14037_/Z sky130_fd_sc_hd__buf_12
Xrepeater82 peripheralBus_data[31] vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__buf_12
XFILLER_158_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater93 peripheralBus_data[27] vssd1 vssd1 vccd1 vccd1 _13994_/Z sky130_fd_sc_hd__buf_12
XFILLER_164_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07151_ _07205_/A vssd1 vssd1 vccd1 vccd1 _07163_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__11402__B _13935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07082_ _07533_/A vssd1 vssd1 vccd1 vccd1 _07137_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07984_ _07984_/A vssd1 vssd1 vccd1 vccd1 _07984_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09723_ _12344_/Q _13554_/A vssd1 vssd1 vccd1 vccd1 _09725_/C sky130_fd_sc_hd__xor2_1
X_06935_ _06935_/A vssd1 vssd1 vccd1 vccd1 _06935_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09052__S0 _08911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09654_ _13469_/A _09640_/X _09653_/X _09649_/X vssd1 vssd1 vccd1 vccd1 _12339_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06866_ _06877_/A _06870_/B _06870_/C vssd1 vssd1 vccd1 vccd1 _06867_/A sky130_fd_sc_hd__or3_1
XANTENNA__10688__B _11924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08605_ _12427_/Q vssd1 vssd1 vccd1 vccd1 _09997_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06797_ _06801_/A _06806_/B _06806_/C vssd1 vssd1 vccd1 vccd1 _06798_/A sky130_fd_sc_hd__or3_1
X_09585_ _11443_/A vssd1 vssd1 vccd1 vccd1 _12200_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08536_ _08423_/X _08428_/X _08427_/X _08430_/X _08470_/X _09152_/A vssd1 vssd1 vccd1
+ vccd1 _08536_/X sky130_fd_sc_hd__mux4_1
X_08467_ _08479_/A vssd1 vssd1 vccd1 vccd1 _08467_/X sky130_fd_sc_hd__buf_2
XFILLER_11_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07418_ _07418_/A vssd1 vssd1 vccd1 vccd1 _07418_/X sky130_fd_sc_hd__clkbuf_1
X_08398_ _12233_/Q _12234_/Q _12235_/Q _12236_/Q _08396_/X _08397_/X vssd1 vssd1 vccd1
+ vccd1 _08398_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_93_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13334__490 vssd1 vssd1 vccd1 vccd1 _13334__490/HI _14087_/A sky130_fd_sc_hd__conb_1
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07349_ _09875_/B vssd1 vssd1 vccd1 vccd1 _07403_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08866__S0 _08733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06406__B _06412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10360_ _12504_/Q _13746_/A vssd1 vssd1 vccd1 vccd1 _10362_/C sky130_fd_sc_hd__xor2_1
XFILLER_136_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ _08948_/X _08951_/X _08950_/X _08955_/X _09057_/A _09013_/X vssd1 vssd1 vccd1
+ vccd1 _09019_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09717__B _13552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10291_ _13629_/A _10291_/B vssd1 vssd1 vccd1 vccd1 _10291_/X sky130_fd_sc_hd__or2_1
XFILLER_136_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12030_ _12030_/A _12030_/B vssd1 vssd1 vccd1 vccd1 _12031_/A sky130_fd_sc_hd__and2_1
XFILLER_105_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10750__B1 _10749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_clk_A _12759_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13981_ _13981_/A _06337_/X vssd1 vssd1 vccd1 vccd1 _14077_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_74_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12932_ _12952_/CLK _12932_/D vssd1 vssd1 vccd1 vccd1 _12932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _12867_/CLK _12863_/D vssd1 vssd1 vccd1 vccd1 _12863_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11058__A1 _10408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _11814_/A vssd1 vssd1 vccd1 vccd1 _12877_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12799_/CLK _12794_/D vssd1 vssd1 vccd1 vccd1 _13968_/A sky130_fd_sc_hd__dfxtp_2
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11745_/A vssd1 vssd1 vccd1 vccd1 _12863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11503__A _11680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11676_ _11676_/A _11676_/B _11676_/C vssd1 vssd1 vccd1 vccd1 _11677_/C sky130_fd_sc_hd__and3_1
XANTENNA__08084__A _08084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13415_ _13415_/A _08165_/X vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__ebufn_8
X_10627_ _10627_/A _10627_/B _10627_/C _10627_/D vssd1 vssd1 vccd1 vccd1 _10633_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_104_clk_A _12217_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10558_ _10567_/A _10558_/B vssd1 vssd1 vccd1 vccd1 _10559_/A sky130_fd_sc_hd__and2_1
XFILLER_5_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10489_ _10484_/Y _10485_/X _10486_/X _10487_/Y _10488_/Y vssd1 vssd1 vccd1 vccd1
+ _10489_/X sky130_fd_sc_hd__o221a_1
X_12228_ _12295_/CLK _12228_/D vssd1 vssd1 vccd1 vccd1 _12228_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12053__B _13363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12159_ _12966_/Q _13372_/A vssd1 vssd1 vccd1 vccd1 _12161_/C sky130_fd_sc_hd__xor2_1
XFILLER_123_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06720_ _06720_/A vssd1 vssd1 vccd1 vccd1 _06720_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06651_ _06659_/A _06651_/B _06651_/C vssd1 vssd1 vccd1 vccd1 _06652_/A sky130_fd_sc_hd__or3_1
X_13277__433 vssd1 vssd1 vccd1 vccd1 _13277__433/HI _13982_/A sky130_fd_sc_hd__conb_1
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09370_ _09370_/A _09377_/C _09382_/B vssd1 vssd1 vccd1 vccd1 _09370_/X sky130_fd_sc_hd__and3_1
XFILLER_24_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06582_ _06584_/A _06589_/B _06589_/C vssd1 vssd1 vccd1 vccd1 _06583_/A sky130_fd_sc_hd__or3_1
XFILLER_33_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08321_ _08324_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__or2_1
X_13318__474 vssd1 vssd1 vccd1 vccd1 _13318__474/HI _14055_/A sky130_fd_sc_hd__conb_1
XFILLER_33_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08252_ _08252_/A vssd1 vssd1 vccd1 vccd1 _08252_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07203_ _07206_/A _07203_/B _07213_/C vssd1 vssd1 vccd1 vccd1 _07204_/A sky130_fd_sc_hd__or3_1
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12991__147 vssd1 vssd1 vccd1 vccd1 _12991__147/HI _13388_/A sky130_fd_sc_hd__conb_1
XANTENNA__11132__B _13946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ _08183_/A vssd1 vssd1 vccd1 vccd1 _08183_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_12_0_clk/X
+ sky130_fd_sc_hd__clkbuf_2
X_07134_ _07615_/A vssd1 vssd1 vccd1 vccd1 _07145_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_145_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07065_ _07120_/A vssd1 vssd1 vccd1 vccd1 _07076_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07338__A _07406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07057__B _07979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07967_ _08075_/A _08075_/B _07977_/C vssd1 vssd1 vccd1 vccd1 _07968_/A sky130_fd_sc_hd__or3_1
XFILLER_102_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11288__A1 _11153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _09706_/A vssd1 vssd1 vccd1 vccd1 _12354_/D sky130_fd_sc_hd__clkbuf_1
X_06918_ _06955_/A vssd1 vssd1 vccd1 vccd1 _06929_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07898_ _07898_/A vssd1 vssd1 vccd1 vccd1 _07898_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09637_ _13463_/A _09627_/X _09636_/X _09634_/X vssd1 vssd1 vccd1 vccd1 _12333_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06849_ _06849_/A vssd1 vssd1 vccd1 vccd1 _06849_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11026__C _11410_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _09568_/A vssd1 vssd1 vccd1 vccd1 _12318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08519_ _13396_/A vssd1 vssd1 vccd1 vccd1 _09162_/A sky130_fd_sc_hd__buf_2
XFILLER_24_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09499_ _13427_/A _09483_/X _09498_/X _09496_/X vssd1 vssd1 vccd1 vccd1 _12296_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10799__B1 _10798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11530_ _11530_/A _11530_/B vssd1 vssd1 vccd1 vccd1 _12812_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13070__226 vssd1 vssd1 vccd1 vccd1 _13070__226/HI _13545_/A sky130_fd_sc_hd__conb_1
X_11461_ _11474_/A vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__clkbuf_2
X_10412_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10412_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11392_ _12774_/Q _13949_/A vssd1 vssd1 vccd1 vccd1 _11395_/B sky130_fd_sc_hd__xor2_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10343_ _10349_/A _10343_/B vssd1 vssd1 vccd1 vccd1 _10344_/A sky130_fd_sc_hd__and2_1
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13111__267 vssd1 vssd1 vccd1 vccd1 _13111__267/HI _13636_/A sky130_fd_sc_hd__conb_1
XANTENNA__07248__A _07248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10274_ _13623_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10274_/X sky130_fd_sc_hd__or2_1
XFILLER_140_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12013_ _12013_/A _12013_/B vssd1 vssd1 vccd1 vccd1 _12014_/A sky130_fd_sc_hd__and2_1
XFILLER_105_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10723__A0 _13976_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13964_ _13964_/A _06386_/X vssd1 vssd1 vccd1 vccd1 _14028_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12915_ _12918_/CLK _12915_/D vssd1 vssd1 vccd1 vccd1 _14042_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13895_ _13895_/A _06570_/X vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__ebufn_8
X_13005__161 vssd1 vssd1 vccd1 vccd1 _13005__161/HI _13416_/A sky130_fd_sc_hd__conb_1
X_12846_ _12850_/CLK _12846_/D vssd1 vssd1 vccd1 vccd1 _12846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ _12782_/CLK _12777_/D vssd1 vssd1 vccd1 vccd1 _13903_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ _11728_/A vssd1 vssd1 vccd1 vccd1 _12858_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11451__A1 _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12048__B _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11659_ _11659_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _12841_/D sky130_fd_sc_hd__nor2_1
XFILLER_128_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09638__A _09638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08870_ _08783_/X _08787_/X _08790_/X _08791_/X _08826_/X _08859_/X vssd1 vssd1 vccd1
+ vccd1 _08870_/X sky130_fd_sc_hd__mux4_1
XANTENNA__06997__A _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07821_ _07821_/A vssd1 vssd1 vccd1 vccd1 _07821_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11408__A _11408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ _07752_/A vssd1 vssd1 vccd1 vccd1 _07752_/X sky130_fd_sc_hd__clkbuf_1
X_06703_ _06748_/A vssd1 vssd1 vccd1 vccd1 _06714_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__11127__B _13944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ _07686_/A _07683_/B _07691_/C vssd1 vssd1 vccd1 vccd1 _07684_/A sky130_fd_sc_hd__or3_1
XANTENNA__09883__A1 _09750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ _09422_/A _09422_/B vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__and2_1
X_06634_ _06646_/A _06651_/B _07995_/B vssd1 vssd1 vccd1 vccd1 _06635_/A sky130_fd_sc_hd__or3_1
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ _09353_/A _09355_/B vssd1 vssd1 vccd1 vccd1 _12263_/D sky130_fd_sc_hd__nor2_1
X_06565_ _06569_/A _06574_/B _06574_/C vssd1 vssd1 vccd1 vccd1 _06566_/A sky130_fd_sc_hd__or3_1
X_08304_ _08304_/A vssd1 vssd1 vccd1 vccd1 _08304_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09284_ _09322_/A _09322_/B _09321_/C _09284_/D vssd1 vssd1 vccd1 vccd1 _09331_/A
+ sky130_fd_sc_hd__and4_1
X_06496_ _06523_/A vssd1 vssd1 vccd1 vccd1 _06507_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08235_ _08238_/A _08235_/B _08238_/C vssd1 vssd1 vccd1 vccd1 _08236_/A sky130_fd_sc_hd__or3_1
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08166_ _08166_/A vssd1 vssd1 vccd1 vccd1 _08364_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_07117_ _07162_/A vssd1 vssd1 vccd1 vccd1 _07128_/C sky130_fd_sc_hd__clkbuf_1
X_08097_ _08101_/A _08101_/B _08105_/C vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__or3_1
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07068__A _08177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07048_ _07048_/A vssd1 vssd1 vccd1 vccd1 _07048_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08999_ _11631_/C _12827_/Q _11632_/A _11641_/D _08911_/X _08913_/X vssd1 vssd1 vccd1
+ vccd1 _08999_/X sky130_fd_sc_hd__mux4_2
XFILLER_29_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10961_ _10961_/A vssd1 vssd1 vccd1 vccd1 _12665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12700_ _12704_/CLK _12700_/D vssd1 vssd1 vccd1 vccd1 _12700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11681__A1 _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ _13680_/A _07146_/X vssd1 vssd1 vccd1 vccd1 _14096_/Z sky130_fd_sc_hd__ebufn_8
X_10892_ _10897_/C _10897_/D _10891_/Y _10749_/X vssd1 vssd1 vccd1 vccd1 _12647_/D
+ sky130_fd_sc_hd__o211a_1
X_12631_ _12634_/CLK _12631_/D vssd1 vssd1 vccd1 vccd1 _12631_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11053__A _11195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11433__A1 _10662_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12562_ _12565_/CLK _12562_/D vssd1 vssd1 vccd1 vccd1 _13690_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11513_ _11513_/A vssd1 vssd1 vccd1 vccd1 _12808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12493_ _12522_/CLK _12493_/D vssd1 vssd1 vccd1 vccd1 _13623_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11444_ _12084_/A vssd1 vssd1 vccd1 vccd1 _11444_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08362__A _08364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11375_ _11375_/A vssd1 vssd1 vccd1 vccd1 _12773_/D sky130_fd_sc_hd__clkbuf_1
X_10326_ _10326_/A vssd1 vssd1 vccd1 vccd1 _12509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14094_ _14094_/A _08157_/X vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__ebufn_8
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _09139_/X _10249_/X _10255_/X _10256_/X vssd1 vssd1 vccd1 vccd1 _12486_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07706__A _09484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ _10191_/A _10188_/B vssd1 vssd1 vccd1 vccd1 _10189_/A sky130_fd_sc_hd__and2_1
X_13947_ _13947_/A _06429_/X vssd1 vssd1 vccd1 vccd1 _13979_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_35_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ _13878_/A _06617_/X vssd1 vssd1 vccd1 vccd1 _14070_/Z sky130_fd_sc_hd__ebufn_8
X_12829_ _12829_/CLK _12829_/D vssd1 vssd1 vccd1 vccd1 _12829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09617__A1 _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06350_ _06350_/A vssd1 vssd1 vccd1 vccd1 _06350_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11424__A1 _10652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06281_ input26/X input25/X vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__or2b_2
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08020_ _08025_/A _08020_/B _08030_/C vssd1 vssd1 vccd1 vccd1 _08021_/A sky130_fd_sc_hd__or3_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11410__B _11412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09971_ _09971_/A vssd1 vssd1 vccd1 vccd1 _12421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ _13969_/A vssd1 vssd1 vccd1 vccd1 _08922_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater89_A peripheralBus_data[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ _12651_/Q vssd1 vssd1 vccd1 vccd1 _10907_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07804_ _07809_/A _07806_/B _07815_/C vssd1 vssd1 vccd1 vccd1 _07805_/A sky130_fd_sc_hd__or3_1
X_08784_ _12629_/Q vssd1 vssd1 vccd1 vccd1 _10864_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07735_ _07742_/A _07737_/B _07748_/C vssd1 vssd1 vccd1 vccd1 _07736_/A sky130_fd_sc_hd__or3_1
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07666_ _07693_/A vssd1 vssd1 vccd1 vccd1 _07678_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07989__C _07993_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09405_ _09405_/A vssd1 vssd1 vccd1 vccd1 _12275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06617_ _06617_/A vssd1 vssd1 vccd1 vccd1 _06617_/X sky130_fd_sc_hd__clkbuf_1
X_12997__153 vssd1 vssd1 vccd1 vccd1 _12997__153/HI _13408_/A sky130_fd_sc_hd__conb_1
X_07597_ _07597_/A vssd1 vssd1 vccd1 vccd1 _07597_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11415__A1 _11153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ _09336_/A _09336_/B _09336_/C vssd1 vssd1 vccd1 vccd1 _09343_/D sky130_fd_sc_hd__and3_1
X_06548_ _06548_/A _12059_/A _06548_/C _09096_/C vssd1 vssd1 vccd1 vccd1 _06577_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_139_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09267_ _09328_/C _09332_/B _09266_/Y vssd1 vssd1 vccd1 vccd1 _12244_/D sky130_fd_sc_hd__a21oi_1
XFILLER_139_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06479_ _06481_/A _06486_/B _06486_/C vssd1 vssd1 vccd1 vccd1 _06480_/A sky130_fd_sc_hd__or3_1
XFILLER_138_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ _08225_/A _08222_/B _08225_/C vssd1 vssd1 vccd1 vccd1 _08219_/A sky130_fd_sc_hd__or3_1
XFILLER_126_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09198_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09380_/A sky130_fd_sc_hd__buf_2
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08149_ _08149_/A vssd1 vssd1 vccd1 vccd1 _08149_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10926__B1 _10798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11160_ _11160_/A vssd1 vssd1 vccd1 vccd1 _11160_/X sky130_fd_sc_hd__buf_4
XANTENNA__08690__S1 _08603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10111_ _10111_/A _10111_/B _10111_/C vssd1 vssd1 vccd1 vccd1 _10133_/C sky130_fd_sc_hd__and3_1
XFILLER_106_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11091_ _13844_/A _12699_/Q _11101_/S vssd1 vssd1 vccd1 vccd1 _11092_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13182__338 vssd1 vssd1 vccd1 vccd1 _13182__338/HI _13789_/A sky130_fd_sc_hd__conb_1
XFILLER_96_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07526__A _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ _12439_/Q vssd1 vssd1 vccd1 vccd1 _10052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06430__A _06442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13223__379 vssd1 vssd1 vccd1 vccd1 _13223__379/HI _13862_/A sky130_fd_sc_hd__conb_1
XANTENNA__09741__A _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13801_ _13801_/A _06835_/X vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input18_A peripheralBus_address[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11993_ _11996_/A _11993_/B vssd1 vssd1 vccd1 vccd1 _11994_/A sky130_fd_sc_hd__and2_1
XANTENNA__09460__B _13555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13732_ _13732_/A _07012_/X vssd1 vssd1 vccd1 vccd1 _13988_/Z sky130_fd_sc_hd__ebufn_8
X_10944_ _10996_/S vssd1 vssd1 vccd1 vccd1 _10955_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13663_ _13663_/A _07191_/X vssd1 vssd1 vccd1 vccd1 _14079_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_32_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10875_ _10875_/A _10875_/B _10875_/C vssd1 vssd1 vccd1 vccd1 _10877_/C sky130_fd_sc_hd__and3_1
X_13076__232 vssd1 vssd1 vccd1 vccd1 _13076__232/HI _13571_/A sky130_fd_sc_hd__conb_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12614_ _12660_/CLK _12614_/D vssd1 vssd1 vccd1 vccd1 _12614_/Q sky130_fd_sc_hd__dfxtp_1
X_13594_ _13594_/A _07381_/X vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_12_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12545_ _12565_/CLK _12545_/D vssd1 vssd1 vccd1 vccd1 _12545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09480__C1 _09192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14094__A _14094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13117__273 vssd1 vssd1 vccd1 vccd1 _13117__273/HI _13642_/A sky130_fd_sc_hd__conb_1
XFILLER_129_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12476_ _12656_/CLK _12476_/D vssd1 vssd1 vccd1 vccd1 _12476_/Q sky130_fd_sc_hd__dfxtp_1
X_11427_ _13908_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11427_/X sky130_fd_sc_hd__or2_1
XANTENNA__10127__A _10146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11358_ _11358_/A vssd1 vssd1 vccd1 vccd1 _12768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10393__A1 _09756_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ _10309_/A vssd1 vssd1 vccd1 vccd1 _12504_/D sky130_fd_sc_hd__clkbuf_1
X_14077_ _14077_/A _08031_/X vssd1 vssd1 vccd1 vccd1 _14077_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11289_ _13872_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11289_/X sky130_fd_sc_hd__or2_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09651__A _11064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07520_ _08210_/A vssd1 vssd1 vccd1 vccd1 _08197_/A sky130_fd_sc_hd__buf_4
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08267__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07451_ _07451_/A vssd1 vssd1 vccd1 vccd1 _07451_/X sky130_fd_sc_hd__clkbuf_2
X_06402_ _07845_/B vssd1 vssd1 vccd1 vccd1 _06412_/B sky130_fd_sc_hd__clkbuf_4
X_07382_ _07382_/A _07391_/B _07388_/C vssd1 vssd1 vccd1 vccd1 _07383_/A sky130_fd_sc_hd__or3_1
XFILLER_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ _14110_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _09121_/X sky130_fd_sc_hd__or2_1
X_06333_ _06333_/A _06336_/B _06336_/C vssd1 vssd1 vccd1 vccd1 _06334_/A sky130_fd_sc_hd__or3_1
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09052_ _11676_/A _11688_/A _12847_/Q _12848_/Q _08911_/X _08913_/X vssd1 vssd1 vccd1
+ vccd1 _09052_/X sky130_fd_sc_hd__mux4_1
X_06264_ input19/X _09096_/B vssd1 vssd1 vccd1 vccd1 _06548_/C sky130_fd_sc_hd__or2_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06515__A _08210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08003_ _08003_/A vssd1 vssd1 vccd1 vccd1 _08003_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11140__B _13950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10384__A1 _10377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09954_ _10700_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _09955_/A sky130_fd_sc_hd__or2_1
XANTENNA__13615__TE_B _07994_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08905_ _10928_/B _12658_/Q _12659_/Q _12660_/Q _10697_/A _08887_/X vssd1 vssd1 vccd1
+ vccd1 _08905_/X sky130_fd_sc_hd__mux4_2
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _09753_/X _09874_/X _09884_/X _09878_/X vssd1 vssd1 vccd1 vccd1 _12394_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08836_ _10162_/A vssd1 vssd1 vccd1 vccd1 _13747_/A sky130_fd_sc_hd__buf_6
XANTENNA__09561__A _09582_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08767_ _13777_/A vssd1 vssd1 vccd1 vccd1 _08767_/X sky130_fd_sc_hd__buf_2
XFILLER_122_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ _07718_/A vssd1 vssd1 vccd1 vccd1 _07718_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _12461_/Q vssd1 vssd1 vccd1 vccd1 _10148_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08177__A _08177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07081__A _07603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07649_ _07659_/A _07654_/B _07649_/C vssd1 vssd1 vccd1 vccd1 _07650_/A sky130_fd_sc_hd__or3_1
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13811__A _13811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ _13717_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10660_/X sky130_fd_sc_hd__or2_1
XFILLER_15_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09319_ _09329_/B _09329_/C vssd1 vssd1 vccd1 vccd1 _09323_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_114_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _12295_/CLK sky130_fd_sc_hd__clkbuf_16
X_10591_ _10591_/A vssd1 vssd1 vccd1 vccd1 _12576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12330_ _12331_/CLK _12330_/D vssd1 vssd1 vccd1 vccd1 _13460_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12261_ _12264_/CLK _12261_/D vssd1 vssd1 vccd1 vccd1 _12261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14000_ _14000_/A _07984_/X vssd1 vssd1 vccd1 vccd1 _14096_/Z sky130_fd_sc_hd__ebufn_8
X_11212_ _11212_/A vssd1 vssd1 vccd1 vccd1 _12729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12192_ _10652_/A _12182_/X _12191_/X _12187_/X vssd1 vssd1 vccd1 vccd1 _12974_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput31 _13977_/A vssd1 vssd1 vccd1 vccd1 pwm_en[12] sky130_fd_sc_hd__buf_2
XFILLER_134_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput42 _13785_/A vssd1 vssd1 vccd1 vccd1 pwm_en[8] sky130_fd_sc_hd__buf_2
X_11143_ _11143_/A _11143_/B _11143_/C _11143_/D vssd1 vssd1 vccd1 vccd1 _11149_/B
+ sky130_fd_sc_hd__or4_1
Xoutput53 _13378_/A vssd1 vssd1 vccd1 vccd1 pwm_out[3] sky130_fd_sc_hd__buf_2
XFILLER_122_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11074_ _13839_/A _12694_/Q _11151_/B vssd1 vssd1 vccd1 vccd1 _11075_/B sky130_fd_sc_hd__mux2_1
X_10025_ _10022_/A _10030_/C _10029_/B vssd1 vssd1 vccd1 vccd1 _10026_/C sky130_fd_sc_hd__a21o_1
XFILLER_49_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11976_ _11976_/A vssd1 vssd1 vccd1 vccd1 _12918_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10410__A _10423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13715_ _13715_/A _07052_/X vssd1 vssd1 vccd1 vccd1 _14099_/Z sky130_fd_sc_hd__ebufn_8
X_10927_ _10927_/A _10927_/B vssd1 vssd1 vccd1 vccd1 _12657_/D sky130_fd_sc_hd__nor2_1
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13646_ _13646_/A _07235_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_158_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10858_ _10875_/A _10859_/B vssd1 vssd1 vccd1 vccd1 _10860_/B sky130_fd_sc_hd__or2_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_105_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _12969_/CLK sky130_fd_sc_hd__clkbuf_16
X_13577_ _13577_/A _07427_/X vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10789_ _12625_/Q vssd1 vssd1 vccd1 vccd1 _10865_/A sky130_fd_sc_hd__clkbuf_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11241__A _11363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12528_ _12583_/CLK _12528_/D vssd1 vssd1 vccd1 vccd1 _13657_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ _12461_/CLK _12459_/D vssd1 vssd1 vccd1 vccd1 _12459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09646__A _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__S1 _08557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06951_ _06960_/A _06953_/B vssd1 vssd1 vccd1 vccd1 _06952_/A sky130_fd_sc_hd__or2_1
XFILLER_113_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09670_ _09670_/A vssd1 vssd1 vccd1 vccd1 _12344_/D sky130_fd_sc_hd__clkbuf_1
X_06882_ _06890_/A _06884_/B _06884_/C vssd1 vssd1 vccd1 vccd1 _06883_/A sky130_fd_sc_hd__or3_1
XFILLER_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08621_ _08613_/X _08620_/X _08682_/S vssd1 vssd1 vccd1 vccd1 _09397_/C sky130_fd_sc_hd__mux2_1
XFILLER_82_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08552_ _12421_/Q _12422_/Q _12423_/Q _09981_/A _08549_/X _08551_/X vssd1 vssd1 vccd1
+ vccd1 _08552_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07503_ _07503_/A vssd1 vssd1 vccd1 vccd1 _07503_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11135__B _13949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ _08428_/X _08431_/X _08430_/X _08482_/X _08517_/A _08467_/X vssd1 vssd1 vccd1
+ vccd1 _08483_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07434_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07434_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07365_ _07365_/A vssd1 vssd1 vccd1 vccd1 _07365_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11151__A _11151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ _14107_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _09104_/X sky130_fd_sc_hd__or2_1
XANTENNA__10693__C _10693_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09995__B1 _09994_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06316_ _06320_/A _06323_/B _06323_/C vssd1 vssd1 vccd1 vccd1 _06317_/A sky130_fd_sc_hd__or3_1
X_07296_ _07307_/A _07303_/B _07300_/C vssd1 vssd1 vccd1 vccd1 _07297_/A sky130_fd_sc_hd__or3_1
X_09035_ _12845_/Q vssd1 vssd1 vccd1 vccd1 _11676_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09937_ _09937_/A vssd1 vssd1 vccd1 vccd1 _09953_/S sky130_fd_sc_hd__buf_2
XFILLER_131_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _09868_/A _09868_/B _09868_/C _09868_/D vssd1 vssd1 vccd1 vccd1 _09869_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_58_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08819_ _12641_/Q vssd1 vssd1 vccd1 vccd1 _10876_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09799_ _13521_/A _12376_/Q _09871_/B vssd1 vssd1 vccd1 vccd1 _09800_/B sky130_fd_sc_hd__mux2_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ peripheralBus_data[11] _14010_/A _11840_/S vssd1 vssd1 vccd1 vccd1 _11831_/B
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11799_/A _11761_/B vssd1 vssd1 vccd1 vccd1 _11762_/A sky130_fd_sc_hd__and2_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13500_/A _07622_/X vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_8
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10394_/X _10690_/X _10710_/X _10711_/X vssd1 vssd1 vccd1 vccd1 _12605_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11695_/B _11695_/C vssd1 vssd1 vccd1 vccd1 _11694_/A sky130_fd_sc_hd__and2_1
XFILLER_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _13431_/A _07802_/X vssd1 vssd1 vccd1 vccd1 _13623_/Z sky130_fd_sc_hd__ebufn_8
X_10643_ _13712_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10643_/X sky130_fd_sc_hd__or2_1
XFILLER_139_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08354__B _08358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__A _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ _13362_/A _08284_/X vssd1 vssd1 vccd1 vccd1 _14098_/Z sky130_fd_sc_hd__ebufn_8
X_10574_ _10574_/A vssd1 vssd1 vccd1 vccd1 _12571_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_5_clk_A _12917_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12313_ _12313_/CLK _12313_/D vssd1 vssd1 vccd1 vccd1 _12313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13188__344 vssd1 vssd1 vccd1 vccd1 _13188__344/HI _13795_/A sky130_fd_sc_hd__conb_1
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12244_ _12251_/CLK _12244_/D vssd1 vssd1 vccd1 vccd1 _12244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11545__B1 _11540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ _12953_/Q _13359_/A vssd1 vssd1 vccd1 vccd1 _12176_/D sky130_fd_sc_hd__xor2_1
XFILLER_3_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11126_ _11126_/A vssd1 vssd1 vccd1 vccd1 _12709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13229__385 vssd1 vssd1 vccd1 vccd1 _13229__385/HI _13868_/A sky130_fd_sc_hd__conb_1
XFILLER_96_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11057_ _13817_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11057_/X sky130_fd_sc_hd__or2_1
XANTENNA__09061__S1 _08942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10008_ _10021_/D _10029_/C _10029_/D _10008_/D vssd1 vssd1 vccd1 vccd1 _10016_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA_output49_A _13953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11959_ _11959_/A vssd1 vssd1 vccd1 vccd1 _12913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13629_ _13629_/A _07283_/X vssd1 vssd1 vccd1 vccd1 _14077_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_158_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater61 _14072_/Z vssd1 vssd1 vccd1 vccd1 _14104_/Z sky130_fd_sc_hd__buf_12
Xrepeater72 _14100_/Z vssd1 vssd1 vccd1 vccd1 _14068_/Z sky130_fd_sc_hd__buf_12
Xrepeater83 _14125_/Z vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__buf_12
XFILLER_164_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07150_ _09614_/A vssd1 vssd1 vccd1 vccd1 _07205_/A sky130_fd_sc_hd__clkbuf_2
Xrepeater94 _14121_/Z vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__buf_12
XFILLER_158_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07081_ _07603_/A vssd1 vssd1 vccd1 vccd1 _07533_/A sky130_fd_sc_hd__buf_2
XFILLER_161_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07983_ _07983_/A _08062_/B _08002_/C vssd1 vssd1 vccd1 vccd1 _07984_/A sky130_fd_sc_hd__or3_1
XFILLER_141_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09722_ _12347_/Q _13557_/A vssd1 vssd1 vccd1 vccd1 _09725_/B sky130_fd_sc_hd__xor2_1
XFILLER_86_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06934_ _06936_/A _06941_/B vssd1 vssd1 vccd1 vccd1 _06935_/A sky130_fd_sc_hd__or2_1
XANTENNA__09052__S1 _08913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater71_A peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ _14109_/Z _09653_/B vssd1 vssd1 vccd1 vccd1 _09653_/X sky130_fd_sc_hd__or2_1
XFILLER_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06865_ _06879_/A vssd1 vssd1 vccd1 vccd1 _06877_/A sky130_fd_sc_hd__clkbuf_1
X_08604_ _09981_/B _12424_/Q _12425_/Q _12426_/Q _08602_/X _08603_/X vssd1 vssd1 vccd1
+ vccd1 _08604_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10688__C _10688_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09584_ _09584_/A vssd1 vssd1 vccd1 vccd1 _12323_/D sky130_fd_sc_hd__clkbuf_1
X_06796_ _06809_/A vssd1 vssd1 vccd1 vccd1 _06806_/C sky130_fd_sc_hd__clkbuf_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _11708_/B vssd1 vssd1 vccd1 vccd1 _13372_/A sky130_fd_sc_hd__buf_6
XFILLER_70_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13022__178 vssd1 vssd1 vccd1 vccd1 _13022__178/HI _13449_/A sky130_fd_sc_hd__conb_1
XANTENNA__13361__A _13361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08466_ _13395_/A vssd1 vssd1 vccd1 vccd1 _08517_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07417_ _07417_/A _07423_/B vssd1 vssd1 vccd1 vccd1 _07418_/A sky130_fd_sc_hd__or2_1
X_08397_ _13393_/A vssd1 vssd1 vccd1 vccd1 _08397_/X sky130_fd_sc_hd__buf_2
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07348_ _07348_/A vssd1 vssd1 vccd1 vccd1 _07348_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08866__S1 _08735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07279_ _07279_/A _07289_/B _07286_/C vssd1 vssd1 vccd1 vccd1 _07280_/A sky130_fd_sc_hd__or3_1
XFILLER_128_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09018_ _10938_/A vssd1 vssd1 vccd1 vccd1 _13939_/A sky130_fd_sc_hd__buf_6
XFILLER_3_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10290_ _10288_/X _10278_/X _10289_/X _10283_/X vssd1 vssd1 vccd1 vccd1 _12498_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09733__B _13559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13980_ _13980_/A _06341_/X vssd1 vssd1 vccd1 vccd1 _14012_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_93_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07534__A _07590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12931_ _12952_/CLK _12931_/D vssd1 vssd1 vccd1 vccd1 _12931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11056__A _11070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__B _08349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12862_ _12873_/CLK _12862_/D vssd1 vssd1 vccd1 vccd1 _12862_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _11816_/A _11813_/B vssd1 vssd1 vccd1 vccd1 _11814_/A sky130_fd_sc_hd__and2_1
XFILLER_73_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10895__A _10895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _12799_/CLK _12793_/D vssd1 vssd1 vccd1 vccd1 _13967_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11757_/A _11744_/B vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__and2_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11503__B _11503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11675_ _11688_/A _11672_/X _11576_/X vssd1 vssd1 vccd1 vccd1 _11679_/A sky130_fd_sc_hd__o21ai_1
XFILLER_14_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13414_ _13414_/A _08179_/X vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10626_ _12574_/Q _13750_/A vssd1 vssd1 vccd1 vccd1 _10627_/D sky130_fd_sc_hd__xor2_1
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10557_ _13711_/A _12567_/Q _10635_/B vssd1 vssd1 vccd1 vccd1 _10558_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09196__A _09269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10488_ _12547_/Q _13756_/A vssd1 vssd1 vccd1 vccd1 _10488_/Y sky130_fd_sc_hd__xnor2_1
X_12227_ _12325_/CLK _12227_/D vssd1 vssd1 vccd1 vccd1 _13404_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_142_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09924__A _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ _12964_/Q _13370_/A vssd1 vssd1 vccd1 vccd1 _12161_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07147__C _07969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11109_ _11112_/A _11109_/B vssd1 vssd1 vccd1 vccd1 _11110_/A sky130_fd_sc_hd__and2_1
XFILLER_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12089_ _12101_/B vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_96_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07444__A _07468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06650_ _06650_/A vssd1 vssd1 vccd1 vccd1 _06650_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06581_ _06581_/A vssd1 vssd1 vccd1 vccd1 _06581_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08320_ _08320_/A vssd1 vssd1 vccd1 vccd1 _08320_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08251_ _08251_/A _08261_/B _08251_/C vssd1 vssd1 vccd1 vccd1 _08252_/A sky130_fd_sc_hd__or3_1
X_07202_ _07230_/A vssd1 vssd1 vccd1 vccd1 _07213_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_158_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08182_ _08184_/A _08182_/B _08184_/C vssd1 vssd1 vccd1 vccd1 _08183_/A sky130_fd_sc_hd__or3_1
XFILLER_118_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07133_ _08035_/A vssd1 vssd1 vccd1 vccd1 _07615_/A sky130_fd_sc_hd__buf_2
XANTENNA__09965__A3 _09867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07064_ _08035_/A vssd1 vssd1 vccd1 vccd1 _07120_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07966_ _08004_/A vssd1 vssd1 vccd1 vccd1 _07977_/C sky130_fd_sc_hd__buf_2
XFILLER_114_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09705_ _09705_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _09706_/A sky130_fd_sc_hd__and2_1
XFILLER_56_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06917_ _06917_/A vssd1 vssd1 vccd1 vccd1 _06917_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07897_ _07908_/A _07903_/B _07903_/C vssd1 vssd1 vccd1 vccd1 _07898_/A sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_94_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _12386_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09636_ _09636_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09636_/X sky130_fd_sc_hd__or2_1
XFILLER_71_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06848_ _06850_/A _06857_/B _06857_/C vssd1 vssd1 vccd1 vccd1 _06849_/A sky130_fd_sc_hd__or3_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09567_ _09579_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__and2_1
X_06779_ _06779_/A vssd1 vssd1 vccd1 vccd1 _06779_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08518_ _08458_/X _08461_/X _08488_/X _08516_/X _08511_/X _08517_/X vssd1 vssd1 vccd1
+ vccd1 _08518_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09498_ _09625_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _09498_/X sky130_fd_sc_hd__or2_1
XFILLER_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08449_ _13395_/A vssd1 vssd1 vccd1 vccd1 _08449_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11460_ _11460_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _11474_/A sky130_fd_sc_hd__nand2_1
XFILLER_137_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ _13657_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10411_/X sky130_fd_sc_hd__or2_1
XFILLER_137_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11391_ _12770_/Q _13945_/A vssd1 vssd1 vccd1 vccd1 _11395_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09728__B _13566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10881__C _10881_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10342_ _13660_/A _12514_/Q _10342_/S vssd1 vssd1 vccd1 vccd1 _10343_/B sky130_fd_sc_hd__mux2_1
XFILLER_136_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10273_ _09767_/X _10264_/X _10272_/X _10270_/X vssd1 vssd1 vccd1 vccd1 _12492_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12012_ _12929_/Q _14072_/A _12012_/S vssd1 vssd1 vccd1 vccd1 _12013_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09744__A _09789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09463__B _13557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13963_ _13963_/A _06388_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12914_ _12914_/CLK _12914_/D vssd1 vssd1 vccd1 vccd1 _14041_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13894_ _13894_/A _06573_/X vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12845_ _12850_/CLK _12845_/D vssd1 vssd1 vccd1 vccd1 _12845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12776_/CLK _12776_/D vssd1 vssd1 vccd1 vccd1 _13951_/A sky130_fd_sc_hd__dfxtp_4
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08095__A _08110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13350__506 vssd1 vssd1 vccd1 vccd1 _13350__506/HI _14119_/A sky130_fd_sc_hd__conb_1
X_11727_ _11740_/A _11727_/B vssd1 vssd1 vccd1 vccd1 _11728_/A sky130_fd_sc_hd__and2_1
XFILLER_159_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11658_ _11658_/A _11688_/B _11676_/C vssd1 vssd1 vccd1 vccd1 _11659_/B sky130_fd_sc_hd__and3_1
XFILLER_30_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10609_ _10952_/A _10609_/B vssd1 vssd1 vccd1 vccd1 _10610_/A sky130_fd_sc_hd__and2_1
X_11589_ _11631_/C _11587_/A _11540_/X vssd1 vssd1 vccd1 vccd1 _11590_/B sky130_fd_sc_hd__o21ai_1
XFILLER_143_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13244__400 vssd1 vssd1 vccd1 vccd1 _13244__400/HI _13899_/A sky130_fd_sc_hd__conb_1
XFILLER_111_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07820_ _07868_/A _07820_/B _08110_/C vssd1 vssd1 vccd1 vccd1 _07821_/A sky130_fd_sc_hd__or3_1
XFILLER_38_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07751_ _07756_/A _07753_/B _07761_/C vssd1 vssd1 vccd1 vccd1 _07752_/A sky130_fd_sc_hd__or3_1
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_92_clk_A _12438_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_76_clk _12555_/CLK vssd1 vssd1 vccd1 vccd1 _12656_/CLK sky130_fd_sc_hd__clkbuf_16
X_06702_ _06702_/A vssd1 vssd1 vccd1 vccd1 _06702_/X sky130_fd_sc_hd__clkbuf_1
X_07682_ _07682_/A vssd1 vssd1 vccd1 vccd1 _07682_/X sky130_fd_sc_hd__clkbuf_1
X_09421_ _13428_/A _12280_/Q _09431_/S vssd1 vssd1 vccd1 vccd1 _09422_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06633_ _06633_/A vssd1 vssd1 vccd1 vccd1 _07995_/B sky130_fd_sc_hd__buf_2
XFILLER_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09352_ _09362_/D _09352_/B _09352_/C _09352_/D vssd1 vssd1 vccd1 vccd1 _09355_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_80_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06564_ _08182_/B vssd1 vssd1 vccd1 vccd1 _06574_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_21_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08303_ _08312_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08304_/A sky130_fd_sc_hd__or2_1
X_13093__249 vssd1 vssd1 vccd1 vccd1 _13093__249/HI _13602_/A sky130_fd_sc_hd__conb_1
XFILLER_21_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09283_ _09322_/B _09276_/X _09282_/Y vssd1 vssd1 vccd1 vccd1 _12248_/D sky130_fd_sc_hd__a21oi_1
X_06495_ _06495_/A vssd1 vssd1 vccd1 vccd1 _06495_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08234_ _08234_/A vssd1 vssd1 vccd1 vccd1 _08234_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_30_clk_A _12759_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08165_ _08165_/A vssd1 vssd1 vccd1 vccd1 _08165_/X sky130_fd_sc_hd__clkbuf_1
X_07116_ _07116_/A vssd1 vssd1 vccd1 vccd1 _07116_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08096_ _08096_/A vssd1 vssd1 vccd1 vccd1 _08096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07047_ _07055_/A _07055_/B vssd1 vssd1 vccd1 vccd1 _07048_/A sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_45_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08998_ _12826_/Q vssd1 vssd1 vccd1 vccd1 _11631_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07949_ _08064_/A vssd1 vssd1 vccd1 vccd1 _07971_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13028__184 vssd1 vssd1 vccd1 vccd1 _13028__184/HI _13471_/A sky130_fd_sc_hd__conb_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_67_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _12515_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10960_ _10969_/A _10960_/B vssd1 vssd1 vccd1 vccd1 _10961_/A sky130_fd_sc_hd__and2_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07812__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09619_ _13456_/A _09613_/X _09618_/X _09522_/X vssd1 vssd1 vccd1 vccd1 _12326_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10891_ _10897_/C _10891_/B vssd1 vssd1 vccd1 vccd1 _10891_/Y sky130_fd_sc_hd__nand2_1
X_12630_ _12634_/CLK _12630_/D vssd1 vssd1 vccd1 vccd1 _12630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_118_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12561_ _12565_/CLK _12561_/D vssd1 vssd1 vccd1 vccd1 _13689_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ _11514_/B _11512_/B _11682_/B vssd1 vssd1 vccd1 vccd1 _11513_/A sky130_fd_sc_hd__and3b_1
XFILLER_129_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12492_ _12492_/CLK _12492_/D vssd1 vssd1 vccd1 vccd1 _13622_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11443_ _11443_/A vssd1 vssd1 vccd1 vccd1 _12084_/A sky130_fd_sc_hd__buf_4
XANTENNA__09458__B _13552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08362__B _08364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11374_ _11377_/A _11374_/B vssd1 vssd1 vccd1 vccd1 _11375_/A sky130_fd_sc_hd__and2_1
XFILLER_137_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10325_ _10332_/A _10325_/B vssd1 vssd1 vccd1 vccd1 _10326_/A sky130_fd_sc_hd__and2_1
XFILLER_113_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14093_ _14093_/A _08155_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[30] sky130_fd_sc_hd__ebufn_8
XFILLER_124_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10256_ _10256_/A vssd1 vssd1 vccd1 vccd1 _10256_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater102_A _14117_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ _13620_/A _12473_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__mux2_1
XFILLER_79_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_58_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _12835_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_clk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_81_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13946_ _13946_/A _06432_/X vssd1 vssd1 vccd1 vccd1 _13978_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output31_A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13877_ _13877_/A _06622_/X vssd1 vssd1 vccd1 vccd1 _14069_/Z sky130_fd_sc_hd__ebufn_8
X_12828_ _12829_/CLK _12828_/D vssd1 vssd1 vccd1 vccd1 _12828_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06338__A _06462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12759_ _12759_/CLK _12759_/D vssd1 vssd1 vccd1 vccd1 _13886_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06280_ _06442_/A vssd1 vssd1 vccd1 vccd1 _07845_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11188__A1 _11184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11410__C _11410_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09970_ _12421_/Q _10160_/A vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__and2b_1
XFILLER_115_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08921_ _13968_/A vssd1 vssd1 vccd1 vccd1 _08921_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10699__A0 _14097_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ _12650_/Q vssd1 vssd1 vccd1 vccd1 _10907_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08987__S0 _08911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07803_ _07817_/A vssd1 vssd1 vccd1 vccd1 _07815_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08783_ _12624_/Q _12625_/Q _12626_/Q _12627_/Q _08739_/X _08740_/X vssd1 vssd1 vccd1
+ vccd1 _08783_/X sky130_fd_sc_hd__mux4_2
XFILLER_111_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _12593_/CLK sky130_fd_sc_hd__clkbuf_16
X_07734_ _07763_/A vssd1 vssd1 vccd1 vccd1 _07748_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07665_ _07665_/A vssd1 vssd1 vccd1 vccd1 _07665_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ _09404_/A _09404_/B vssd1 vssd1 vccd1 vccd1 _09405_/A sky130_fd_sc_hd__and2_1
X_06616_ _06625_/A _06616_/B _06616_/C vssd1 vssd1 vccd1 vccd1 _06617_/A sky130_fd_sc_hd__or3_1
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07596_ _07601_/A _07598_/B _07608_/C vssd1 vssd1 vccd1 vccd1 _07597_/A sky130_fd_sc_hd__or3_1
XFILLER_71_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ _09368_/B vssd1 vssd1 vccd1 vccd1 _09363_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06547_ _06547_/A vssd1 vssd1 vccd1 vccd1 _07323_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ _09328_/C _09332_/B _09206_/X vssd1 vssd1 vccd1 vccd1 _09266_/Y sky130_fd_sc_hd__o21ai_1
X_06478_ _06478_/A vssd1 vssd1 vccd1 vccd1 _06478_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08217_ _08217_/A vssd1 vssd1 vccd1 vccd1 _08217_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09197_ _09281_/A vssd1 vssd1 vccd1 vccd1 _09263_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__09278__B _09389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08148_ _08148_/A _08151_/B _08151_/C vssd1 vssd1 vccd1 vccd1 _08149_/A sky130_fd_sc_hd__or3_1
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08079_ _09484_/A vssd1 vssd1 vccd1 vccd1 _11026_/B sky130_fd_sc_hd__buf_6
XFILLER_161_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10110_ _10111_/B _10108_/B _10109_/Y vssd1 vssd1 vccd1 vccd1 _12454_/D sky130_fd_sc_hd__a21oi_1
XFILLER_134_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11090_ _11090_/A vssd1 vssd1 vccd1 vccd1 _12698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11329__A _11381_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _10041_/A vssd1 vssd1 vccd1 vccd1 _12438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11763__S _11763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13544__A _13544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13800_ _13800_/A _06837_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
X_11992_ _12923_/Q _14066_/A _11995_/S vssd1 vssd1 vccd1 vccd1 _11993_/B sky130_fd_sc_hd__mux2_1
X_10943_ _13980_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _10996_/S sky130_fd_sc_hd__and2_2
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13731_ _13731_/A _07014_/X vssd1 vssd1 vccd1 vccd1 _13987_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11064__A _11064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_13662_ _13662_/A _07194_/X vssd1 vssd1 vccd1 vccd1 _14078_/Z sky130_fd_sc_hd__ebufn_8
X_10874_ _10874_/A _10874_/B _10874_/C vssd1 vssd1 vccd1 vccd1 _10877_/B sky130_fd_sc_hd__and3_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11999__A _12033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12613_ _12802_/CLK _12613_/D vssd1 vssd1 vccd1 vccd1 _13788_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13593_ _13593_/A _07383_/X vssd1 vssd1 vccd1 vccd1 _13625_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12544_ _12599_/CLK _12544_/D vssd1 vssd1 vccd1 vccd1 _12544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12475_ _12656_/CLK _12475_/D vssd1 vssd1 vccd1 vccd1 _12475_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10408__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11426_ _11452_/B vssd1 vssd1 vccd1 vccd1 _11436_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11357_ _11361_/A _11357_/B vssd1 vssd1 vccd1 vccd1 _11358_/A sky130_fd_sc_hd__and2_1
XFILLER_125_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ _10315_/A _10308_/B vssd1 vssd1 vccd1 vccd1 _10309_/A sky130_fd_sc_hd__and2_1
XFILLER_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14076_ _14076_/A _08029_/X vssd1 vssd1 vccd1 vccd1 _14108_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_152_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11288_ _11153_/X _11284_/X _11287_/X _11195_/X vssd1 vssd1 vccd1 vccd1 _12744_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08969__S0 _08967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ _12472_/Q _13747_/A vssd1 vssd1 vccd1 vccd1 _10242_/B sky130_fd_sc_hd__xor2_1
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09932__A _09939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13356__512 vssd1 vssd1 vccd1 vccd1 _13356__512/HI _14125_/A sky130_fd_sc_hd__conb_1
X_13929_ _13929_/A _06478_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[26] sky130_fd_sc_hd__ebufn_8
XFILLER_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07450_ _07454_/A _07459_/B vssd1 vssd1 vccd1 vccd1 _07451_/A sky130_fd_sc_hd__or2_1
XFILLER_62_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06401_ _06401_/A vssd1 vssd1 vccd1 vccd1 _06401_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07381_ _07381_/A vssd1 vssd1 vccd1 vccd1 _07381_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09120_ _10552_/A vssd1 vssd1 vccd1 vccd1 _09120_/X sky130_fd_sc_hd__buf_4
XANTENNA__09379__A _09379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06332_ _06332_/A vssd1 vssd1 vccd1 vccd1 _06332_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09051_ _12846_/Q vssd1 vssd1 vccd1 vccd1 _11688_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06263_ input20/X input22/X input21/X _06263_/D vssd1 vssd1 vccd1 vccd1 _09096_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_129_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08002_ _08010_/A _08005_/B _08002_/C vssd1 vssd1 vccd1 vccd1 _08003_/A sky130_fd_sc_hd__or3_1
XFILLER_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11581__A1 _11634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09953_ _14104_/Z _13592_/A _09953_/S vssd1 vssd1 vccd1 vccd1 _09954_/B sky130_fd_sc_hd__mux2_1
XFILLER_58_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08904_ _08809_/X _08818_/X _08815_/X _08822_/X _08769_/X _08850_/X vssd1 vssd1 vccd1
+ vccd1 _08904_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10053__A _13583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _13522_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09884_/X sky130_fd_sc_hd__or2_1
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _08832_/X _08834_/X _13780_/A vssd1 vssd1 vccd1 vccd1 _10162_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10988__A _10988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13364__A _13364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ _13776_/A vssd1 vssd1 vccd1 vccd1 _08766_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ _07727_/A _07724_/B _07719_/C vssd1 vssd1 vccd1 vccd1 _07718_/A sky130_fd_sc_hd__or3_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _12460_/Q vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13099__255 vssd1 vssd1 vccd1 vccd1 _13099__255/HI _13608_/A sky130_fd_sc_hd__conb_1
XANTENNA__10500__B _13751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07648_ _07648_/A vssd1 vssd1 vccd1 vccd1 _07648_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07579_ _07579_/A vssd1 vssd1 vccd1 vccd1 _07579_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09318_ _09318_/A _09318_/B _09318_/C _09318_/D vssd1 vssd1 vccd1 vccd1 _09336_/B
+ sky130_fd_sc_hd__and4_1
X_10590_ _10602_/A _10590_/B vssd1 vssd1 vccd1 vccd1 _10591_/A sky130_fd_sc_hd__and2_1
X_09249_ _09315_/B _09253_/C _09248_/X vssd1 vssd1 vccd1 vccd1 _09251_/A sky130_fd_sc_hd__o21ai_1
X_12260_ _12264_/CLK _12260_/D vssd1 vssd1 vccd1 vccd1 _12260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11211_ _11221_/A _11211_/B vssd1 vssd1 vccd1 vccd1 _11212_/A sky130_fd_sc_hd__and2_1
XFILLER_107_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12191_ _14099_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12191_/X sky130_fd_sc_hd__or2_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput32 _13978_/A vssd1 vssd1 vccd1 vccd1 pwm_en[13] sky130_fd_sc_hd__buf_2
X_11142_ _12696_/Q _13937_/A vssd1 vssd1 vccd1 vccd1 _11143_/D sky130_fd_sc_hd__xor2_1
Xoutput43 _13786_/A vssd1 vssd1 vccd1 vccd1 pwm_en[9] sky130_fd_sc_hd__buf_2
Xoutput54 _13567_/A vssd1 vssd1 vccd1 vccd1 pwm_out[4] sky130_fd_sc_hd__buf_2
XFILLER_1_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12162__B _13362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _11124_/S vssd1 vssd1 vccd1 vccd1 _11151_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_49_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11324__A1 _10548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10024_ _10029_/B _10024_/B _10024_/C vssd1 vssd1 vccd1 vccd1 _10024_/X sky130_fd_sc_hd__and3_1
XFILLER_48_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09471__B _13566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11975_ _11978_/A _11975_/B vssd1 vssd1 vccd1 vccd1 _11976_/A sky130_fd_sc_hd__and2_1
XFILLER_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13714_ _13714_/A _07054_/X vssd1 vssd1 vccd1 vccd1 _14098_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_32_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926_ _10928_/B _10928_/C _10798_/X vssd1 vssd1 vccd1 vccd1 _10927_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13645_ _13645_/A _07240_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
X_10857_ _10857_/A vssd1 vssd1 vccd1 vccd1 _12641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13576_ _13576_/A _07429_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
X_10788_ _10788_/A vssd1 vssd1 vccd1 vccd1 _12624_/D sky130_fd_sc_hd__clkbuf_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12527_ _12583_/CLK _12527_/D vssd1 vssd1 vccd1 vccd1 _13656_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09927__A _09982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ _12461_/CLK _12458_/D vssd1 vssd1 vccd1 vccd1 _12458_/Q sky130_fd_sc_hd__dfxtp_1
X_11409_ _11409_/A vssd1 vssd1 vccd1 vccd1 _12776_/D sky130_fd_sc_hd__clkbuf_1
X_12389_ _12400_/CLK _12389_/D vssd1 vssd1 vccd1 vccd1 _12389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06351__A _06462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06950_ _06974_/A vssd1 vssd1 vccd1 vccd1 _06960_/A sky130_fd_sc_hd__clkbuf_1
X_14059_ _14059_/A _07940_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
XANTENNA__11315__A1 _11184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06881_ _06881_/A vssd1 vssd1 vccd1 vccd1 _06881_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08620_ _08614_/X _08615_/X _08617_/X _08619_/X _08583_/X _08584_/X vssd1 vssd1 vccd1
+ vccd1 _08620_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08551_ _08709_/A vssd1 vssd1 vccd1 vccd1 _08551_/X sky130_fd_sc_hd__buf_2
XFILLER_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07502_ _07504_/A _07504_/B _07510_/C vssd1 vssd1 vccd1 vccd1 _07503_/A sky130_fd_sc_hd__or3_1
XFILLER_23_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08482_ _09352_/B _09362_/D _12264_/Q _12265_/Q _08373_/X _08374_/X vssd1 vssd1 vccd1
+ vccd1 _08482_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07433_ _07442_/A _07435_/B vssd1 vssd1 vccd1 vccd1 _07434_/A sky130_fd_sc_hd__or2_1
XANTENNA__07910__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07364_ _07369_/A _07364_/B _07374_/C vssd1 vssd1 vccd1 vccd1 _07365_/A sky130_fd_sc_hd__or3_1
X_09103_ _12208_/B vssd1 vssd1 vccd1 vccd1 _12180_/B sky130_fd_sc_hd__clkbuf_2
X_06315_ _06315_/A vssd1 vssd1 vccd1 vccd1 _06315_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07295_ _07519_/A vssd1 vssd1 vccd1 vccd1 _07307_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_164_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09034_ _12844_/Q vssd1 vssd1 vccd1 vccd1 _11676_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13359__A _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06261__A input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09936_ _09936_/A vssd1 vssd1 vccd1 vccd1 _12410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _12378_/Q _09867_/B vssd1 vssd1 vccd1 vccd1 _09868_/D sky130_fd_sc_hd__xor2_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08818_ _10876_/C _12638_/Q _10875_/B _10876_/B _08807_/X _08808_/X vssd1 vssd1 vccd1
+ vccd1 _08818_/X sky130_fd_sc_hd__mux4_2
XFILLER_133_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09798_ _09798_/A vssd1 vssd1 vccd1 vccd1 _12375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08188__A _08228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _13779_/A vssd1 vssd1 vccd1 vccd1 _08749_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10230__B _13746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _12868_/Q _14013_/A _11760_/S vssd1 vssd1 vccd1 vccd1 _11761_/B sky130_fd_sc_hd__mux2_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08486__A1 _08447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07820__A _07868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _11039_/A vssd1 vssd1 vccd1 vccd1 _10711_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11691_ _11691_/A vssd1 vssd1 vccd1 vccd1 _12849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11342__A _11381_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13430_ _13430_/A _07805_/X vssd1 vssd1 vccd1 vccd1 _14102_/Z sky130_fd_sc_hd__ebufn_8
X_10642_ _10377_/X _10638_/X _10641_/X _10550_/X vssd1 vssd1 vccd1 vccd1 _12584_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12157__B _13368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__C _08360_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ _13361_/A _08282_/X vssd1 vssd1 vccd1 vccd1 _14065_/Z sky130_fd_sc_hd__ebufn_8
X_10573_ _10585_/A _10573_/B vssd1 vssd1 vccd1 vccd1 _10574_/A sky130_fd_sc_hd__and2_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12312_ _12313_/CLK _12312_/D vssd1 vssd1 vccd1 vccd1 _12312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12243_ _12251_/CLK _12243_/D vssd1 vssd1 vccd1 vccd1 _12243_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09466__B _13565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12174_ _12957_/Q _13363_/A vssd1 vssd1 vccd1 vccd1 _12176_/C sky130_fd_sc_hd__xor2_1
XFILLER_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11125_ _11204_/A _11125_/B vssd1 vssd1 vccd1 vccd1 _11126_/A sky130_fd_sc_hd__and2_1
XFILLER_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09482__A _11026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ _11070_/B vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__09910__A1 _09092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _10022_/A _10007_/B vssd1 vssd1 vccd1 vccd1 _12430_/D sky130_fd_sc_hd__nor2_1
XFILLER_92_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11958_ _11962_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11959_/A sky130_fd_sc_hd__and2_1
XFILLER_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11652__C_N _11515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10284__A1 _09186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ _10909_/A _10909_/B _10922_/C vssd1 vssd1 vccd1 vccd1 _10909_/X sky130_fd_sc_hd__and3_1
X_11889_ _12899_/Q _14043_/A _11895_/S vssd1 vssd1 vccd1 vccd1 _11890_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13628_ _13628_/A _07285_/X vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_8
Xrepeater62 peripheralBus_data[9] vssd1 vssd1 vccd1 vccd1 _14072_/Z sky130_fd_sc_hd__buf_12
Xrepeater73 peripheralBus_data[5] vssd1 vssd1 vccd1 vccd1 _14100_/Z sky130_fd_sc_hd__buf_12
Xrepeater84 peripheralBus_data[30] vssd1 vssd1 vccd1 vccd1 _14125_/Z sky130_fd_sc_hd__buf_12
Xrepeater95 peripheralBus_data[26] vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__buf_12
X_13559_ _13559_/A _07470_/X vssd1 vssd1 vccd1 vccd1 _13623_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_9_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09657__A _13594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07080_ _07080_/A vssd1 vssd1 vccd1 vccd1 _07080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07982_ _08004_/A vssd1 vssd1 vccd1 vccd1 _08002_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09392__A _09392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ _12351_/Q _13561_/A vssd1 vssd1 vccd1 vccd1 _09725_/A sky130_fd_sc_hd__xor2_1
X_06933_ _06933_/A vssd1 vssd1 vccd1 vccd1 _06933_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09901__A1 _09773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _13468_/A _09640_/X _09651_/X _09649_/X vssd1 vssd1 vccd1 vccd1 _12338_/D
+ sky130_fd_sc_hd__o211a_1
X_06864_ _06864_/A vssd1 vssd1 vccd1 vccd1 _06864_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater64_A peripheralBus_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ _08709_/A vssd1 vssd1 vccd1 vccd1 _08603_/X sky130_fd_sc_hd__buf_2
XFILLER_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11146__B _13943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09583_ _09669_/A _09583_/B vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__and2_1
X_06795_ _06832_/A vssd1 vssd1 vccd1 vccd1 _06806_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08534_ _08530_/X _08533_/X _09162_/A vssd1 vssd1 vccd1 vccd1 _11708_/B sky130_fd_sc_hd__mux2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10275__A1 _09770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ _11706_/D vssd1 vssd1 vccd1 vccd1 _13362_/A sky130_fd_sc_hd__buf_4
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07416_ _07416_/A vssd1 vssd1 vccd1 vccd1 _07416_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08396_ _13392_/A vssd1 vssd1 vccd1 vccd1 _08396_/X sky130_fd_sc_hd__clkbuf_4
X_07347_ _07356_/A _07351_/B _07347_/C vssd1 vssd1 vccd1 vccd1 _07348_/A sky130_fd_sc_hd__or3_1
XFILLER_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07278_ _07291_/A vssd1 vssd1 vccd1 vccd1 _07289_/B sky130_fd_sc_hd__clkbuf_1
X_09017_ _09014_/X _09016_/X _13972_/A vssd1 vssd1 vccd1 vccd1 _10938_/A sky130_fd_sc_hd__mux2_2
XFILLER_128_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10225__B _13752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13261__417 vssd1 vssd1 vccd1 vccd1 _13261__417/HI _13932_/A sky130_fd_sc_hd__conb_1
XANTENNA__07815__A _07868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ _09925_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09937_/A sky130_fd_sc_hd__nand2_2
XFILLER_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12930_ _12952_/CLK _12930_/D vssd1 vssd1 vccd1 vccd1 _12930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13302__458 vssd1 vssd1 vccd1 vccd1 _13302__458/HI _14023_/A sky130_fd_sc_hd__conb_1
XFILLER_160_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12867_/CLK _12861_/D vssd1 vssd1 vccd1 vccd1 _12861_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13552__A _13552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _09631_/A _14005_/A _11823_/S vssd1 vssd1 vccd1 vccd1 _11813_/B sky130_fd_sc_hd__mux2_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12938_/CLK _12792_/D vssd1 vssd1 vccd1 vccd1 _13918_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _12863_/Q _14008_/A _11743_/S vssd1 vssd1 vccd1 vccd1 _11744_/B sky130_fd_sc_hd__mux2_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13155__311 vssd1 vssd1 vccd1 vccd1 _13155__311/HI _13728_/A sky130_fd_sc_hd__conb_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11072__A _13979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _11670_/Y _11668_/C _11673_/X vssd1 vssd1 vccd1 vccd1 _12845_/D sky130_fd_sc_hd__a21oi_1
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13413_ _13413_/A _08175_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
XFILLER_155_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10625_ _12569_/Q _13745_/A vssd1 vssd1 vccd1 vccd1 _10627_/C sky130_fd_sc_hd__xor2_1
XFILLER_127_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10556_ _10608_/S vssd1 vssd1 vccd1 vccd1 _10635_/B sky130_fd_sc_hd__buf_2
XFILLER_10_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09196__B _11503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater132_A peripheralBus_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10487_ _12535_/Q _13744_/A vssd1 vssd1 vccd1 vccd1 _10487_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12226_ _12325_/CLK _12226_/D vssd1 vssd1 vccd1 vccd1 _13403_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__11923__D1 _13403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _12962_/Q _13368_/A vssd1 vssd1 vccd1 vccd1 _12161_/A sky130_fd_sc_hd__xor2_1
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ _13849_/A _12704_/Q _11118_/S vssd1 vssd1 vccd1 vccd1 _11109_/B sky130_fd_sc_hd__mux2_1
XFILLER_150_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12088_ _12088_/A vssd1 vssd1 vccd1 vccd1 _12088_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11039_ _11039_/A vssd1 vssd1 vccd1 vccd1 _11039_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06580_ _06584_/A _06589_/B _06589_/C vssd1 vssd1 vccd1 vccd1 _06581_/A sky130_fd_sc_hd__or3_1
XANTENNA__10257__A1 _09139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08250_ _08263_/A vssd1 vssd1 vccd1 vccd1 _08261_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07201_ _07201_/A vssd1 vssd1 vccd1 vccd1 _07201_/X sky130_fd_sc_hd__clkbuf_1
X_08181_ _08181_/A vssd1 vssd1 vccd1 vccd1 _08181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07132_ _07132_/A vssd1 vssd1 vccd1 vccd1 _07132_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06804__A _07857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07063_ _08177_/A vssd1 vssd1 vccd1 vccd1 _08180_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11509__A1 _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07965_ _08084_/A vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_68_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11157__A _11199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _13500_/A _12354_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09705_/B sky130_fd_sc_hd__mux2_1
XFILLER_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06916_ _06923_/A _06916_/B vssd1 vssd1 vccd1 vccd1 _06917_/A sky130_fd_sc_hd__or2_1
XFILLER_56_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07896_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07908_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__11693__B1 _11569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _13462_/A _09627_/X _09633_/X _09634_/X vssd1 vssd1 vccd1 vccd1 _12332_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_4_clk_A _12917_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06847_ _06967_/A vssd1 vssd1 vccd1 vccd1 _06857_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_82_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13372__A _13372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ _13465_/A _12318_/Q _09575_/S vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__mux2_1
XFILLER_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06778_ _06788_/A _06780_/B _06780_/C vssd1 vssd1 vccd1 vccd1 _06779_/A sky130_fd_sc_hd__or3_1
XFILLER_70_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11604__B _11604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ _08517_/A vssd1 vssd1 vccd1 vccd1 _08517_/X sky130_fd_sc_hd__clkbuf_2
X_09497_ _13426_/A _09483_/X _09492_/X _09496_/X vssd1 vssd1 vccd1 vccd1 _12295_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ _13394_/A vssd1 vssd1 vccd1 vccd1 _08448_/X sky130_fd_sc_hd__buf_2
XFILLER_135_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08379_ _13392_/A vssd1 vssd1 vccd1 vccd1 _08379_/X sky130_fd_sc_hd__buf_2
X_10410_ _10423_/B vssd1 vssd1 vccd1 vccd1 _10421_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_136_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ _11385_/Y _11386_/X _11387_/Y _11388_/X _11389_/Y vssd1 vssd1 vccd1 vccd1
+ _11390_/X sky130_fd_sc_hd__o221a_1
XFILLER_99_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10341_ _10341_/A vssd1 vssd1 vccd1 vccd1 _12513_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10420__A1 _10288_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10272_ _13622_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10272_/X sky130_fd_sc_hd__or2_1
XFILLER_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12011_ _12011_/A vssd1 vssd1 vccd1 vccd1 _12928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12170__B _13371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13962_ _13962_/A _06392_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
XFILLER_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09760__A _09789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ _12914_/CLK _12913_/D vssd1 vssd1 vccd1 vccd1 _14040_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11684__B1 _11505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ _13893_/A _06575_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
XFILLER_62_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _12850_/CLK _12844_/D vssd1 vssd1 vccd1 vccd1 _12844_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12775_/CLK _12775_/D vssd1 vssd1 vccd1 vccd1 _12775_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _12858_/Q _14003_/A _11726_/S vssd1 vssd1 vccd1 vccd1 _11727_/B sky130_fd_sc_hd__mux2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11657_ _11661_/B _11657_/B _11657_/C vssd1 vssd1 vccd1 vccd1 _11676_/C sky130_fd_sc_hd__and3_1
XFILLER_30_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09919__B _09919_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11739__A1 _14007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10608_ _13726_/A _12582_/Q _10608_/S vssd1 vssd1 vccd1 vccd1 _10609_/B sky130_fd_sc_hd__mux2_1
X_11588_ _11631_/C _11631_/D _11602_/C vssd1 vssd1 vccd1 vccd1 _11590_/A sky130_fd_sc_hd__and3_1
XFILLER_127_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10146__A _10146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10539_ _10553_/B vssd1 vssd1 vccd1 vccd1 _10549_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09935__A _09939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12209_ _11189_/X _12195_/A _12208_/X _12200_/X vssd1 vssd1 vccd1 vccd1 _12981_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13324__480 vssd1 vssd1 vccd1 vccd1 _13324__480/HI _14061_/A sky130_fd_sc_hd__conb_1
XFILLER_111_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07750_ _07763_/A vssd1 vssd1 vccd1 vccd1 _07761_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_96_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06701_ _06701_/A _06706_/B _06706_/C vssd1 vssd1 vccd1 vccd1 _06702_/A sky130_fd_sc_hd__or3_1
XANTENNA__11675__B1 _11576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ _07686_/A _07683_/B _07691_/C vssd1 vssd1 vccd1 vccd1 _07682_/A sky130_fd_sc_hd__or3_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09420_ _09420_/A vssd1 vssd1 vccd1 vccd1 _12279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06632_ _06680_/A vssd1 vssd1 vccd1 vccd1 _06651_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09351_ _09362_/D _09347_/X _09248_/X vssd1 vssd1 vccd1 vccd1 _09353_/A sky130_fd_sc_hd__o21ai_1
X_06563_ _06604_/A vssd1 vssd1 vccd1 vccd1 _06574_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_33_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08302_ _08314_/A vssd1 vssd1 vccd1 vccd1 _08312_/A sky130_fd_sc_hd__clkbuf_1
X_09282_ _09322_/B _09276_/X _09392_/A vssd1 vssd1 vccd1 vccd1 _09282_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06494_ _06494_/A _06499_/B _06499_/C vssd1 vssd1 vccd1 vccd1 _06495_/A sky130_fd_sc_hd__or3_1
X_08233_ _08238_/A _08235_/B _08238_/C vssd1 vssd1 vccd1 vccd1 _08234_/A sky130_fd_sc_hd__or3_1
XFILLER_159_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08164_ _08174_/A _08174_/B _08164_/C vssd1 vssd1 vccd1 vccd1 _08165_/A sky130_fd_sc_hd__or3_1
X_07115_ _07121_/A _07118_/B _07115_/C vssd1 vssd1 vccd1 vccd1 _07116_/A sky130_fd_sc_hd__or3_1
XFILLER_107_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08095_ _08110_/A _08113_/B _08105_/C vssd1 vssd1 vccd1 vccd1 _08096_/A sky130_fd_sc_hd__or3_1
XFILLER_69_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07046_ _10637_/A vssd1 vssd1 vccd1 vccd1 _07055_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__13367__A _13367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10503__B _13743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _08985_/X _08987_/X _08991_/X _08993_/X _08994_/X _08996_/X vssd1 vssd1 vccd1
+ vccd1 _08997_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07948_ _07948_/A vssd1 vssd1 vccd1 vccd1 _07948_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07879_ _07892_/A vssd1 vssd1 vccd1 vccd1 _07890_/B sky130_fd_sc_hd__clkbuf_1
X_09618_ _11160_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09618_/X sky130_fd_sc_hd__or2_1
XFILLER_83_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10890_ _13775_/A _10908_/C _10909_/A _10909_/B vssd1 vssd1 vccd1 vccd1 _10897_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__06709__A _06722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09549_ _13460_/A _12313_/Q _09558_/S vssd1 vssd1 vccd1 vccd1 _09550_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12560_ _12565_/CLK _12560_/D vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _11576_/A vssd1 vssd1 vccd1 vccd1 _11682_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_12_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12491_ _12492_/CLK _12491_/D vssd1 vssd1 vccd1 vccd1 _13621_/A sky130_fd_sc_hd__dfxtp_1
X_11442_ _13914_/A _11450_/B vssd1 vssd1 vccd1 vccd1 _11442_/X sky130_fd_sc_hd__or2_1
XFILLER_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12165__B _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11373_ _13916_/A _12773_/Q _11373_/S vssd1 vssd1 vccd1 vccd1 _11374_/B sky130_fd_sc_hd__mux2_1
X_13267__423 vssd1 vssd1 vccd1 vccd1 _13267__423/HI _13958_/A sky130_fd_sc_hd__conb_1
XFILLER_164_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10324_ _13655_/A _12509_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10325_/B sky130_fd_sc_hd__mux2_1
XFILLER_152_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14092_ _14092_/A _08152_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[29] sky130_fd_sc_hd__ebufn_8
XANTENNA__09474__B _13561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _13616_/A _10262_/B vssd1 vssd1 vccd1 vccd1 _10255_/X sky130_fd_sc_hd__or2_1
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13308__464 vssd1 vssd1 vccd1 vccd1 _13308__464/HI _14029_/A sky130_fd_sc_hd__conb_1
X_10186_ _10186_/A vssd1 vssd1 vccd1 vccd1 _12472_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08770__A0 _08763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09490__A _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13945_ _13945_/A _06434_/X vssd1 vssd1 vccd1 vccd1 _14009_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13876_ _13876_/A _06624_/X vssd1 vssd1 vccd1 vccd1 _14068_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__06619__A _06680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12827_ _12829_/CLK _12827_/D vssd1 vssd1 vccd1 vccd1 _12827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12758_/CLK _12758_/D vssd1 vssd1 vccd1 vccd1 _13885_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _11709_/A _11709_/B _11709_/C _11709_/D vssd1 vssd1 vccd1 vccd1 _12103_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_148_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12689_ _12710_/CLK _12689_/D vssd1 vssd1 vccd1 vccd1 _13818_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_155_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08920_ _12815_/Q _12816_/Q _12817_/Q _12818_/Q _08918_/X _08919_/X vssd1 vssd1 vccd1
+ vccd1 _08920_/X sky130_fd_sc_hd__mux4_2
XANTENNA__10604__A _10971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08851_ _08802_/X _08809_/X _08805_/X _08815_/X _08837_/X _08850_/X vssd1 vssd1 vccd1
+ vccd1 _08851_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08987__S1 _08913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07802_ _07802_/A vssd1 vssd1 vccd1 vccd1 _07802_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08782_ _10773_/B _12621_/Q _12622_/Q _12623_/Q _08739_/X _08740_/X vssd1 vssd1 vccd1
+ vccd1 _08782_/X sky130_fd_sc_hd__mux4_2
X_13060__216 vssd1 vssd1 vccd1 vccd1 _13060__216/HI _13535_/A sky130_fd_sc_hd__conb_1
X_07733_ _07733_/A vssd1 vssd1 vccd1 vccd1 _07733_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07664_ _07672_/A _07669_/B _07664_/C vssd1 vssd1 vccd1 vccd1 _07665_/A sky130_fd_sc_hd__or3_1
XANTENNA__06529__A _07507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09403_ _13423_/A _12275_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _09404_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11154__B _11154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06615_ _06615_/A vssd1 vssd1 vccd1 vccd1 _06615_/X sky130_fd_sc_hd__clkbuf_1
X_13101__257 vssd1 vssd1 vccd1 vccd1 _13101__257/HI _13610_/A sky130_fd_sc_hd__conb_1
XFILLER_41_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07595_ _07623_/A vssd1 vssd1 vccd1 vccd1 _07608_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_111_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09334_ _09343_/C _09336_/A _09334_/C _09334_/D vssd1 vssd1 vccd1 vccd1 _09368_/B
+ sky130_fd_sc_hd__and4_1
X_06546_ _06546_/A vssd1 vssd1 vccd1 vccd1 _06546_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11820__A0 _09636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _09322_/D vssd1 vssd1 vccd1 vccd1 _09328_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_06477_ _06481_/A _06486_/B _06486_/C vssd1 vssd1 vccd1 vccd1 _06478_/A sky130_fd_sc_hd__or3_1
XANTENNA__11170__A _11170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08216_ _08225_/A _08222_/B _08225_/C vssd1 vssd1 vccd1 vccd1 _08217_/A sky130_fd_sc_hd__or3_1
X_09196_ _09269_/A _11503_/B _09196_/C vssd1 vssd1 vccd1 vccd1 _09281_/A sky130_fd_sc_hd__and3_2
XANTENNA__06264__A input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08147_ _08147_/A vssd1 vssd1 vccd1 vccd1 _08147_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08078_ _08078_/A vssd1 vssd1 vccd1 vccd1 _08078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07029_ _07031_/A _07031_/B vssd1 vssd1 vccd1 vccd1 _07030_/A sky130_fd_sc_hd__or2_1
XANTENNA__09294__B _09389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _10045_/C _10040_/B _10049_/A vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__and3b_1
XANTENNA__10233__B _13758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11991_ _11991_/A vssd1 vssd1 vccd1 vccd1 _12922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _13730_/A _07016_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
X_10942_ _10942_/A _10942_/B _10942_/C _10942_/D vssd1 vssd1 vccd1 vccd1 _11328_/B
+ sky130_fd_sc_hd__or4_2
XANTENNA__06439__A _06913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ _13661_/A _07197_/X vssd1 vssd1 vccd1 vccd1 _14077_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10873_ _10862_/Y _10860_/C _10872_/X _10895_/A vssd1 vssd1 vccd1 vccd1 _12643_/D
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__13560__A _13560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12802_/CLK _12612_/D vssd1 vssd1 vccd1 vccd1 _13787_/A sky130_fd_sc_hd__dfxtp_2
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _13592_/A _07387_/X vssd1 vssd1 vccd1 vccd1 _14104_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_12_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12543_ _12565_/CLK _12543_/D vssd1 vssd1 vccd1 vccd1 _12543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09469__B _13551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09480__A1 _13570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11080__A _11206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12474_ _12656_/CLK _12474_/D vssd1 vssd1 vccd1 vccd1 _12474_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_91_clk_A _12438_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ _11438_/A vssd1 vssd1 vccd1 vccd1 _11425_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08666__S0 _08575_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11356_ _13911_/A _12768_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _11357_/B sky130_fd_sc_hd__mux2_1
XANTENNA__06902__A _07328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10307_ _13650_/A _12504_/Q _10375_/B vssd1 vssd1 vccd1 vccd1 _10308_/B sky130_fd_sc_hd__mux2_1
X_14075_ _14075_/A _08026_/X vssd1 vssd1 vccd1 vccd1 _14075_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10424__A _10667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11287_ _13871_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11287_/X sky130_fd_sc_hd__or2_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _12476_/Q _13751_/A vssd1 vssd1 vccd1 vccd1 _10242_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08969__S1 _08968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10169_ _13615_/A _12468_/Q _10180_/S vssd1 vssd1 vccd1 vccd1 _10170_/B sky130_fd_sc_hd__mux2_1
XFILLER_121_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13928_ _13928_/A _06480_/X vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_35_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13859_ _13859_/A _06672_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[20] sky130_fd_sc_hd__ebufn_8
XANTENNA_clkbuf_leaf_44_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06400_ _06403_/A _06400_/B vssd1 vssd1 vccd1 vccd1 _06401_/A sky130_fd_sc_hd__or2_1
XANTENNA__13470__A _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07380_ _07382_/A _07391_/B _07388_/C vssd1 vssd1 vccd1 vccd1 _07381_/A sky130_fd_sc_hd__or3_1
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11802__A0 _09623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06331_ _06333_/A _06336_/B _06336_/C vssd1 vssd1 vccd1 vccd1 _06332_/A sky130_fd_sc_hd__or3_1
X_09050_ _08970_/X _08972_/X _08975_/X _08976_/X _08952_/X _08953_/X vssd1 vssd1 vccd1
+ vccd1 _09050_/X sky130_fd_sc_hd__mux4_1
X_06262_ input24/X input23/X input3/X input2/X vssd1 vssd1 vccd1 vccd1 _06263_/D sky130_fd_sc_hd__or4_1
XFILLER_129_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_59_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08001_ _08001_/A vssd1 vssd1 vccd1 vccd1 _08001_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09395__A _09846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09952_ _09952_/A vssd1 vssd1 vccd1 vccd1 _12415_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10334__A _10988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ _10165_/C vssd1 vssd1 vccd1 vccd1 _13757_/A sky130_fd_sc_hd__buf_4
XFILLER_131_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater94_A _14121_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_117_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09750_/X _09874_/X _09882_/X _09878_/X vssd1 vssd1 vccd1 vccd1 _12393_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08834_ _08754_/X _08757_/X _08756_/X _08833_/X _08876_/A _08831_/X vssd1 vssd1 vccd1
+ vccd1 _08834_/X sky130_fd_sc_hd__mux4_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07643__A _08022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08765_ _12623_/Q _12624_/Q _12625_/Q _12626_/Q _08745_/X _08746_/X vssd1 vssd1 vccd1
+ vccd1 _08765_/X sky130_fd_sc_hd__mux4_2
XFILLER_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _07729_/A vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ _08628_/X _08631_/X _08637_/X _08640_/X _08694_/X _08695_/X vssd1 vssd1 vccd1
+ vccd1 _08696_/X sky130_fd_sc_hd__mux4_1
X_07647_ _07659_/A _07654_/B _07649_/C vssd1 vssd1 vccd1 vccd1 _07648_/A sky130_fd_sc_hd__or3_1
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07578_ _07588_/A _07585_/B _07580_/C vssd1 vssd1 vccd1 vccd1 _07579_/A sky130_fd_sc_hd__or3_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09317_ _09317_/A _09317_/B _09317_/C _09317_/D vssd1 vssd1 vccd1 vccd1 _09318_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_139_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06529_ _07507_/A vssd1 vssd1 vccd1 vccd1 _06540_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__10509__A _12062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ _09271_/C vssd1 vssd1 vccd1 vccd1 _09248_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10228__B _13753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_10_0_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _12759_/CLK sky130_fd_sc_hd__clkbuf_2
X_09179_ _13400_/A _09179_/B vssd1 vssd1 vccd1 vccd1 _09179_/X sky130_fd_sc_hd__and2_1
XFILLER_135_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11210_ _13873_/A _12729_/Q _11281_/B vssd1 vssd1 vccd1 vccd1 _11211_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07818__A _07868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12190_ _10648_/A _12182_/X _12189_/X _12187_/X vssd1 vssd1 vccd1 vccd1 _12973_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06722__A _06722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11141_ _12706_/Q _13947_/A vssd1 vssd1 vccd1 vccd1 _11143_/C sky130_fd_sc_hd__xor2_1
Xoutput33 _13979_/A vssd1 vssd1 vccd1 vccd1 pwm_en[14] sky130_fd_sc_hd__buf_2
Xoutput44 _13375_/A vssd1 vssd1 vccd1 vccd1 pwm_out[0] sky130_fd_sc_hd__buf_2
XFILLER_150_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput55 _13568_/A vssd1 vssd1 vccd1 vccd1 pwm_out[5] sky130_fd_sc_hd__buf_2
X_11072_ _13979_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11124_/S sky130_fd_sc_hd__and2_4
XFILLER_1_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10023_ _10024_/B _10024_/C _10022_/Y _09987_/X vssd1 vssd1 vccd1 vccd1 _12434_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13555__A _13555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07553__A _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A peripheralBus_address[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11974_ _14109_/Z _14045_/A _11974_/S vssd1 vssd1 vccd1 vccd1 _11975_/B sky130_fd_sc_hd__mux2_1
XFILLER_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13713_ _13713_/A _07056_/X vssd1 vssd1 vccd1 vccd1 _14097_/Z sky130_fd_sc_hd__ebufn_8
X_10925_ _10928_/B _10928_/C vssd1 vssd1 vccd1 vccd1 _10927_/A sky130_fd_sc_hd__and2_1
X_13644_ _13644_/A _07243_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
X_10856_ _10859_/B _10917_/B _10856_/C vssd1 vssd1 vccd1 vccd1 _10857_/A sky130_fd_sc_hd__and3b_1
XFILLER_32_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09199__B _09380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13575_ _13575_/A _07431_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10794_/C _10812_/B _10787_/C vssd1 vssd1 vccd1 vccd1 _10788_/A sky130_fd_sc_hd__and3b_1
XFILLER_40_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12526_ _12533_/CLK _12526_/D vssd1 vssd1 vccd1 vccd1 _13655_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12457_ _12457_/CLK _12457_/D vssd1 vssd1 vccd1 vccd1 _12457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11408_ _11408_/A _11408_/B _11408_/C vssd1 vssd1 vccd1 vccd1 _11409_/A sky130_fd_sc_hd__and3_1
X_12388_ _12414_/CLK _12388_/D vssd1 vssd1 vccd1 vccd1 _12388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06632__A _06680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11339_ _13906_/A _12763_/Q _11408_/B vssd1 vssd1 vccd1 vccd1 _11340_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12987__143 vssd1 vssd1 vccd1 vccd1 _12987__143/HI _13384_/A sky130_fd_sc_hd__conb_1
XFILLER_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09943__A _11490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ _14058_/A _07937_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06880_ _06890_/A _06884_/B _06884_/C vssd1 vssd1 vccd1 vccd1 _06881_/A sky130_fd_sc_hd__or3_1
XFILLER_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08550_ _13585_/A vssd1 vssd1 vccd1 vccd1 _08709_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07501_ _07501_/A vssd1 vssd1 vccd1 vccd1 _07501_/X sky130_fd_sc_hd__clkbuf_1
X_08481_ _12263_/Q vssd1 vssd1 vccd1 vccd1 _09362_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_63_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07432_ _07468_/A vssd1 vssd1 vccd1 vccd1 _07442_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_149_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13172__328 vssd1 vssd1 vccd1 vccd1 _13172__328/HI _13765_/A sky130_fd_sc_hd__conb_1
XFILLER_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ _07403_/A vssd1 vssd1 vccd1 vccd1 _07374_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09102_ _09102_/A _12062_/A _12059_/B _12062_/B vssd1 vssd1 vccd1 vccd1 _12208_/B
+ sky130_fd_sc_hd__nor4_2
X_06314_ _06320_/A _06323_/B _06323_/C vssd1 vssd1 vccd1 vccd1 _06315_/A sky130_fd_sc_hd__or3_1
X_07294_ _07533_/A vssd1 vssd1 vccd1 vccd1 _07519_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09033_ _12843_/Q vssd1 vssd1 vccd1 vccd1 _11677_/A sky130_fd_sc_hd__clkbuf_1
X_13213__369 vssd1 vssd1 vccd1 vccd1 _13213__369/HI _13836_/A sky130_fd_sc_hd__conb_1
XFILLER_117_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06542__A _06694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13066__222 vssd1 vssd1 vccd1 vccd1 _13066__222/HI _13541_/A sky130_fd_sc_hd__conb_1
X_09935_ _09939_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__or2_1
XANTENNA__13375__A _13375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _12382_/Q _13559_/A vssd1 vssd1 vccd1 vccd1 _09868_/C sky130_fd_sc_hd__xor2_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08802__S0 _08733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08817_ _12639_/Q vssd1 vssd1 vccd1 vccd1 _10875_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13107__263 vssd1 vssd1 vccd1 vccd1 _13107__263/HI _13632_/A sky130_fd_sc_hd__conb_1
XFILLER_100_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09797_ _09800_/A _09797_/B vssd1 vssd1 vccd1 vccd1 _09798_/A sky130_fd_sc_hd__and2_1
XFILLER_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _13778_/A vssd1 vssd1 vccd1 vccd1 _08748_/X sky130_fd_sc_hd__buf_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _08558_/X _08561_/X _08565_/X _08566_/X _08678_/X _08584_/X vssd1 vssd1 vccd1
+ vccd1 _08679_/X sky130_fd_sc_hd__mux4_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11623__A _11703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10710_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10710_/X sky130_fd_sc_hd__or2_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11703_/A _11690_/B _11690_/C vssd1 vssd1 vccd1 vccd1 _11691_/A sky130_fd_sc_hd__and3_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10641_ _13711_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10641_/X sky130_fd_sc_hd__or2_1
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13360_ _13360_/A _08280_/X vssd1 vssd1 vccd1 vccd1 _14096_/Z sky130_fd_sc_hd__ebufn_8
X_10572_ _13715_/A _12571_/Q _10584_/S vssd1 vssd1 vccd1 vccd1 _10573_/B sky130_fd_sc_hd__mux2_1
X_12311_ _12334_/CLK _12311_/D vssd1 vssd1 vccd1 vccd1 _12311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07548__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ _12242_/CLK _12242_/D vssd1 vssd1 vccd1 vccd1 _12242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12173__B _13367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12173_ _12961_/Q _13367_/A vssd1 vssd1 vccd1 vccd1 _12176_/B sky130_fd_sc_hd__xor2_1
XFILLER_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11124_ _13854_/A _12709_/Q _11124_/S vssd1 vssd1 vccd1 vccd1 _11125_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09763__A _10659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09046__S0 _08967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11055_ _11055_/A vssd1 vssd1 vccd1 vccd1 _11055_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10702__A input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ _10029_/C _10004_/A _09994_/X vssd1 vssd1 vccd1 vccd1 _10007_/B sky130_fd_sc_hd__o21ai_1
XFILLER_92_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11957_ _09638_/A _14040_/A _11957_/S vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__mux2_1
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10908_ _10908_/A _10908_/B _10908_/C _10908_/D vssd1 vssd1 vccd1 vccd1 _10922_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11888_ _11888_/A vssd1 vssd1 vccd1 vccd1 _11927_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13627_ _13627_/A _07287_/X vssd1 vssd1 vccd1 vccd1 _14075_/Z sky130_fd_sc_hd__ebufn_8
X_10839_ _10869_/B _10833_/X _10838_/Y vssd1 vssd1 vccd1 vccd1 _12636_/D sky130_fd_sc_hd__a21oi_1
Xrepeater63 _13623_/Z vssd1 vssd1 vccd1 vccd1 _14103_/Z sky130_fd_sc_hd__buf_12
Xrepeater74 peripheralBus_data[5] vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__buf_12
XFILLER_158_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13558_ _13558_/A _07472_/X vssd1 vssd1 vccd1 vccd1 _14102_/Z sky130_fd_sc_hd__ebufn_8
Xrepeater85 _14065_/Z vssd1 vssd1 vccd1 vccd1 _14097_/Z sky130_fd_sc_hd__buf_12
XFILLER_146_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater96 _14120_/Z vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__buf_12
XFILLER_158_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12509_ _12515_/CLK _12509_/D vssd1 vssd1 vccd1 vccd1 _12509_/Q sky130_fd_sc_hd__dfxtp_1
X_13489_ _13489_/A _07653_/X vssd1 vssd1 vccd1 vccd1 _14033_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_126_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07981_ _08064_/A vssd1 vssd1 vccd1 vccd1 _08062_/B sky130_fd_sc_hd__buf_2
XFILLER_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09720_ _09715_/X _09716_/Y _09717_/Y _09718_/X _09719_/Y vssd1 vssd1 vccd1 vccd1
+ _09720_/X sky130_fd_sc_hd__o221a_1
X_06932_ _06936_/A _06941_/B vssd1 vssd1 vccd1 vccd1 _06933_/A sky130_fd_sc_hd__or2_1
XFILLER_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09651_ _11064_/A _09653_/B vssd1 vssd1 vccd1 vccd1 _09651_/X sky130_fd_sc_hd__or2_1
XFILLER_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06863_ _06863_/A _06870_/B _06870_/C vssd1 vssd1 vccd1 vccd1 _06864_/A sky130_fd_sc_hd__or3_1
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08602_ _08708_/A vssd1 vssd1 vccd1 vccd1 _08602_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09582_ _13470_/A _12323_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09583_/B sky130_fd_sc_hd__mux2_1
X_06794_ _06794_/A vssd1 vssd1 vccd1 vccd1 _06794_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08533_ _08411_/X _08475_/X _08502_/X _08532_/X _08511_/X _08517_/X vssd1 vssd1 vccd1
+ vccd1 _08533_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11443__A _11443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ _08450_/X _08462_/X _08528_/S vssd1 vssd1 vccd1 vccd1 _11706_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07415_ _07417_/A _07423_/B vssd1 vssd1 vccd1 vccd1 _07416_/A sky130_fd_sc_hd__or2_1
XFILLER_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08395_ _12229_/Q _12230_/Q _12231_/Q _12232_/Q _08368_/X _08370_/X vssd1 vssd1 vccd1
+ vccd1 _08395_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ _07346_/A vssd1 vssd1 vccd1 vccd1 _07346_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07277_ _07277_/A vssd1 vssd1 vccd1 vccd1 _07277_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09016_ _08931_/X _08932_/X _08933_/X _09015_/X _09030_/A _08934_/X vssd1 vssd1 vccd1
+ vccd1 _09016_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10735__A0 _10614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09918_ _11457_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09925_/A sky130_fd_sc_hd__nor2_2
XFILLER_120_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09849_ _12385_/Q _13562_/A vssd1 vssd1 vccd1 vccd1 _09849_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10241__B _13743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13341__497 vssd1 vssd1 vccd1 vccd1 _13341__497/HI _14094_/A sky130_fd_sc_hd__conb_1
XFILLER_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12860_ _12867_/CLK _12860_/D vssd1 vssd1 vccd1 vccd1 _12860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11811_/A vssd1 vssd1 vccd1 vccd1 _12876_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09656__A1 _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12791_ _12923_/CLK _12791_/D vssd1 vssd1 vccd1 vccd1 _13917_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11801_/A vssd1 vssd1 vccd1 vccd1 _11757_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13194__350 vssd1 vssd1 vccd1 vccd1 _13194__350/HI _13801_/A sky130_fd_sc_hd__conb_1
XANTENNA__12168__B _13374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11689_/A _11672_/X _11582_/C vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__a21bo_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13412_ _13412_/A _08173_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
X_10624_ _12579_/Q _13755_/A vssd1 vssd1 vccd1 vccd1 _10627_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13235__391 vssd1 vssd1 vccd1 vccd1 _13235__391/HI _13890_/A sky130_fd_sc_hd__conb_1
XFILLER_139_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09477__B _13558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10555_ _13785_/A _10555_/B vssd1 vssd1 vccd1 vccd1 _10608_/S sky130_fd_sc_hd__and2_2
XFILLER_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07278__A _07291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09196__C _09196_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10486_ _12535_/Q _10614_/B vssd1 vssd1 vccd1 vccd1 _10486_/X sky130_fd_sc_hd__and2_1
XFILLER_6_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12225_ _12969_/CLK _12225_/D vssd1 vssd1 vccd1 vccd1 _13402_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_108_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11923__C1 _09404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A _09967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ _12156_/A vssd1 vssd1 vccd1 vccd1 _12968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11107_ _11107_/A vssd1 vssd1 vccd1 vccd1 _12703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12087_ _10670_/A _12075_/X _12086_/X _12084_/X vssd1 vssd1 vccd1 vccd1 _12946_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_output54_A _13567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11038_ _13811_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11038_/X sky130_fd_sc_hd__or2_1
XFILLER_65_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09895__A1 _09763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10151__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13743__A _13743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07200_ _07206_/A _07203_/B _07200_/C vssd1 vssd1 vccd1 vccd1 _07201_/A sky130_fd_sc_hd__or3_1
XFILLER_165_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08180_ _08180_/A _08180_/B _08180_/C vssd1 vssd1 vccd1 vccd1 _08181_/A sky130_fd_sc_hd__or3_1
XFILLER_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07131_ _07135_/A _07131_/B _07142_/C vssd1 vssd1 vccd1 vccd1 _07132_/A sky130_fd_sc_hd__or3_1
XFILLER_118_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07062_ _07406_/A vssd1 vssd1 vccd1 vccd1 _08177_/A sky130_fd_sc_hd__buf_2
XFILLER_118_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06820__A _07248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07964_ _07964_/A vssd1 vssd1 vccd1 vccd1 _08075_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__12033__S _12033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09703_ _09703_/A vssd1 vssd1 vccd1 vccd1 _12353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06915_ _06915_/A vssd1 vssd1 vccd1 vccd1 _06915_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07895_ _07895_/A vssd1 vssd1 vccd1 vccd1 _07895_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09634_ _09634_/A vssd1 vssd1 vccd1 vccd1 _09634_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09850__B _13552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ _06900_/A vssd1 vssd1 vccd1 vccd1 _06857_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_83_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09565_ _09671_/A vssd1 vssd1 vccd1 vccd1 _09579_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13178__334 vssd1 vssd1 vccd1 vccd1 _13178__334/HI _13771_/A sky130_fd_sc_hd__conb_1
X_06777_ _06803_/A vssd1 vssd1 vccd1 vccd1 _06788_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_82_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08516_ _09368_/A _09377_/C _12269_/Q _09377_/A _08417_/X _08418_/X vssd1 vssd1 vccd1
+ vccd1 _08516_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11445__A1 _11189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ _09634_/A vssd1 vssd1 vccd1 vccd1 _09496_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__06267__A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08447_ _09316_/A _09322_/D _09328_/B _09321_/D _08445_/X _08446_/X vssd1 vssd1 vccd1
+ vccd1 _08447_/X sky130_fd_sc_hd__mux4_2
X_13219__375 vssd1 vssd1 vccd1 vccd1 _13219__375/HI _13858_/A sky130_fd_sc_hd__conb_1
XFILLER_23_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08378_ _12236_/Q _12237_/Q _12238_/Q _12239_/Q _08376_/X _08377_/X vssd1 vssd1 vccd1
+ vccd1 _08378_/X sky130_fd_sc_hd__mux4_2
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07329_ _07329_/A vssd1 vssd1 vccd1 vccd1 _07329_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10340_ _10349_/A _10340_/B vssd1 vssd1 vccd1 vccd1 _10341_/A sky130_fd_sc_hd__and2_1
XFILLER_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10236__B _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10271_ _09763_/X _10264_/X _10268_/X _10270_/X vssd1 vssd1 vccd1 vccd1 _12491_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12010_ _12013_/A _12010_/B vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__and2_1
XANTENNA__07826__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10252__A _10293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13961_ _13961_/A _06395_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[26] sky130_fd_sc_hd__ebufn_8
XFILLER_120_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13563__A _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ _12912_/CLK _12912_/D vssd1 vssd1 vccd1 vccd1 _14039_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892_ _13892_/A _06581_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[21] sky130_fd_sc_hd__ebufn_8
XANTENNA__08657__A _09867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07561__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ _12850_/CLK _12843_/D vssd1 vssd1 vccd1 vccd1 _12843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10892__C1 _10749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12938_/CLK _12774_/D vssd1 vssd1 vccd1 vccd1 _12774_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _11801_/A vssd1 vssd1 vccd1 vccd1 _11740_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09488__A _11160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11656_ _11661_/B _11661_/C _11569_/X vssd1 vssd1 vccd1 vccd1 _11659_/A sky130_fd_sc_hd__o21ai_1
X_10607_ _10607_/A vssd1 vssd1 vccd1 vccd1 _12581_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10427__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11587_ _11587_/A _11587_/B vssd1 vssd1 vccd1 vccd1 _12825_/D sky130_fd_sc_hd__nor2_1
XFILLER_127_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10538_ _10538_/A vssd1 vssd1 vccd1 vccd1 _10538_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10469_ _10469_/A vssd1 vssd1 vccd1 vccd1 _12545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13012__168 vssd1 vssd1 vccd1 vccd1 _13012__168/HI _13439_/A sky130_fd_sc_hd__conb_1
X_12208_ _14106_/A _12208_/B vssd1 vssd1 vccd1 vccd1 _12208_/X sky130_fd_sc_hd__or2_1
XANTENNA__06640__A _11156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11258__A _12740_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12139_ _12963_/Q _14105_/A _12151_/S vssd1 vssd1 vccd1 vccd1 _12140_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09951__A _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06700_ _06700_/A vssd1 vssd1 vccd1 vccd1 _06700_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07680_ _07693_/A vssd1 vssd1 vccd1 vccd1 _07691_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_53_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06631_ _06631_/A vssd1 vssd1 vccd1 vccd1 _06631_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09350_ _09350_/A vssd1 vssd1 vccd1 vccd1 _12262_/D sky130_fd_sc_hd__clkbuf_1
X_06562_ _06562_/A vssd1 vssd1 vccd1 vccd1 _06562_/X sky130_fd_sc_hd__clkbuf_1
X_08301_ _08301_/A vssd1 vssd1 vccd1 vccd1 _08301_/X sky130_fd_sc_hd__clkbuf_1
X_09281_ _09281_/A vssd1 vssd1 vccd1 vccd1 _09392_/A sky130_fd_sc_hd__buf_2
XFILLER_21_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06493_ _06493_/A vssd1 vssd1 vccd1 vccd1 _06493_/X sky130_fd_sc_hd__clkbuf_1
X_08232_ _08232_/A vssd1 vssd1 vccd1 vccd1 _08232_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06815__A _06983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ _08163_/A vssd1 vssd1 vccd1 vccd1 _08163_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07114_ _07114_/A vssd1 vssd1 vccd1 vccd1 _07114_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ _08153_/A vssd1 vssd1 vccd1 vccd1 _08105_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_119_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07045_ _07045_/A vssd1 vssd1 vccd1 vccd1 _07055_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_161_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06550__A _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08996_ _09057_/A vssd1 vssd1 vccd1 vccd1 _08996_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07947_ _08180_/A _07947_/B _08349_/B vssd1 vssd1 vccd1 vccd1 _07948_/A sky130_fd_sc_hd__or3_2
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07878_ _07878_/A vssd1 vssd1 vccd1 vccd1 _07878_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09617_ _13455_/A _09613_/X _09616_/X _09522_/X vssd1 vssd1 vccd1 vccd1 _12325_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06829_ _06829_/A vssd1 vssd1 vccd1 vccd1 _06829_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11418__A1 _11160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09548_ _09671_/A vssd1 vssd1 vccd1 vccd1 _09563_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12091__A1 _11184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ _09479_/A _09479_/B _09479_/C vssd1 vssd1 vccd1 vccd1 _09479_/X sky130_fd_sc_hd__and3_1
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11510_ _11520_/A vssd1 vssd1 vccd1 vccd1 _11576_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12490_ _12492_/CLK _12490_/D vssd1 vssd1 vccd1 vccd1 _13620_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11441_ _11184_/X _11438_/X _11440_/X _11430_/X vssd1 vssd1 vccd1 vccd1 _12787_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10247__A _10688_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11372_ _11372_/A vssd1 vssd1 vccd1 vccd1 _12772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13558__A _13558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10323_ _10323_/A vssd1 vssd1 vccd1 vccd1 _12508_/D sky130_fd_sc_hd__clkbuf_1
X_14091_ _14091_/A _08149_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
XFILLER_124_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10254_ _09124_/X _10249_/X _10253_/X _09959_/X vssd1 vssd1 vccd1 vccd1 _12485_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06460__A _07822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10185_ _10191_/A _10185_/B vssd1 vssd1 vccd1 vccd1 _10186_/A sky130_fd_sc_hd__and2_1
XFILLER_120_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08770__A1 _08764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__A _13495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13944_ _13944_/A _06436_/X vssd1 vssd1 vccd1 vccd1 _13976_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07291__A _07291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13875_ _13875_/A _06626_/X vssd1 vssd1 vccd1 vccd1 _14067_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12826_ _12829_/CLK _12826_/D vssd1 vssd1 vccd1 vccd1 _12826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12757_ _12758_/CLK _12757_/D vssd1 vssd1 vccd1 vccd1 _13884_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12082__A1 _10662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11708_/A _11708_/B _11708_/C _11708_/D vssd1 vssd1 vccd1 vccd1 _11709_/D
+ sky130_fd_sc_hd__or4_1
X_12688_ _12710_/CLK _12688_/D vssd1 vssd1 vccd1 vccd1 _13817_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11260__B _13936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11639_ _11639_/A _11639_/B _11639_/C vssd1 vssd1 vccd1 vccd1 _11642_/B sky130_fd_sc_hd__and3_1
XFILLER_162_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_3_clk_A _12917_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08850_ _08850_/A vssd1 vssd1 vccd1 vccd1 _08850_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07801_ _07809_/A _07806_/B _07801_/C vssd1 vssd1 vccd1 vccd1 _07802_/A sky130_fd_sc_hd__or3_1
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08781_ _10806_/B _12617_/Q _10773_/D _12619_/Q _08779_/X _08780_/X vssd1 vssd1 vccd1
+ vccd1 _08781_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07732_ _07742_/A _07737_/B _07732_/C vssd1 vssd1 vccd1 vccd1 _07733_/A sky130_fd_sc_hd__or3_1
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08513__A1 _08447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07663_ _07663_/A vssd1 vssd1 vccd1 vccd1 _07663_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09402_ _09454_/S vssd1 vssd1 vccd1 vccd1 _09414_/S sky130_fd_sc_hd__clkbuf_2
X_06614_ _06625_/A _06616_/B _06616_/C vssd1 vssd1 vccd1 vccd1 _06615_/A sky130_fd_sc_hd__or3_1
X_13140__296 vssd1 vssd1 vccd1 vccd1 _13140__296/HI _13697_/A sky130_fd_sc_hd__conb_1
XANTENNA__12058__D1 _13402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11154__C _11410_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07594_ _07594_/A vssd1 vssd1 vccd1 vccd1 _07594_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ _09336_/A _09324_/X _09332_/Y _09263_/X vssd1 vssd1 vccd1 vccd1 _12258_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06545_ _06556_/A _06561_/B _08180_/B vssd1 vssd1 vccd1 vccd1 _06546_/A sky130_fd_sc_hd__or3_1
XFILLER_139_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09264_ _09316_/A _09257_/B _09262_/Y _09263_/X vssd1 vssd1 vccd1 vccd1 _12243_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11820__A1 _14007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06476_ _08276_/B vssd1 vssd1 vccd1 vccd1 _06486_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_21_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08215_ _08228_/A vssd1 vssd1 vccd1 vccd1 _08225_/C sky130_fd_sc_hd__clkbuf_1
X_09195_ _13400_/A _13399_/A _09194_/X vssd1 vssd1 vccd1 vccd1 _09196_/C sky130_fd_sc_hd__or3b_2
XANTENNA__06264__B _09096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ _08148_/A _08151_/B _08151_/C vssd1 vssd1 vccd1 vccd1 _08147_/A sky130_fd_sc_hd__or3_1
XFILLER_20_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10387__A1 _10385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13378__A _13378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034__190 vssd1 vssd1 vccd1 vccd1 _13034__190/HI _13477_/A sky130_fd_sc_hd__conb_1
XFILLER_107_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08077_ _08081_/A _08077_/B _08087_/C vssd1 vssd1 vccd1 vccd1 _08078_/A sky130_fd_sc_hd__or3_1
XFILLER_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07376__A _07403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07028_ _07028_/A vssd1 vssd1 vccd1 vccd1 _07028_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06280__A _06442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08979_ _12838_/Q vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11990_ _11996_/A _11990_/B vssd1 vssd1 vccd1 vccd1 _11991_/A sky130_fd_sc_hd__and2_1
XFILLER_17_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10941_ _10941_/A _10941_/B _10941_/C _10941_/D vssd1 vssd1 vccd1 vccd1 _10942_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_45_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13660_ _13660_/A _07199_/X vssd1 vssd1 vccd1 vccd1 _14108_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_32_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10872_ _10872_/A _10881_/B _10881_/C vssd1 vssd1 vccd1 vccd1 _10872_/X sky130_fd_sc_hd__and3_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _12802_/CLK _12611_/D vssd1 vssd1 vccd1 vccd1 _13786_/A sky130_fd_sc_hd__dfxtp_2
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_117_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _12258_/CLK sky130_fd_sc_hd__clkbuf_16
X_13591_ _13591_/A _07389_/X vssd1 vssd1 vccd1 vccd1 _13623_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_40_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12542_ _12554_/CLK _12542_/D vssd1 vssd1 vccd1 vccd1 _12542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06455__A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12473_ _12659_/CLK _12473_/D vssd1 vssd1 vccd1 vccd1 _12473_/Q sky130_fd_sc_hd__dfxtp_1
X_11424_ _10652_/X _11411_/X _11423_/X _11417_/X vssd1 vssd1 vccd1 vccd1 _12781_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08666__S1 _08576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ _11355_/A vssd1 vssd1 vccd1 vccd1 _12767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06902__B _07336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ _10306_/A vssd1 vssd1 vccd1 vccd1 _12503_/D sky130_fd_sc_hd__clkbuf_1
X_14074_ _14074_/A _08024_/X vssd1 vssd1 vccd1 vccd1 _14106_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_3_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11286_ _11325_/B vssd1 vssd1 vccd1 vccd1 _11297_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_140_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10237_ _10237_/A _10237_/B _10237_/C _10237_/D vssd1 vssd1 vccd1 vccd1 _10243_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13083__239 vssd1 vssd1 vccd1 vccd1 _13083__239/HI _13578_/A sky130_fd_sc_hd__conb_1
XFILLER_126_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10168_ _10220_/S vssd1 vssd1 vccd1 vccd1 _10180_/S sky130_fd_sc_hd__buf_2
XFILLER_66_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10099_ _10099_/A _10099_/B _10099_/C _10099_/D vssd1 vssd1 vccd1 vccd1 _10100_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13927_ _13927_/A _06482_/X vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13751__A _13751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _13858_/A _06674_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
XFILLER_35_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12809_ _12811_/CLK _12809_/D vssd1 vssd1 vccd1 vccd1 _12809_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_108_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _12334_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13789_ _13789_/A _06867_/X vssd1 vssd1 vccd1 vccd1 _14077_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06330_ _06330_/A vssd1 vssd1 vccd1 vccd1 _06330_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06261_ input17/X vssd1 vssd1 vccd1 vccd1 _09102_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08000_ _08010_/A _08005_/B _08002_/C vssd1 vssd1 vccd1 vccd1 _08001_/A sky130_fd_sc_hd__or3_1
XFILLER_163_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13018__174 vssd1 vssd1 vccd1 vccd1 _13018__174/HI _13445_/A sky130_fd_sc_hd__conb_1
XFILLER_129_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09951_ _10700_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__or2_1
XANTENNA__11581__A3 _11649_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ _08898_/X _08901_/X _10710_/A vssd1 vssd1 vccd1 vccd1 _10165_/C sky130_fd_sc_hd__mux2_1
XFILLER_103_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _13521_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09882_/X sky130_fd_sc_hd__or2_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09931__A0 _14033_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater87_A peripheralBus_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08833_ _12646_/Q _12647_/Q _12648_/Q _12649_/Q _08785_/X _08786_/X vssd1 vssd1 vccd1
+ vccd1 _08833_/X sky130_fd_sc_hd__mux4_1
XANTENNA__07924__A _07999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10541__A1 _10408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08764_ _12619_/Q _12620_/Q _12621_/Q _12622_/Q _08745_/X _08746_/X vssd1 vssd1 vccd1
+ vccd1 _08764_/X sky130_fd_sc_hd__mux4_2
XFILLER_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ _07715_/A vssd1 vssd1 vccd1 vccd1 _07715_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _08695_/A vssd1 vssd1 vccd1 vccd1 _08695_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07646_ _07661_/A vssd1 vssd1 vccd1 vccd1 _07659_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_81_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07577_ _07590_/A vssd1 vssd1 vccd1 vccd1 _07588_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09316_ _09316_/A _09316_/B _09316_/C _09316_/D vssd1 vssd1 vccd1 vccd1 _09318_/C
+ sky130_fd_sc_hd__and4_1
X_06528_ _06528_/A vssd1 vssd1 vccd1 vccd1 _06540_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_139_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09247_ _12240_/Q vssd1 vssd1 vccd1 vccd1 _09315_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06459_ _08276_/B vssd1 vssd1 vccd1 vccd1 _06472_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_21_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09178_ _09638_/A vssd1 vssd1 vccd1 vccd1 _10670_/A sky130_fd_sc_hd__buf_4
XFILLER_5_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ _08129_/A vssd1 vssd1 vccd1 vccd1 _08129_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ _12709_/Q _13950_/A vssd1 vssd1 vccd1 vccd1 _11143_/B sky130_fd_sc_hd__xor2_1
Xoutput34 _13980_/A vssd1 vssd1 vccd1 vccd1 pwm_en[15] sky130_fd_sc_hd__buf_2
XFILLER_162_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput45 _13761_/A vssd1 vssd1 vccd1 vccd1 pwm_out[10] sky130_fd_sc_hd__buf_2
XFILLER_163_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput56 _13569_/A vssd1 vssd1 vccd1 vccd1 pwm_out[6] sky130_fd_sc_hd__buf_2
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11071_ _10552_/X _11055_/A _11070_/X _11068_/X vssd1 vssd1 vccd1 vccd1 _12693_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10022_ _10022_/A _10030_/C vssd1 vssd1 vccd1 vccd1 _10022_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10532__A1 _09767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input16_A peripheralBus_address[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08489__A0 _08455_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _11973_/A vssd1 vssd1 vccd1 vccd1 _12917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10924_ _10872_/A _10928_/C _10923_/Y _10895_/A vssd1 vssd1 vccd1 vccd1 _12656_/D
+ sky130_fd_sc_hd__a211oi_1
X_13712_ _13712_/A _07058_/X vssd1 vssd1 vccd1 vccd1 _14064_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__12438__CLK _12438_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13643_ _13643_/A _07245_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
X_10855_ _10868_/D _10854_/C _10876_/A vssd1 vssd1 vccd1 vccd1 _10856_/C sky130_fd_sc_hd__a21o_1
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12187__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13574_ _13574_/A _07434_/X vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10786_ _10865_/B _10790_/C vssd1 vssd1 vccd1 vccd1 _10787_/C sky130_fd_sc_hd__or2_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ _12583_/CLK _12525_/D vssd1 vssd1 vccd1 vccd1 _13654_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09496__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ _12457_/CLK _12456_/D vssd1 vssd1 vccd1 vccd1 _12456_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06913__A _06913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ _11384_/Y _11390_/X _11406_/Y _13951_/A vssd1 vssd1 vccd1 vccd1 _11408_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12387_ _12400_/CLK _12387_/D vssd1 vssd1 vccd1 vccd1 _12387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14126_ _14126_/A _08277_/X vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__ebufn_8
X_11338_ _11338_/A vssd1 vssd1 vccd1 vccd1 _12762_/D sky130_fd_sc_hd__clkbuf_1
X_14057_ _14057_/A _07932_/X vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__13746__A _13746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ _12734_/Q _13942_/A vssd1 vssd1 vccd1 vccd1 _11273_/A sky130_fd_sc_hd__xor2_1
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07744__A _07923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10170__A _10173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ _07504_/A _07504_/B _07510_/C vssd1 vssd1 vccd1 vccd1 _07501_/A sky130_fd_sc_hd__or3_1
X_08480_ _08420_/X _08423_/X _08421_/X _08427_/X _08470_/X _09152_/A vssd1 vssd1 vccd1
+ vccd1 _08480_/X sky130_fd_sc_hd__mux4_1
X_07431_ _07431_/A vssd1 vssd1 vccd1 vccd1 _07431_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__12097__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07362_ _07362_/A vssd1 vssd1 vccd1 vccd1 _07362_/X sky130_fd_sc_hd__clkbuf_1
X_09101_ _10250_/A vssd1 vssd1 vccd1 vccd1 _12062_/A sky130_fd_sc_hd__clkbuf_4
X_06313_ _07045_/A vssd1 vssd1 vccd1 vccd1 _06323_/C sky130_fd_sc_hd__clkbuf_1
X_07293_ _07293_/A vssd1 vssd1 vccd1 vccd1 _07293_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06281__B_N input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09032_ _12842_/Q vssd1 vssd1 vccd1 vccd1 _11677_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07919__A _11154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09934_ _14034_/Z _08670_/X _09934_/S vssd1 vssd1 vccd1 vccd1 _09935_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10999__B _13944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09865_ _12379_/Q _13556_/A vssd1 vssd1 vccd1 vccd1 _09868_/B sky130_fd_sc_hd__xor2_1
XANTENNA_input8_A peripheralBus_address[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08802__S1 _08735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08816_ _12637_/Q vssd1 vssd1 vccd1 vccd1 _10876_/C sky130_fd_sc_hd__clkbuf_1
X_09796_ _13520_/A _12375_/Q _09871_/B vssd1 vssd1 vccd1 vccd1 _09797_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_90_clk_A _12438_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08747_ _12626_/Q _12627_/Q _12628_/Q _12629_/Q _08745_/X _08746_/X vssd1 vssd1 vccd1
+ vccd1 _08747_/X sky130_fd_sc_hd__mux4_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08566__S0 _08559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13391__A _13391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _13586_/A vssd1 vssd1 vccd1 vccd1 _08678_/X sky130_fd_sc_hd__buf_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08486__A3 _08452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07629_ _08022_/A vssd1 vssd1 vccd1 vccd1 _07641_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07820__C _08110_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10686_/B vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10239__B _13747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10571_ _10608_/S vssd1 vssd1 vccd1 vccd1 _10584_/S sky130_fd_sc_hd__clkbuf_2
X_12310_ _12320_/CLK _12310_/D vssd1 vssd1 vccd1 vccd1 _12310_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07829__A _07964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12241_ _12242_/CLK _12241_/D vssd1 vssd1 vccd1 vccd1 _12241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13346__502 vssd1 vssd1 vccd1 vccd1 _13346__502/HI _14115_/A sky130_fd_sc_hd__conb_1
XFILLER_135_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12172_ _12958_/Q _13364_/A vssd1 vssd1 vccd1 vccd1 _12176_/A sky130_fd_sc_hd__xor2_1
XFILLER_162_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ _11123_/A vssd1 vssd1 vccd1 vccd1 _12708_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13566__A _13566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_43_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09046__S1 _08968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11054_ _10670_/X _11041_/X _11051_/X _11053_/X vssd1 vssd1 vccd1 vccd1 _12687_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09482__C _10637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09371__A1 _09347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _10029_/C _10029_/D _10008_/D vssd1 vssd1 vccd1 vccd1 _10022_/A sky130_fd_sc_hd__and3_1
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_58_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_101_clk_A _12555_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11956_ _11956_/A vssd1 vssd1 vccd1 vccd1 _12912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ _10907_/A _10907_/B _10907_/C _10907_/D vssd1 vssd1 vccd1 vccd1 _10908_/D
+ sky130_fd_sc_hd__and4_1
X_11887_ _11887_/A vssd1 vssd1 vccd1 vccd1 _12898_/D sky130_fd_sc_hd__clkbuf_1
X_13626_ _13626_/A _07290_/X vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_8
X_10838_ _10869_/B _10833_/X _10803_/X vssd1 vssd1 vccd1 vccd1 _10838_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_116_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater64 peripheralBus_data[8] vssd1 vssd1 vccd1 vccd1 _13623_/Z sky130_fd_sc_hd__buf_12
Xrepeater75 _14067_/Z vssd1 vssd1 vccd1 vccd1 _14099_/Z sky130_fd_sc_hd__buf_12
X_13557_ _13557_/A _07475_/X vssd1 vssd1 vccd1 vccd1 _14037_/Z sky130_fd_sc_hd__ebufn_8
Xrepeater86 _14033_/Z vssd1 vssd1 vccd1 vccd1 _14065_/Z sky130_fd_sc_hd__buf_12
X_10769_ _10864_/D _10767_/C _10864_/C vssd1 vssd1 vccd1 vccd1 _10770_/C sky130_fd_sc_hd__a21o_1
XFILLER_157_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater97 peripheralBus_data[25] vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__buf_12
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12508_ _12515_/CLK _12508_/D vssd1 vssd1 vccd1 vccd1 _12508_/Q sky130_fd_sc_hd__dfxtp_1
X_13488_ _13488_/A _07655_/X vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_157_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12439_ _12443_/CLK _12439_/D vssd1 vssd1 vccd1 vccd1 _12439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13089__245 vssd1 vssd1 vccd1 vccd1 _13089__245/HI _13598_/A sky130_fd_sc_hd__conb_1
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09954__A _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14109_ _14109_/A _08234_/X vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__ebufn_8
X_07980_ _07980_/A vssd1 vssd1 vccd1 vccd1 _07980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06931_ _06955_/A vssd1 vssd1 vccd1 vccd1 _06941_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_68_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10612__B _13754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _13467_/A _09640_/X _09646_/X _09649_/X vssd1 vssd1 vccd1 vccd1 _12337_/D
+ sky130_fd_sc_hd__o211a_1
X_06862_ _06862_/A vssd1 vssd1 vccd1 vccd1 _06862_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08601_ _12423_/Q vssd1 vssd1 vccd1 vccd1 _09981_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09581_ _09671_/A vssd1 vssd1 vccd1 vccd1 _09669_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06793_ _06801_/A _06793_/B _06793_/C vssd1 vssd1 vccd1 vccd1 _06794_/A sky130_fd_sc_hd__or3_1
XFILLER_82_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09114__A1 _09112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08532_ _09377_/B _12270_/Q _12271_/Q _12272_/Q _09140_/A _09146_/A vssd1 vssd1 vccd1
+ vccd1 _08532_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08463_ _13396_/A vssd1 vssd1 vccd1 vccd1 _08528_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07414_ _07414_/A vssd1 vssd1 vccd1 vccd1 _07414_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08394_ _11706_/A vssd1 vssd1 vccd1 vccd1 _13359_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07345_ _07356_/A _07351_/B _07347_/C vssd1 vssd1 vccd1 vccd1 _07346_/A sky130_fd_sc_hd__or3_1
XANTENNA__09848__B _09848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_clk _12759_/CLK vssd1 vssd1 vccd1 vccd1 _12768_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08720__S0 _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07276_ _07279_/A _07276_/B _07286_/C vssd1 vssd1 vccd1 vccd1 _07277_/A sky130_fd_sc_hd__or3_1
X_09015_ _12839_/Q _12840_/Q _12841_/Q _12842_/Q _08915_/X _08916_/X vssd1 vssd1 vccd1
+ vccd1 _09015_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07384__A _09125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__B _11682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ _09120_/X _09902_/A _09915_/X _09916_/X vssd1 vssd1 vccd1 vccd1 _12406_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_97_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _12349_/CLK sky130_fd_sc_hd__clkbuf_16
X_09848_ _12385_/Q _09848_/B vssd1 vssd1 vccd1 vccd1 _09848_/X sky130_fd_sc_hd__and2_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09779_ _09182_/X _09776_/X _09778_/X _09765_/X vssd1 vssd1 vccd1 vccd1 _12368_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11634__A _11634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11810_ _11816_/A _11810_/B vssd1 vssd1 vccd1 vccd1 _11811_/A sky130_fd_sc_hd__and2_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12938_/CLK _12790_/D vssd1 vssd1 vccd1 vccd1 _13916_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09656__A2 _09640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11741_/A vssd1 vssd1 vccd1 vccd1 _12862_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11672_ _11672_/A _11676_/C _11672_/C vssd1 vssd1 vccd1 vccd1 _11672_/X sky130_fd_sc_hd__and3_1
XFILLER_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _12582_/Q _13758_/A vssd1 vssd1 vccd1 vccd1 _10627_/A sky130_fd_sc_hd__xor2_1
X_13411_ _13411_/A _08163_/X vssd1 vssd1 vccd1 vccd1 _13987_/Z sky130_fd_sc_hd__ebufn_8
Xclkbuf_leaf_21_clk _12881_/CLK vssd1 vssd1 vccd1 vccd1 _12935_/CLK sky130_fd_sc_hd__clkbuf_16
X_10554_ _10552_/X _10538_/A _10553_/X _10550_/X vssd1 vssd1 vccd1 vccd1 _12566_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06463__A _06547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10485_ _12545_/Q _10613_/B vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__and2_1
X_12224_ _12969_/CLK _12224_/D vssd1 vssd1 vccd1 vccd1 _13401_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ _12155_/A _12155_/B vssd1 vssd1 vccd1 vccd1 _12156_/A sky130_fd_sc_hd__and2_1
XANTENNA_repeater118_A peripheralBus_data[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ _11112_/A _11106_/B vssd1 vssd1 vccd1 vccd1 _11107_/A sky130_fd_sc_hd__and2_1
XFILLER_150_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07294__A _07533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12086_ _14072_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12086_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_88_clk _12438_/CLK vssd1 vssd1 vccd1 vccd1 _12457_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11037_ _10648_/X _11027_/X _11036_/X _11024_/X vssd1 vssd1 vccd1 vccd1 _12681_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output47_A _13951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06638__A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11939_ _11939_/A vssd1 vssd1 vccd1 vccd1 _12907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ _13609_/A _07341_/X vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_119_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_clk _12217_/CLK vssd1 vssd1 vccd1 vccd1 _12903_/CLK sky130_fd_sc_hd__clkbuf_16
X_07130_ _07162_/A vssd1 vssd1 vccd1 vccd1 _07142_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__06373__A _11457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07061_ _07061_/A vssd1 vssd1 vccd1 vccd1 _07061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09341__C_N _09263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07963_ _07963_/A vssd1 vssd1 vccd1 vccd1 _07963_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _12646_/CLK sky130_fd_sc_hd__clkbuf_16
X_09702_ _09705_/A _09702_/B vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__and2_1
X_06914_ _06923_/A _06916_/B vssd1 vssd1 vccd1 vccd1 _06915_/A sky130_fd_sc_hd__or2_1
X_07894_ _07894_/A _07903_/B _07903_/C vssd1 vssd1 vccd1 vccd1 _07895_/A sky130_fd_sc_hd__or3_1
XFILLER_67_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09633_ _09633_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09633_/X sky130_fd_sc_hd__or2_1
XFILLER_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06845_ _07406_/A vssd1 vssd1 vccd1 vccd1 _06900_/A sky130_fd_sc_hd__buf_2
XANTENNA__11454__A _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _09564_/A vssd1 vssd1 vccd1 vccd1 _12317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06776_ _06776_/A vssd1 vssd1 vccd1 vccd1 _06776_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ _12270_/Q vssd1 vssd1 vccd1 vccd1 _09377_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09495_ _12134_/A vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__buf_2
X_08446_ _08525_/A vssd1 vssd1 vccd1 vccd1 _08446_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08377_ _13393_/A vssd1 vssd1 vccd1 vccd1 _08377_/X sky130_fd_sc_hd__buf_2
XANTENNA__11901__B _13368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07379__A _07393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07328_ _07328_/A _07336_/B _07739_/C vssd1 vssd1 vccd1 vccd1 _07329_/A sky130_fd_sc_hd__or3_1
XFILLER_139_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06283__A _08186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07259_ _07259_/A vssd1 vssd1 vccd1 vccd1 _07259_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10270_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10270_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13960_ _13960_/A _06397_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[25] sky130_fd_sc_hd__ebufn_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07842__A _08084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ _12914_/CLK _12911_/D vssd1 vssd1 vccd1 vccd1 _14038_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_101_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13891_ _13891_/A _06583_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[20] sky130_fd_sc_hd__ebufn_8
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _12842_/CLK _12842_/D vssd1 vssd1 vccd1 vccd1 _12842_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06458__A _11412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12780_/CLK _12773_/D vssd1 vssd1 vccd1 vccd1 _12773_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11724_/A vssd1 vssd1 vccd1 vccd1 _12857_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _11655_/A _11661_/C vssd1 vssd1 vccd1 vccd1 _12840_/D sky130_fd_sc_hd__nor2_1
XFILLER_128_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10606_ _10952_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _10607_/A sky130_fd_sc_hd__and2_1
X_11586_ _11631_/D _11595_/A _11540_/X vssd1 vssd1 vccd1 vccd1 _11587_/B sky130_fd_sc_hd__o21ai_1
XFILLER_155_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10537_ _09773_/X _10525_/X _10535_/X _10536_/X vssd1 vssd1 vccd1 vccd1 _12560_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09708__S _09711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10468_ _10477_/A _10468_/B vssd1 vssd1 vccd1 vccd1 _10469_/A sky130_fd_sc_hd__and2_1
XFILLER_124_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12207_ _11184_/X _12195_/X _12206_/X _12200_/X vssd1 vssd1 vccd1 vccd1 _12980_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08999__S0 _08911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10399_ _10394_/X _10395_/X _10397_/X _10398_/X vssd1 vssd1 vccd1 vccd1 _12523_/D
+ sky130_fd_sc_hd__o211a_1
X_12138_ _12154_/S vssd1 vssd1 vccd1 vccd1 _12151_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11258__B _13948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13754__A _13754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12069_ _10645_/A _12061_/X _12068_/X _11497_/X vssd1 vssd1 vccd1 vccd1 _12939_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_1_clk _12917_/CLK vssd1 vssd1 vccd1 vccd1 _12912_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06630_ _06646_/A _06630_/B _06630_/C vssd1 vssd1 vccd1 vccd1 _06631_/A sky130_fd_sc_hd__or3_1
XFILLER_53_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06561_ _06569_/A _06561_/B _06561_/C vssd1 vssd1 vccd1 vccd1 _06562_/A sky130_fd_sc_hd__or3_1
X_08300_ _08300_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08301_/A sky130_fd_sc_hd__or2_1
X_09280_ _12248_/Q vssd1 vssd1 vccd1 vccd1 _09322_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06492_ _06494_/A _06499_/B _06499_/C vssd1 vssd1 vccd1 vccd1 _06493_/A sky130_fd_sc_hd__or3_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08231_ _08238_/A _08235_/B _08238_/C vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__or3_1
X_13251__407 vssd1 vssd1 vccd1 vccd1 _13251__407/HI _13922_/A sky130_fd_sc_hd__conb_1
XFILLER_165_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08162_ _08174_/A _08174_/B _08164_/C vssd1 vssd1 vccd1 vccd1 _08163_/A sky130_fd_sc_hd__or3_1
XFILLER_146_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07113_ _07121_/A _07118_/B _07115_/C vssd1 vssd1 vccd1 vccd1 _07114_/A sky130_fd_sc_hd__or3_1
XFILLER_119_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08093_ _09125_/B vssd1 vssd1 vccd1 vccd1 _08153_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_161_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07044_ _07044_/A vssd1 vssd1 vccd1 vccd1 _07044_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13145__301 vssd1 vssd1 vccd1 vccd1 _13145__301/HI _13702_/A sky130_fd_sc_hd__conb_1
XFILLER_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08995_ _13971_/A vssd1 vssd1 vccd1 vccd1 _09057_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09861__B _13566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07946_ _07946_/A vssd1 vssd1 vccd1 vccd1 _07946_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07877_ _07881_/A _07877_/B _07877_/C vssd1 vssd1 vccd1 vccd1 _07878_/A sky130_fd_sc_hd__or3_1
XANTENNA__11184__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09616_ _11153_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09616_/X sky130_fd_sc_hd__or2_1
XFILLER_141_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06828_ _06836_/A _06830_/B _07234_/C vssd1 vssd1 vccd1 vccd1 _06829_/A sky130_fd_sc_hd__or3_1
XANTENNA__06278__A _11457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09547_ _09547_/A vssd1 vssd1 vccd1 vccd1 _12312_/D sky130_fd_sc_hd__clkbuf_1
X_06759_ _06759_/A vssd1 vssd1 vccd1 vccd1 _06759_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08914__S0 _08911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ _09478_/A _09478_/B _09478_/C _09478_/D vssd1 vssd1 vccd1 vccd1 _09479_/C
+ sky130_fd_sc_hd__and4_1
X_08429_ _12257_/Q vssd1 vssd1 vccd1 vccd1 _09328_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11440_ _13913_/A _11450_/B vssd1 vssd1 vccd1 vccd1 _11440_/X sky130_fd_sc_hd__or2_1
XFILLER_149_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13839__A _13839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _11377_/A _11371_/B vssd1 vssd1 vccd1 vccd1 _11372_/A sky130_fd_sc_hd__and2_1
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10322_ _10332_/A _10322_/B vssd1 vssd1 vccd1 vccd1 _10323_/A sky130_fd_sc_hd__and2_1
XFILLER_125_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14090_ _14090_/A _08147_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
XFILLER_106_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11359__A _11381_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10253_ _13615_/A _10262_/B vssd1 vssd1 vccd1 vccd1 _10253_/X sky130_fd_sc_hd__or2_1
XFILLER_152_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06460__B _07822_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10184_ _13619_/A _12472_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _10185_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08770__A2 _08765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13943_ _13943_/A _06438_/X vssd1 vssd1 vccd1 vccd1 _14007_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_19_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09180__C1 _09939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13874_ _13874_/A _06629_/X vssd1 vssd1 vccd1 vccd1 _14066_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12067__C1 _11497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ _12829_/CLK _12825_/D vssd1 vssd1 vccd1 vccd1 _12825_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08905__S0 _10697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12758_/CLK _12756_/D vssd1 vssd1 vccd1 vccd1 _13883_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11707_/A _11707_/B _11707_/C _11707_/D vssd1 vssd1 vccd1 vccd1 _11709_/C
+ sky130_fd_sc_hd__or4_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _12687_/CLK _12687_/D vssd1 vssd1 vccd1 vccd1 _13816_/A sky130_fd_sc_hd__dfxtp_1
X_11638_ _12837_/Q vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_11_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10157__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09786__A1 _09112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13749__A _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11569_ _11582_/C vssd1 vssd1 vccd1 vccd1 _11569_/X sky130_fd_sc_hd__buf_2
XFILLER_116_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10173__A _10173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07800_ _07800_/A vssd1 vssd1 vccd1 vccd1 _07800_/X sky130_fd_sc_hd__clkbuf_1
X_08780_ _08887_/A vssd1 vssd1 vccd1 vccd1 _08780_/X sky130_fd_sc_hd__buf_2
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07731_ _07731_/A vssd1 vssd1 vccd1 vccd1 _07731_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__07482__A _08089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10620__B _13746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08513__A2 _08452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07662_ _07672_/A _07669_/B _07664_/C vssd1 vssd1 vccd1 vccd1 _07663_/A sky130_fd_sc_hd__or3_1
XFILLER_65_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09401_ _13596_/A _09791_/B vssd1 vssd1 vccd1 vccd1 _09454_/S sky130_fd_sc_hd__and2_4
XFILLER_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06613_ _06675_/A vssd1 vssd1 vccd1 vccd1 _06625_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__12058__C1 _09404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07593_ _07601_/A _07598_/B _07593_/C vssd1 vssd1 vccd1 vccd1 _07594_/A sky130_fd_sc_hd__or3_1
XFILLER_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09332_ _09336_/A _09332_/B _09334_/D vssd1 vssd1 vccd1 vccd1 _09332_/Y sky130_fd_sc_hd__nand3_1
X_06544_ _07507_/A vssd1 vssd1 vccd1 vccd1 _08180_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09263_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09263_/X sky130_fd_sc_hd__buf_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06475_ _06528_/A vssd1 vssd1 vccd1 vccd1 _06486_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_139_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08214_ _08240_/A vssd1 vssd1 vccd1 vccd1 _08225_/A sky130_fd_sc_hd__clkbuf_1
X_09194_ _11706_/B _11706_/C _11706_/D _11705_/A _13397_/A _13398_/A vssd1 vssd1 vccd1
+ vccd1 _09194_/X sky130_fd_sc_hd__mux4_1
XFILLER_147_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08145_ _08145_/A vssd1 vssd1 vccd1 vccd1 _08145_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09856__B _13554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08076_ _08076_/A vssd1 vssd1 vccd1 vccd1 _08076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07027_ _07031_/A _07031_/B vssd1 vssd1 vccd1 vccd1 _07028_/A sky130_fd_sc_hd__or2_1
XFILLER_161_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09591__B _13564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08978_ _11641_/B _12834_/Q _12835_/Q _11639_/A _08915_/X _08916_/X vssd1 vssd1 vccd1
+ vccd1 _08978_/X sky130_fd_sc_hd__mux4_2
XFILLER_88_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07929_ _07936_/A _07931_/B _07931_/C vssd1 vssd1 vccd1 vccd1 _07930_/A sky130_fd_sc_hd__or3_1
XFILLER_28_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10940_ _10940_/A _11384_/B _10940_/C _10940_/D vssd1 vssd1 vccd1 vccd1 _10942_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10871_ _10871_/A _10871_/B _10871_/C _10871_/D vssd1 vssd1 vccd1 vccd1 _10881_/C
+ sky130_fd_sc_hd__and4_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _12802_/CLK _12610_/D vssd1 vssd1 vccd1 vccd1 _13785_/A sky130_fd_sc_hd__dfxtp_2
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13590_/A _07392_/X vssd1 vssd1 vccd1 vccd1 _14102_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_40_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09112__A _11064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12541_ _12550_/CLK _12541_/D vssd1 vssd1 vccd1 vccd1 _12541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12217__CLK _12217_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ _12659_/CLK _12472_/D vssd1 vssd1 vccd1 vccd1 _12472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13314__470 vssd1 vssd1 vccd1 vccd1 _13314__470/HI _14051_/A sky130_fd_sc_hd__conb_1
XFILLER_138_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13569__A _13569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11423_ _13907_/A _11423_/B vssd1 vssd1 vccd1 vccd1 _11423_/X sky130_fd_sc_hd__or2_1
XFILLER_125_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11354_ _11361_/A _11354_/B vssd1 vssd1 vccd1 vccd1 _11355_/A sky130_fd_sc_hd__and2_1
XFILLER_4_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10305_ _10315_/A _10305_/B vssd1 vssd1 vccd1 vccd1 _10306_/A sky130_fd_sc_hd__and2_1
X_14073_ _14073_/A _08021_/X vssd1 vssd1 vccd1 vccd1 _14105_/Z sky130_fd_sc_hd__ebufn_8
X_11285_ _11412_/A _11285_/B _11412_/C vssd1 vssd1 vccd1 vccd1 _11325_/B sky130_fd_sc_hd__nor3_4
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10236_ _12475_/Q _13750_/A vssd1 vssd1 vccd1 vccd1 _10237_/D sky130_fd_sc_hd__xor2_1
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater100_A _14086_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ _13788_/A _10555_/B vssd1 vssd1 vccd1 vccd1 _10220_/S sky130_fd_sc_hd__and2_2
XFILLER_120_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10098_ _10098_/A _10098_/B _10098_/C vssd1 vssd1 vccd1 vccd1 _10100_/C sky130_fd_sc_hd__and3_1
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10838__B1 _10803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13926_ _13926_/A _06485_/X vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_74_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857_ _13857_/A _06677_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[18] sky130_fd_sc_hd__ebufn_8
XFILLER_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ _12811_/CLK _12808_/D vssd1 vssd1 vccd1 vccd1 _12808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13788_ _13788_/A _06869_/X vssd1 vssd1 vccd1 vccd1 _14108_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11271__B _13947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _12758_/CLK _12739_/D vssd1 vssd1 vccd1 vccd1 _12739_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10168__A _10220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10615__B _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09950_ _13623_/Z _13591_/A _09953_/S vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08901_ _08795_/X _08846_/X _08872_/X _08900_/X _08831_/X _08876_/X vssd1 vssd1 vccd1
+ vccd1 _08901_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _09139_/X _09874_/X _09880_/X _09878_/X vssd1 vssd1 vccd1 vccd1 _12392_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _08741_/X _08747_/X _08744_/X _08752_/X _08876_/A _08831_/X vssd1 vssd1 vccd1
+ vccd1 _08832_/X sky130_fd_sc_hd__mux4_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _12615_/Q _12616_/Q _12617_/Q _12618_/Q _08745_/X _08746_/X vssd1 vssd1 vccd1
+ vccd1 _08763_/X sky130_fd_sc_hd__mux4_2
XANTENNA__13942__A _13942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07714_ _07714_/A _07724_/B _07719_/C vssd1 vssd1 vccd1 vccd1 _07715_/A sky130_fd_sc_hd__or3_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08694_ _13586_/A vssd1 vssd1 vccd1 vccd1 _08694_/X sky130_fd_sc_hd__buf_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257__413 vssd1 vssd1 vccd1 vccd1 _13257__413/HI _13928_/A sky130_fd_sc_hd__conb_1
X_07645_ _07645_/A vssd1 vssd1 vccd1 vccd1 _07645_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07576_ _07576_/A vssd1 vssd1 vccd1 vccd1 _07576_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09315_ _09315_/A _09315_/B _09315_/C _09315_/D vssd1 vssd1 vccd1 vccd1 _09318_/B
+ sky130_fd_sc_hd__and4_1
X_06527_ _06527_/A vssd1 vssd1 vccd1 vccd1 _06527_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09246_ _09246_/A vssd1 vssd1 vccd1 vccd1 _12239_/D sky130_fd_sc_hd__clkbuf_1
X_06458_ _11412_/B vssd1 vssd1 vccd1 vccd1 _08276_/B sky130_fd_sc_hd__buf_2
XFILLER_139_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09586__B _13560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ _14072_/Z vssd1 vssd1 vccd1 vccd1 _09638_/A sky130_fd_sc_hd__buf_4
X_06389_ _08338_/A vssd1 vssd1 vccd1 vccd1 _07845_/B sky130_fd_sc_hd__buf_2
XFILLER_5_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08128_ _08135_/A _08128_/B _08138_/C vssd1 vssd1 vccd1 vccd1 _08129_/A sky130_fd_sc_hd__or3_1
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07818__C _08110_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08059_ _08072_/A vssd1 vssd1 vccd1 vccd1 _08070_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_162_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11309__A1 _10665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput35 _13402_/A vssd1 vssd1 vccd1 vccd1 pwm_en[1] sky130_fd_sc_hd__buf_2
XFILLER_122_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput46 _13762_/A vssd1 vssd1 vccd1 vccd1 pwm_out[11] sky130_fd_sc_hd__buf_2
XFILLER_89_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput57 _13570_/A vssd1 vssd1 vccd1 vccd1 pwm_out[7] sky130_fd_sc_hd__buf_2
X_11070_ _13822_/A _11070_/B vssd1 vssd1 vccd1 vccd1 _11070_/X sky130_fd_sc_hd__or2_1
XFILLER_163_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10021_ _10024_/B _10021_/B _10021_/C _10021_/D vssd1 vssd1 vccd1 vccd1 _10030_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_103_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09107__A _09967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11972_ _11978_/A _11972_/B vssd1 vssd1 vccd1 vccd1 _11973_/A sky130_fd_sc_hd__and2_1
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13711_ _13711_/A _07980_/X vssd1 vssd1 vccd1 vccd1 _14063_/Z sky130_fd_sc_hd__ebufn_8
X_10923_ _10921_/B _10915_/X _10921_/A vssd1 vssd1 vccd1 vccd1 _10923_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13642_ _13642_/A _07247_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
X_10854_ _10876_/A _10868_/D _10854_/C vssd1 vssd1 vccd1 vccd1 _10859_/B sky130_fd_sc_hd__and3_1
XFILLER_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06466__A _06729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13573_ _13573_/A _07436_/X vssd1 vssd1 vccd1 vccd1 _13765_/Z sky130_fd_sc_hd__ebufn_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _10865_/B _10865_/C _10865_/D _10785_/D vssd1 vssd1 vccd1 vccd1 _10794_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_157_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09777__A _09789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ _12533_/CLK _12524_/D vssd1 vssd1 vccd1 vccd1 _13653_/A sky130_fd_sc_hd__dfxtp_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12455_ _12461_/CLK _12455_/D vssd1 vssd1 vccd1 vccd1 _12455_/Q sky130_fd_sc_hd__dfxtp_1
X_13050__206 vssd1 vssd1 vccd1 vccd1 _13050__206/HI _13509_/A sky130_fd_sc_hd__conb_1
X_11406_ _11406_/A _11406_/B _11406_/C vssd1 vssd1 vccd1 vccd1 _11406_/Y sky130_fd_sc_hd__nor3_1
XFILLER_165_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12386_ _12386_/CLK _12386_/D vssd1 vssd1 vccd1 vccd1 _12386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ _14125_/A _08275_/X vssd1 vssd1 vccd1 vccd1 _14125_/Z sky130_fd_sc_hd__ebufn_8
X_11337_ _11344_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11338_/A sky130_fd_sc_hd__and2_1
XFILLER_98_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14056_ _14056_/A _07930_/X vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__ebufn_8
X_11268_ _11268_/A _11268_/B _11268_/C _11268_/D vssd1 vssd1 vccd1 vccd1 _11279_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_95_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10219_ _10219_/A vssd1 vssd1 vccd1 vccd1 _12482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11199_ _13854_/A _11199_/B vssd1 vssd1 vccd1 vccd1 _11199_/X sky130_fd_sc_hd__or2_1
XANTENNA__11266__B _13941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13762__A _13762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09451__S _09454_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10287__A1 _10285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ _13909_/A _06531_/X vssd1 vssd1 vccd1 vccd1 _14069_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07430_ _07430_/A _07435_/B vssd1 vssd1 vccd1 vccd1 _07431_/A sky130_fd_sc_hd__or2_1
XFILLER_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06376__A input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10039__A1 _09982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07361_ _07369_/A _07364_/B _07361_/C vssd1 vssd1 vccd1 vccd1 _07362_/A sky130_fd_sc_hd__or3_1
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09100_ _12195_/A vssd1 vssd1 vccd1 vccd1 _09100_/X sky130_fd_sc_hd__clkbuf_2
X_06312_ _06462_/A vssd1 vssd1 vccd1 vccd1 _06323_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_31_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07292_ _07292_/A _07303_/B _07300_/C vssd1 vssd1 vccd1 vccd1 _07293_/A sky130_fd_sc_hd__or3_1
XFILLER_148_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09031_ _08987_/X _08993_/X _08991_/X _08999_/X _09024_/X _09030_/X vssd1 vssd1 vccd1
+ vccd1 _09031_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13937__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09933_ _09933_/A vssd1 vssd1 vccd1 vccd1 _12409_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07935__A _08004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11457__A _11457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _12374_/Q _13551_/A vssd1 vssd1 vccd1 vccd1 _09868_/A sky130_fd_sc_hd__xor2_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _10869_/C _12634_/Q _10870_/A _10876_/D _08733_/X _08735_/X vssd1 vssd1 vccd1
+ vccd1 _08815_/X sky130_fd_sc_hd__mux4_2
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _09795_/A vssd1 vssd1 vccd1 vccd1 _12374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08746_ _13777_/A vssd1 vssd1 vccd1 vccd1 _08746_/X sky130_fd_sc_hd__buf_2
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08766__A _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11475__A0 _14099_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11904__B _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08566__S1 _08560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _09396_/D vssd1 vssd1 vccd1 vccd1 _13558_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_53_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _08035_/A vssd1 vssd1 vccd1 vccd1 _08022_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07559_ _07559_/A vssd1 vssd1 vccd1 vccd1 _07559_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ _10971_/A vssd1 vssd1 vccd1 vccd1 _10585_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09229_ _09316_/C _09226_/A _09217_/X vssd1 vssd1 vccd1 vccd1 _09230_/B sky130_fd_sc_hd__o21ai_1
XFILLER_139_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10536__A _10650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ _12242_/CLK _12240_/D vssd1 vssd1 vccd1 vccd1 _12240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12171_ _12171_/A _12171_/B _12171_/C _12171_/D vssd1 vssd1 vccd1 vccd1 _12177_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_135_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11122_ _11204_/A _11122_/B vssd1 vssd1 vccd1 vccd1 _11123_/A sky130_fd_sc_hd__and2_1
XFILLER_1_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11053_ _11195_/A vssd1 vssd1 vccd1 vccd1 _11053_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10004_ _10004_/A _10004_/B vssd1 vssd1 vccd1 vccd1 _12429_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09659__A0 _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11955_ _11962_/A _11955_/B vssd1 vssd1 vccd1 vccd1 _11956_/A sky130_fd_sc_hd__and2_1
XFILLER_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12555__CLK _12555_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10906_ _10907_/A vssd1 vssd1 vccd1 vccd1 _10906_/Y sky130_fd_sc_hd__inv_2
X_11886_ _11886_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _11887_/A sky130_fd_sc_hd__and2_1
XFILLER_72_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13625_ _13625_/A _07293_/X vssd1 vssd1 vccd1 vccd1 _13625_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_60_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10837_ _10876_/D vssd1 vssd1 vccd1 vccd1 _10869_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater65 peripheralBus_data[8] vssd1 vssd1 vccd1 vccd1 _14007_/Z sky130_fd_sc_hd__buf_12
X_13556_ _13556_/A _07477_/X vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_13_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater76 _14035_/Z vssd1 vssd1 vccd1 vccd1 _14067_/Z sky130_fd_sc_hd__buf_12
X_10768_ _10768_/A vssd1 vssd1 vccd1 vccd1 _10936_/A sky130_fd_sc_hd__clkbuf_4
Xrepeater87 peripheralBus_data[2] vssd1 vssd1 vccd1 vccd1 _14033_/Z sky130_fd_sc_hd__buf_12
Xrepeater98 _14119_/Z vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__buf_12
XFILLER_157_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12507_ _12515_/CLK _12507_/D vssd1 vssd1 vccd1 vccd1 _12507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07739__B _07947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13487_ _13487_/A _08111_/X vssd1 vssd1 vccd1 vccd1 _13775_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10446__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12179__D1 _13401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10699_ _14097_/Z _08887_/X _10703_/S vssd1 vssd1 vccd1 vccd1 _10700_/B sky130_fd_sc_hd__mux2_1
XFILLER_157_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12438_ _12438_/CLK _12438_/D vssd1 vssd1 vccd1 vccd1 _12438_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12194__A1 _11170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13757__A _13757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12369_ _12369_/CLK _12369_/D vssd1 vssd1 vccd1 vccd1 _13498_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14108_ _14108_/A _08232_/X vssd1 vssd1 vccd1 vccd1 _14108_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_113_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14039_ _14039_/A _07885_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[8] sky130_fd_sc_hd__ebufn_8
X_06930_ _06930_/A vssd1 vssd1 vccd1 vccd1 _06930_/X sky130_fd_sc_hd__clkbuf_1
X_06861_ _06863_/A _06870_/B _06870_/C vssd1 vssd1 vccd1 vccd1 _06862_/A sky130_fd_sc_hd__or3_1
XFILLER_95_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08600_ _09851_/B vssd1 vssd1 vccd1 vccd1 _13552_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__13492__A _13492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06792_ _06792_/A vssd1 vssd1 vccd1 vccd1 _06792_/X sky130_fd_sc_hd__clkbuf_1
X_09580_ _09580_/A vssd1 vssd1 vccd1 vccd1 _12322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08531_ _12269_/Q vssd1 vssd1 vccd1 vccd1 _09377_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08462_ _08452_/X _08455_/X _08458_/X _08461_/X _08448_/X _08449_/X vssd1 vssd1 vccd1
+ vccd1 _08462_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07413_ _08168_/A _07423_/B vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__or2_1
XANTENNA__10680__A1 _10285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08393_ _08384_/X _08391_/X _08498_/S vssd1 vssd1 vccd1 vccd1 _11706_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07344_ _07371_/A vssd1 vssd1 vccd1 vccd1 _07356_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07275_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07286_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_164_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09014_ _08917_/X _08923_/X _08920_/X _08930_/X _09057_/A _09013_/X vssd1 vssd1 vccd1
+ vccd1 _09014_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12185__A1 _11160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09864__B _13551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09916_ _10256_/A vssd1 vssd1 vccd1 vccd1 _09916_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_6_0_clk_A clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ _12383_/Q _13560_/A vssd1 vssd1 vccd1 vccd1 _09847_/Y sky130_fd_sc_hd__xnor2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09778_ _13497_/A _09787_/B vssd1 vssd1 vccd1 vccd1 _09778_/X sky130_fd_sc_hd__or2_1
XFILLER_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _09399_/D vssd1 vssd1 vccd1 vccd1 _13566_/A sky130_fd_sc_hd__buf_6
XFILLER_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11740_ _11740_/A _11740_/B vssd1 vssd1 vccd1 vccd1 _11741_/A sky130_fd_sc_hd__and2_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11676_/A _11676_/B _11677_/A _11677_/B vssd1 vssd1 vccd1 vccd1 _11672_/C
+ sky130_fd_sc_hd__and4_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13410_ _13410_/A _08102_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10622_ _10622_/A _10622_/B _10622_/C _10622_/D vssd1 vssd1 vccd1 vccd1 _10633_/A
+ sky130_fd_sc_hd__or4_1
XANTENNA__09120__A _10552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10553_ _13694_/A _10553_/B vssd1 vssd1 vccd1 vccd1 _10553_/X sky130_fd_sc_hd__or2_1
XFILLER_10_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10484_ _12545_/Q _13754_/A vssd1 vssd1 vccd1 vccd1 _10484_/Y sky130_fd_sc_hd__nor2_1
XFILLER_154_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12223_ _12325_/CLK _12223_/D vssd1 vssd1 vccd1 vccd1 _13400_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11923__A1 _13377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12154_ _12968_/Q _14110_/A _12154_/S vssd1 vssd1 vccd1 vccd1 _12155_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11097__A _11206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _13848_/A _12703_/Q _11118_/S vssd1 vssd1 vccd1 vccd1 _11106_/B sky130_fd_sc_hd__mux2_1
X_13162__318 vssd1 vssd1 vccd1 vccd1 _13162__318/HI _13735_/A sky130_fd_sc_hd__conb_1
X_12085_ _10665_/A _12075_/X _12083_/X _12084_/X vssd1 vssd1 vccd1 vccd1 _12945_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11036_ _13810_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11036_/X sky130_fd_sc_hd__or2_1
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13203__359 vssd1 vssd1 vccd1 vccd1 _13203__359/HI _13826_/A sky130_fd_sc_hd__conb_1
XFILLER_80_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12100__A1 _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11938_ _11945_/A _11938_/B vssd1 vssd1 vccd1 vccd1 _11939_/A sky130_fd_sc_hd__and2_1
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13056__212 vssd1 vssd1 vccd1 vccd1 _13056__212/HI _13515_/A sky130_fd_sc_hd__conb_1
X_11869_ _11869_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _11870_/A sky130_fd_sc_hd__and2_1
X_13608_ _13608_/A _07343_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_158_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06654__A _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11611__B1 _11569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13539_ _13539_/A _07518_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07060_ _08364_/B _07995_/B _07969_/B vssd1 vssd1 vccd1 vccd1 _07061_/A sky130_fd_sc_hd__or3_1
XFILLER_118_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13487__A _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10904__A _10936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10623__B _13758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07962_ _07962_/A _07962_/B _07962_/C vssd1 vssd1 vccd1 vccd1 _07963_/A sky130_fd_sc_hd__or3_1
X_09701_ _13499_/A _12353_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09702_/B sky130_fd_sc_hd__mux2_1
X_06913_ _06913_/A vssd1 vssd1 vccd1 vccd1 _06923_/A sky130_fd_sc_hd__clkbuf_1
X_07893_ _07920_/A vssd1 vssd1 vccd1 vccd1 _07903_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_56_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ _13461_/A _09627_/X _09631_/X _09621_/X vssd1 vssd1 vccd1 vccd1 _12331_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06844_ _06844_/A vssd1 vssd1 vccd1 vccd1 _06844_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09563_ _09563_/A _09563_/B vssd1 vssd1 vccd1 vccd1 _09564_/A sky130_fd_sc_hd__and2_1
X_06775_ _06775_/A _06780_/B _06780_/C vssd1 vssd1 vccd1 vccd1 _06776_/A sky130_fd_sc_hd__or3_1
XFILLER_71_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13950__A _13950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ _12268_/Q vssd1 vssd1 vccd1 vccd1 _09377_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09494_ _11929_/A vssd1 vssd1 vccd1 vccd1 _12134_/A sky130_fd_sc_hd__clkbuf_2
X_08445_ _08524_/A vssd1 vssd1 vccd1 vccd1 _08445_/X sky130_fd_sc_hd__buf_2
XANTENNA__09859__B _13553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08376_ _13392_/A vssd1 vssd1 vccd1 vccd1 _08376_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10405__A1 _09770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07327_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07739_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_109_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09875__A _11412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07258_ _07266_/A _07263_/B _07260_/C vssd1 vssd1 vccd1 vccd1 _07259_/A sky130_fd_sc_hd__or3_1
XFILLER_3_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09594__B _13557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07189_ _07230_/A vssd1 vssd1 vccd1 vccd1 _07200_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_100_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_115_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12910_ _12914_/CLK _12910_/D vssd1 vssd1 vccd1 vccd1 _14037_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13890_ _13890_/A _06585_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09115__A peripheralBus_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ _12842_/CLK _12841_/D vssd1 vssd1 vccd1 vccd1 _12841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12775_/CLK _12772_/D vssd1 vssd1 vccd1 vccd1 _12772_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11723_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11724_/A sky130_fd_sc_hd__and2_1
XANTENNA__10644__A1 _10385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11680_/A _11657_/B _11657_/C _11672_/A vssd1 vssd1 vccd1 vccd1 _11661_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__06474__A _06694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10605_ _13725_/A _12581_/Q _10608_/S vssd1 vssd1 vccd1 vccd1 _10606_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ _11631_/D _11595_/A vssd1 vssd1 vccd1 vccd1 _11587_/A sky130_fd_sc_hd__and2_1
XFILLER_155_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10536_ _10650_/A vssd1 vssd1 vccd1 vccd1 _10536_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater130_A peripheralBus_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _13690_/A _12545_/Q _10473_/S vssd1 vssd1 vccd1 vccd1 _10468_/B sky130_fd_sc_hd__mux2_1
X_12206_ _14105_/A _12206_/B vssd1 vssd1 vccd1 vccd1 _12206_/X sky130_fd_sc_hd__or2_1
XFILLER_89_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08999__S1 _08913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10398_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10398_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ _12137_/A vssd1 vssd1 vccd1 vccd1 _12962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12068_ _14065_/A _12073_/B vssd1 vssd1 vccd1 vccd1 _12068_/X sky130_fd_sc_hd__or2_1
XFILLER_38_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11019_ _12669_/Q _13943_/A vssd1 vssd1 vccd1 vccd1 _11021_/C sky130_fd_sc_hd__xor2_1
XFILLER_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11274__B _13940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06560_ _06560_/A vssd1 vssd1 vccd1 vccd1 _06560_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06491_ _06491_/A vssd1 vssd1 vccd1 vccd1 _06491_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13290__446 vssd1 vssd1 vccd1 vccd1 _13290__446/HI _13995_/A sky130_fd_sc_hd__conb_1
X_08230_ _08230_/A vssd1 vssd1 vccd1 vccd1 _08230_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10618__B _13753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08161_ _08161_/A vssd1 vssd1 vccd1 vccd1 _08161_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11060__A1 _10414_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07112_ _07112_/A vssd1 vssd1 vccd1 vccd1 _07112_/X sky130_fd_sc_hd__clkbuf_1
X_13331__487 vssd1 vssd1 vccd1 vccd1 _13331__487/HI _14084_/A sky130_fd_sc_hd__conb_1
X_08092_ _08150_/A vssd1 vssd1 vccd1 vccd1 _08110_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_118_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07043_ _07043_/A _07043_/B vssd1 vssd1 vccd1 vccd1 _07044_/A sky130_fd_sc_hd__or2_1
XANTENNA__08439__S0 _08417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10353__B _10613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13184__340 vssd1 vssd1 vccd1 vccd1 _13184__340/HI _13791_/A sky130_fd_sc_hd__conb_1
XANTENNA__13945__A _13945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08994_ _13970_/A vssd1 vssd1 vccd1 vccd1 _08994_/X sky130_fd_sc_hd__buf_2
XFILLER_88_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07945_ _07951_/A _07945_/B _07945_/C vssd1 vssd1 vccd1 vccd1 _07946_/A sky130_fd_sc_hd__or3_1
X_13225__381 vssd1 vssd1 vccd1 vccd1 _13225__381/HI _13864_/A sky130_fd_sc_hd__conb_1
X_07876_ _07876_/A vssd1 vssd1 vccd1 vccd1 _07876_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09615_ _09655_/B vssd1 vssd1 vccd1 vccd1 _09625_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06827_ _06827_/A vssd1 vssd1 vccd1 vccd1 _06827_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ _09546_/A _09546_/B vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__and2_1
XFILLER_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06758_ _06760_/A _06765_/B _06765_/C vssd1 vssd1 vccd1 vccd1 _06759_/A sky130_fd_sc_hd__or3_1
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11823__A0 _09638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__B _13374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09589__B _13552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ _12282_/Q _13558_/A vssd1 vssd1 vccd1 vccd1 _09478_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__08914__S1 _08913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06689_ _06748_/A vssd1 vssd1 vccd1 vccd1 _06701_/A sky130_fd_sc_hd__clkbuf_1
X_08428_ _09321_/B _12251_/Q _12252_/Q _12253_/Q _08404_/X _08405_/X vssd1 vssd1 vccd1
+ vccd1 _08428_/X sky130_fd_sc_hd__mux4_2
XANTENNA__06294__A _08186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08359_ _08359_/A vssd1 vssd1 vccd1 vccd1 _08359_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ _13915_/A _12772_/Q _11373_/S vssd1 vssd1 vccd1 vccd1 _11371_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10321_ _13654_/A _12508_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10322_/B sky130_fd_sc_hd__mux2_1
XFILLER_3_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07837__B _07840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10252_ _10293_/B vssd1 vssd1 vccd1 vccd1 _10262_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_117_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10183_ _10220_/S vssd1 vssd1 vccd1 vccd1 _10197_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_105_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_3_0_clk_A clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13942_ _13942_/A _06441_/X vssd1 vssd1 vccd1 vccd1 _14070_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__07572__B _07995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13873_ _13873_/A _06631_/X vssd1 vssd1 vccd1 vccd1 _14065_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12824_ _12829_/CLK _12824_/D vssd1 vssd1 vccd1 vccd1 _12824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12755_ _12758_/CLK _12755_/D vssd1 vssd1 vccd1 vccd1 _13882_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__A1 _11160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11706_ _11706_/A _11706_/B _11706_/C _11706_/D vssd1 vssd1 vccd1 vccd1 _11709_/B
+ sky130_fd_sc_hd__or4_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12806_/CLK _12686_/D vssd1 vssd1 vccd1 vccd1 _13815_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11637_ _11637_/A vssd1 vssd1 vccd1 vccd1 _12836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11568_ _11568_/A vssd1 vssd1 vccd1 vccd1 _12821_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10519_ _09750_/X _10511_/X _10518_/X _10425_/X vssd1 vssd1 vccd1 vccd1 _12553_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11499_ _14012_/Z _11499_/B vssd1 vssd1 vccd1 vccd1 _11499_/X sky130_fd_sc_hd__or2_1
X_13168__324 vssd1 vssd1 vccd1 vccd1 _13168__324/HI _13741_/A sky130_fd_sc_hd__conb_1
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11269__B _13942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09454__S _09454_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209__365 vssd1 vssd1 vccd1 vccd1 _13209__365/HI _13832_/A sky130_fd_sc_hd__conb_1
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07730_ _07742_/A _07737_/B _07732_/C vssd1 vssd1 vccd1 vccd1 _07731_/A sky130_fd_sc_hd__or3_1
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06379__A _07480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08513__A3 _08455_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ _07661_/A vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09400_ _09400_/A _09400_/B _09400_/C _09400_/D vssd1 vssd1 vccd1 vccd1 _09791_/B
+ sky130_fd_sc_hd__or4_1
X_06612_ _06688_/A vssd1 vssd1 vccd1 vccd1 _06675_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07592_ _07592_/A vssd1 vssd1 vccd1 vccd1 _07592_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09331_ _09331_/A _09331_/B _09331_/C _09331_/D vssd1 vssd1 vccd1 vccd1 _09334_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__11805__A0 _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06543_ _06604_/A vssd1 vssd1 vccd1 vccd1 _06561_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09262_ _09332_/B vssd1 vssd1 vccd1 vccd1 _09262_/Y sky130_fd_sc_hd__inv_2
X_06474_ _06694_/A vssd1 vssd1 vccd1 vccd1 _06528_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06545__C _08180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08213_ _08213_/A vssd1 vssd1 vccd1 vccd1 _08213_/X sky130_fd_sc_hd__clkbuf_1
X_09193_ _09112_/X _09152_/B _09191_/X _09192_/X vssd1 vssd1 vccd1 vccd1 _12227_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11033__A1 _10385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07938__A _07999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _08148_/A _08151_/B _08151_/C vssd1 vssd1 vccd1 vccd1 _08145_/A sky130_fd_sc_hd__or3_1
XFILLER_146_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08075_ _08075_/A _08075_/B _08110_/C vssd1 vssd1 vccd1 vccd1 _08076_/A sky130_fd_sc_hd__or3_1
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07026_ _07026_/A vssd1 vssd1 vccd1 vccd1 _07026_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11907__B _13365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08977_ _12836_/Q vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11195__A _11195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07928_ _07928_/A vssd1 vssd1 vccd1 vccd1 _07928_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07859_ _07861_/A _07962_/B _07863_/B vssd1 vssd1 vccd1 vccd1 _07860_/A sky130_fd_sc_hd__or3_1
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10870_ _10870_/A _10870_/B _10874_/B _10870_/D vssd1 vssd1 vccd1 vccd1 _10871_/D
+ sky130_fd_sc_hd__and4_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09671_/A vssd1 vssd1 vccd1 vccd1 _09546_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13002__158 vssd1 vssd1 vccd1 vccd1 _13002__158/HI _13413_/A sky130_fd_sc_hd__conb_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _12550_/CLK _12540_/D vssd1 vssd1 vccd1 vccd1 _12540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12471_ _12492_/CLK _12471_/D vssd1 vssd1 vccd1 vccd1 _12471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11422_ _10648_/X _11411_/X _11421_/X _11417_/X vssd1 vssd1 vccd1 vccd1 _12780_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11353_ _13910_/A _12767_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _11354_/B sky130_fd_sc_hd__mux2_1
X_10304_ _13649_/A _12503_/Q _10375_/B vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__mux2_1
X_14072_ _14072_/A _08017_/X vssd1 vssd1 vccd1 vccd1 _14072_/Z sky130_fd_sc_hd__ebufn_8
X_11284_ _11312_/A vssd1 vssd1 vccd1 vccd1 _11284_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10235_ _12470_/Q _13745_/A vssd1 vssd1 vccd1 vccd1 _10237_/C sky130_fd_sc_hd__xor2_1
XFILLER_106_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10166_ _10166_/A _10166_/B _10166_/C _10166_/D vssd1 vssd1 vccd1 vccd1 _10555_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10097_ _10097_/A _10097_/B _10097_/C vssd1 vssd1 vccd1 vccd1 _10100_/B sky130_fd_sc_hd__and3_1
XFILLER_75_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13925_ _13925_/A _06487_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13856_ _13856_/A _06679_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[17] sky130_fd_sc_hd__ebufn_8
XFILLER_62_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ _12821_/CLK _12807_/D vssd1 vssd1 vccd1 vccd1 _12807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13787_ _13787_/A _06871_/X vssd1 vssd1 vccd1 vccd1 _14075_/Z sky130_fd_sc_hd__ebufn_8
X_10999_ _12670_/Q _13944_/A vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__or2_1
X_12738_ _12753_/CLK _12738_/D vssd1 vssd1 vccd1 vccd1 _12738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12669_ _12853_/CLK _12669_/D vssd1 vssd1 vccd1 vccd1 _12669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08900_ _10921_/A _10928_/B _12658_/Q _12659_/Q _10697_/A _08887_/X vssd1 vssd1 vccd1
+ vccd1 _08900_/X sky130_fd_sc_hd__mux4_2
XANTENNA__13495__A _13495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _13520_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09880_/X sky130_fd_sc_hd__or2_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07493__A _07507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _13778_/A vssd1 vssd1 vccd1 vccd1 _08831_/X sky130_fd_sc_hd__clkbuf_2
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10631__B _13743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08762_ _10163_/A vssd1 vssd1 vccd1 vccd1 _13743_/A sky130_fd_sc_hd__buf_6
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07713_ _07892_/A vssd1 vssd1 vccd1 vccd1 _07724_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_122_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08693_ _09398_/C vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__buf_4
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07644_ _07644_/A _07654_/B _07649_/C vssd1 vssd1 vccd1 vccd1 _07645_/A sky130_fd_sc_hd__or3_1
XFILLER_93_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13296__452 vssd1 vssd1 vccd1 vccd1 _13296__452/HI _14017_/A sky130_fd_sc_hd__conb_1
XFILLER_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09213__A _09281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07575_ _07575_/A _07585_/B _07580_/C vssd1 vssd1 vccd1 vccd1 _07576_/A sky130_fd_sc_hd__or3_1
XFILLER_80_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09314_ _09314_/A vssd1 vssd1 vccd1 vccd1 _12256_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06526_ _06534_/A _06526_/B _06526_/C vssd1 vssd1 vccd1 vccd1 _06527_/A sky130_fd_sc_hd__or3_1
X_13337__493 vssd1 vssd1 vccd1 vccd1 _13337__493/HI _14090_/A sky130_fd_sc_hd__conb_1
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09245_ _09253_/C _09389_/A _09245_/C vssd1 vssd1 vccd1 vccd1 _09246_/A sky130_fd_sc_hd__and3b_1
XANTENNA__09867__B _09867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06457_ _08210_/A vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__buf_4
XFILLER_21_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09176_ _10665_/A _09145_/A _09174_/X _09939_/A vssd1 vssd1 vccd1 vccd1 _12222_/D
+ sky130_fd_sc_hd__a211o_1
X_06388_ _06388_/A vssd1 vssd1 vccd1 vccd1 _06388_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08127_ _08127_/A vssd1 vssd1 vccd1 vccd1 _08127_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10765__B1 _10757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08058_ _08058_/A vssd1 vssd1 vccd1 vccd1 _08058_/X sky130_fd_sc_hd__clkbuf_1
Xoutput36 _13403_/A vssd1 vssd1 vccd1 vccd1 pwm_en[2] sky130_fd_sc_hd__buf_2
X_07009_ _07033_/A vssd1 vssd1 vccd1 vccd1 _07019_/A sky130_fd_sc_hd__clkbuf_1
Xoutput47 _13951_/A vssd1 vssd1 vccd1 vccd1 pwm_out[12] sky130_fd_sc_hd__buf_2
Xoutput58 _13759_/A vssd1 vssd1 vccd1 vccd1 pwm_out[8] sky130_fd_sc_hd__buf_2
XFILLER_163_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08805__S0 _08733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__B1 _09236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _10020_/A vssd1 vssd1 vccd1 vccd1 _12433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11971_ _14108_/Z _14044_/A _11974_/S vssd1 vssd1 vccd1 vccd1 _11972_/B sky130_fd_sc_hd__mux2_1
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13710_ _13710_/A _07061_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11493__A1 _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07850__B _07854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ _10922_/A _10922_/B _10922_/C _10922_/D vssd1 vssd1 vccd1 vccd1 _10928_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_72_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09123__A _13775_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13641_ _13641_/A _07251_/X vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_8
X_10853_ _10868_/D _10854_/C _10852_/Y vssd1 vssd1 vccd1 vccd1 _12640_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__10269__A _10667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _13572_/A _07439_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _12624_/Q vssd1 vssd1 vccd1 vccd1 _10865_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12523_ _12533_/CLK _12523_/D vssd1 vssd1 vccd1 vccd1 _13652_/A sky130_fd_sc_hd__dfxtp_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12454_ _12457_/CLK _12454_/D vssd1 vssd1 vccd1 vccd1 _12454_/Q sky130_fd_sc_hd__dfxtp_1
X_11405_ _11405_/A _11405_/B _11405_/C _11405_/D vssd1 vssd1 vccd1 vccd1 _11406_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_125_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12385_ _12400_/CLK _12385_/D vssd1 vssd1 vccd1 vccd1 _12385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14124_ _14124_/A _08273_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[29] sky130_fd_sc_hd__ebufn_8
XFILLER_126_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11336_ _13905_/A _12762_/Q _11408_/B vssd1 vssd1 vccd1 vccd1 _11337_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13130__286 vssd1 vssd1 vccd1 vccd1 _13130__286/HI _13671_/A sky130_fd_sc_hd__conb_1
XFILLER_153_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14055_ _14055_/A _07928_/X vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11828__A _11834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ _12730_/Q _13938_/A vssd1 vssd1 vccd1 vccd1 _11268_/D sky130_fd_sc_hd__xor2_1
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10732__A _13788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09374__B1 _09392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10218_ _10298_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10219_/A sky130_fd_sc_hd__and2_1
X_11198_ _10548_/X _11185_/X _11197_/X _11195_/X vssd1 vssd1 vccd1 vccd1 _12725_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10149_ _10149_/A _10149_/B _10149_/C vssd1 vssd1 vccd1 vccd1 _10155_/C sky130_fd_sc_hd__and3_1
XFILLER_94_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _13908_/A _06533_/X vssd1 vssd1 vccd1 vccd1 _14068_/Z sky130_fd_sc_hd__ebufn_8
X_13024__180 vssd1 vssd1 vccd1 vccd1 _13024__180/HI _13451_/A sky130_fd_sc_hd__conb_1
XFILLER_90_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13839_ _13839_/A _07860_/X vssd1 vssd1 vccd1 vccd1 _14063_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09968__A _09977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07360_ _07360_/A vssd1 vssd1 vccd1 vccd1 _07360_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06311_ _06688_/A vssd1 vssd1 vccd1 vccd1 _06462_/A sky130_fd_sc_hd__buf_2
X_07291_ _07291_/A vssd1 vssd1 vccd1 vccd1 _07303_/B sky130_fd_sc_hd__clkbuf_1
X_09030_ _09030_/A vssd1 vssd1 vccd1 vccd1 _09030_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10626__B _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09932_ _09939_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__or2_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater92_A _13994_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11457__B _11457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _09863_/A _09863_/B _09863_/C _09863_/D vssd1 vssd1 vccd1 vccd1 _09869_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10361__B _13757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _12633_/Q vssd1 vssd1 vccd1 vccd1 _10869_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13953__A _13953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09800_/A _09794_/B vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__and2_1
XFILLER_39_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater130 peripheralBus_data[11] vssd1 vssd1 vccd1 vccd1 _13978_/Z sky130_fd_sc_hd__buf_12
X_08745_ _13776_/A vssd1 vssd1 vccd1 vccd1 _08745_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_54_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08676_ _08671_/X _08675_/X _08712_/S vssd1 vssd1 vccd1 vccd1 _09396_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07627_/A vssd1 vssd1 vccd1 vccd1 _07627_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07558_ _07558_/A _07558_/B _07564_/C vssd1 vssd1 vccd1 vccd1 _07559_/A sky130_fd_sc_hd__or3_1
XFILLER_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_2_0_clk_A clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073__229 vssd1 vssd1 vccd1 vccd1 _13073__229/HI _13548_/A sky130_fd_sc_hd__conb_1
X_06509_ _06523_/A vssd1 vssd1 vccd1 vccd1 _06521_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_158_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10817__A _13775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07489_ _07489_/A vssd1 vssd1 vccd1 vccd1 _07489_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09228_ _13391_/A _09318_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _09235_/C sky130_fd_sc_hd__and3_1
XANTENNA__07398__A _07964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09159_ _14100_/Z vssd1 vssd1 vccd1 vccd1 _11170_/A sky130_fd_sc_hd__buf_4
X_12170_ _12965_/Q _13371_/A vssd1 vssd1 vccd1 vccd1 _12171_/D sky130_fd_sc_hd__xor2_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11121_ _13853_/A _12708_/Q _11124_/S vssd1 vssd1 vccd1 vccd1 _11122_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07845__B _07845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__A _10552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11052_ _11443_/A vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__buf_2
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08022__A _08022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10003_ _10029_/D _10008_/D _09994_/X vssd1 vssd1 vccd1 vccd1 _10004_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__07861__A _07861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A peripheralBus_address[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008__164 vssd1 vssd1 vccd1 vccd1 _13008__164/HI _13419_/A sky130_fd_sc_hd__conb_1
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13_0_clk_A clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11954_ _09636_/A _14039_/A _11957_/S vssd1 vssd1 vccd1 vccd1 _11955_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06477__A _06481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10905_ _10905_/A vssd1 vssd1 vccd1 vccd1 _12651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11885_ _12898_/Q _14042_/A _11895_/S vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__mux2_1
X_13624_ _13624_/A _07297_/X vssd1 vssd1 vccd1 vccd1 _14072_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10836_ _10836_/A vssd1 vssd1 vccd1 vccd1 _12635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13555_ _13555_/A _07479_/X vssd1 vssd1 vccd1 vccd1 _14035_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ _10864_/C _10864_/D _10767_/C vssd1 vssd1 vccd1 vccd1 _10785_/D sky130_fd_sc_hd__and3_1
Xrepeater66 _14102_/Z vssd1 vssd1 vccd1 vccd1 _13974_/Z sky130_fd_sc_hd__buf_12
Xrepeater77 peripheralBus_data[4] vssd1 vssd1 vccd1 vccd1 _14035_/Z sky130_fd_sc_hd__buf_12
XFILLER_158_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater88 _14028_/Z vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__buf_12
XFILLER_146_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ _12515_/CLK _12506_/D vssd1 vssd1 vccd1 vccd1 _12506_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater99 peripheralBus_data[24] vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__buf_12
X_13486_ _13486_/A _07657_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__07739__C _07739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10698_ _10385_/X _10690_/X _10697_/X _10682_/X vssd1 vssd1 vccd1 vccd1 _12601_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12179__C1 _09404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12437_ _12443_/CLK _12437_/D vssd1 vssd1 vccd1 vccd1 _12437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12368_ _12369_/CLK _12368_/D vssd1 vssd1 vccd1 vccd1 _13497_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _14107_/A _08230_/X vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_114_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11319_ _11430_/A vssd1 vssd1 vccd1 vccd1 _11319_/X sky130_fd_sc_hd__buf_2
X_12299_ _12301_/CLK _12299_/D vssd1 vssd1 vccd1 vccd1 _13430_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_141_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14038_ _14038_/A _07882_/X vssd1 vssd1 vccd1 vccd1 _14070_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11277__B _13939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09970__B _10160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06860_ _06967_/A vssd1 vssd1 vccd1 vccd1 _06870_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06791_ _06801_/A _06793_/B _06793_/C vssd1 vssd1 vccd1 vccd1 _06792_/A sky130_fd_sc_hd__or3_1
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08530_ _08401_/X _08406_/X _08407_/X _08409_/X _08511_/X _08517_/X vssd1 vssd1 vccd1
+ vccd1 _08530_/X sky130_fd_sc_hd__mux4_1
XANTENNA__07490__B _08180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08461_ _09343_/C _09346_/C _12261_/Q _09352_/B _08445_/X _08446_/X vssd1 vssd1 vccd1
+ vccd1 _08461_/X sky130_fd_sc_hd__mux4_2
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07412_ _08131_/C vssd1 vssd1 vccd1 vccd1 _07423_/B sky130_fd_sc_hd__clkbuf_1
X_08392_ _13396_/A vssd1 vssd1 vccd1 vccd1 _08498_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07343_ _07343_/A vssd1 vssd1 vccd1 vccd1 _07343_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10637__A _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07274_ _07274_/A vssd1 vssd1 vccd1 vccd1 _07274_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10356__B _13756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09013_ _09030_/A vssd1 vssd1 vccd1 vccd1 _09013_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13948__A _13948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_1_clk_A _12917_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09915_ _13534_/A _09915_/B vssd1 vssd1 vccd1 vccd1 _09915_/X sky130_fd_sc_hd__or2_1
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09846_ _09846_/A vssd1 vssd1 vccd1 vccd1 _11151_/A sky130_fd_sc_hd__buf_8
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09777_ _09789_/B vssd1 vssd1 vccd1 vccd1 _09787_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_74_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06989_ _06995_/A _06995_/B vssd1 vssd1 vccd1 vccd1 _06990_/A sky130_fd_sc_hd__or2_1
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08728_ _08724_/X _08727_/X _09941_/A vssd1 vssd1 vccd1 vccd1 _09399_/D sky130_fd_sc_hd__mux2_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _12454_/Q _10111_/A _12456_/Q _12457_/Q _08578_/X _08579_/X vssd1 vssd1 vccd1
+ vccd1 _08659_/X sky130_fd_sc_hd__mux4_2
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11676_/A vssd1 vssd1 vccd1 vccd1 _11670_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09401__A _13596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10621_ _12581_/Q _13757_/A vssd1 vssd1 vccd1 vccd1 _10622_/D sky130_fd_sc_hd__xor2_1
XANTENNA__10959__A0 _13811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10552_ _10552_/A vssd1 vssd1 vccd1 vccd1 _10552_/X sky130_fd_sc_hd__buf_6
XFILLER_6_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10483_ _12543_/Q _13752_/A vssd1 vssd1 vccd1 vccd1 _10483_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12222_ _12325_/CLK _12222_/D vssd1 vssd1 vccd1 vccd1 _13399_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07856__A _08084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ _12153_/A vssd1 vssd1 vccd1 vccd1 _12967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _11124_/S vssd1 vssd1 vccd1 vccd1 _11118_/S sky130_fd_sc_hd__clkbuf_2
X_12084_ _12084_/A vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13593__A _13593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11035_ _10645_/X _11027_/X _11034_/X _11024_/X vssd1 vssd1 vccd1 vccd1 _12680_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13242__398 vssd1 vssd1 vccd1 vccd1 _13242__398/HI _13897_/A sky130_fd_sc_hd__conb_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11937_ _09623_/A _14034_/A _11940_/S vssd1 vssd1 vccd1 vccd1 _11938_/B sky130_fd_sc_hd__mux2_1
XFILLER_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11841__A _11852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11868_ _12893_/Q _14037_/A _11878_/S vssd1 vssd1 vccd1 vccd1 _11869_/B sky130_fd_sc_hd__mux2_1
X_13095__251 vssd1 vssd1 vccd1 vccd1 _13095__251/HI _13604_/A sky130_fd_sc_hd__conb_1
X_13607_ _13607_/A _07346_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
X_10819_ _10885_/A _10870_/D _10880_/C _10874_/B vssd1 vssd1 vccd1 vccd1 _10820_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11560__B _11604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11799_ _11799_/A _11799_/B vssd1 vssd1 vccd1 vccd1 _11800_/A sky130_fd_sc_hd__and2_1
XFILLER_158_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13538_ _13538_/A _07523_/X vssd1 vssd1 vccd1 vccd1 _13666_/Z sky130_fd_sc_hd__ebufn_8
X_13136__292 vssd1 vssd1 vccd1 vccd1 _13136__292/HI _13677_/A sky130_fd_sc_hd__conb_1
X_13469_ _13469_/A _07703_/X vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_145_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07961_ _07961_/A vssd1 vssd1 vccd1 vccd1 _07961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _09700_/A vssd1 vssd1 vccd1 vccd1 _12352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06912_ _06912_/A vssd1 vssd1 vccd1 vccd1 _06912_/X sky130_fd_sc_hd__clkbuf_1
X_07892_ _07892_/A vssd1 vssd1 vccd1 vccd1 _07903_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09631_ _09631_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09631_/X sky130_fd_sc_hd__or2_1
XFILLER_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06843_ _06850_/A _06843_/B _06843_/C vssd1 vssd1 vccd1 vccd1 _06844_/A sky130_fd_sc_hd__or3_1
XFILLER_95_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09562_ _13464_/A _12317_/Q _09575_/S vssd1 vssd1 vccd1 vccd1 _09563_/B sky130_fd_sc_hd__mux2_1
X_06774_ _06774_/A vssd1 vssd1 vccd1 vccd1 _06774_/X sky130_fd_sc_hd__clkbuf_1
X_08513_ _08443_/X _08447_/X _08452_/X _08455_/X _08511_/X _09157_/A vssd1 vssd1 vccd1
+ vccd1 _08513_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ _09967_/B vssd1 vssd1 vccd1 vccd1 _11929_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08444_ _12245_/Q vssd1 vssd1 vccd1 vccd1 _09328_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06845__A _07406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ _12232_/Q _12233_/Q _12234_/Q _09316_/C _08373_/X _08374_/X vssd1 vssd1 vccd1
+ vccd1 _08375_/X sky130_fd_sc_hd__mux4_1
X_07326_ _09875_/B vssd1 vssd1 vccd1 vccd1 _07473_/A sky130_fd_sc_hd__buf_2
XFILLER_149_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07257_ _07257_/A vssd1 vssd1 vccd1 vccd1 _07257_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07188_ _07188_/A vssd1 vssd1 vccd1 vccd1 _07188_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09891__A _10667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09829_ _09829_/A vssd1 vssd1 vccd1 vccd1 _12384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _12842_/CLK _12840_/D vssd1 vssd1 vccd1 vccd1 _12840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079__235 vssd1 vssd1 vccd1 vccd1 _13079__235/HI _13574_/A sky130_fd_sc_hd__conb_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12780_/CLK _12771_/D vssd1 vssd1 vccd1 vccd1 _12771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _12857_/Q _14002_/A _11726_/S vssd1 vssd1 vccd1 vccd1 _11723_/B sky130_fd_sc_hd__mux2_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06755__A _06809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09131__A _13391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11653_ _11657_/B _11652_/B _11569_/X vssd1 vssd1 vccd1 vccd1 _11655_/A sky130_fd_sc_hd__o21ai_1
XFILLER_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10604_ _10971_/A vssd1 vssd1 vccd1 vccd1 _10952_/A sky130_fd_sc_hd__buf_2
X_11584_ _12825_/Q vssd1 vssd1 vccd1 vccd1 _11631_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10535_ _13688_/A _10535_/B vssd1 vssd1 vccd1 vccd1 _10535_/X sky130_fd_sc_hd__or2_1
XFILLER_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10466_ _10466_/A vssd1 vssd1 vccd1 vccd1 _12544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12205_ _10670_/A _12195_/X _12204_/X _12200_/X vssd1 vssd1 vccd1 vccd1 _12979_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater123_A peripheralBus_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ _13652_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10397_/X sky130_fd_sc_hd__or2_1
XFILLER_151_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12136_ _12149_/A _12136_/B vssd1 vssd1 vccd1 vccd1 _12137_/A sky130_fd_sc_hd__and2_1
XFILLER_96_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12067_ _11160_/X _12061_/X _12066_/X _11497_/X vssd1 vssd1 vccd1 vccd1 _12938_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output52_A _13377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ _12661_/Q _13935_/A vssd1 vssd1 vccd1 vccd1 _11021_/B sky130_fd_sc_hd__xor2_1
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08210__A _08210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12085__A1 _10665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ _12969_/CLK _12969_/D vssd1 vssd1 vccd1 vccd1 _13375_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06490_ _06494_/A _06499_/B _06499_/C vssd1 vssd1 vccd1 vccd1 _06491_/A sky130_fd_sc_hd__or3_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09398__D _09848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08160_ _08174_/A _08174_/B _08164_/C vssd1 vssd1 vccd1 vccd1 _08161_/A sky130_fd_sc_hd__or3_4
XANTENNA__10399__A1 _10394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07111_ _07121_/A _07118_/B _07115_/C vssd1 vssd1 vccd1 vccd1 _07112_/A sky130_fd_sc_hd__or3_1
X_08091_ _08186_/A vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07042_ _07042_/A vssd1 vssd1 vccd1 vccd1 _07042_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08439__S1 _08418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_1_0_clk_A clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08993_ _11626_/A _11639_/C _11639_/B _12825_/Q _08946_/X _08947_/X vssd1 vssd1 vccd1
+ vccd1 _08993_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11746__A _11763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ _07944_/A vssd1 vssd1 vccd1 vccd1 _07944_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10650__A _10650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09216__A _09269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ _07881_/A _07877_/B _07877_/C vssd1 vssd1 vccd1 vccd1 _07876_/A sky130_fd_sc_hd__or3_1
XANTENNA__08120__A _08122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09614_ _09614_/A _09918_/B _12062_/A vssd1 vssd1 vccd1 vccd1 _09655_/B sky130_fd_sc_hd__or3_4
X_06826_ _06836_/A _06830_/B _07234_/C vssd1 vssd1 vccd1 vccd1 _06827_/A sky130_fd_sc_hd__or3_1
XFILLER_44_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09545_ _13459_/A _12312_/Q _09558_/S vssd1 vssd1 vccd1 vccd1 _09546_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06757_ _06757_/A vssd1 vssd1 vccd1 vccd1 _06757_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08375__S0 _08373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09476_ _12286_/Q _13562_/A vssd1 vssd1 vccd1 vccd1 _09478_/C sky130_fd_sc_hd__xnor2_1
X_06688_ _06688_/A vssd1 vssd1 vccd1 vccd1 _06748_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08427_ _09321_/D _12247_/Q _12248_/Q _09322_/A _08396_/X _08397_/X vssd1 vssd1 vccd1
+ vccd1 _08427_/X sky130_fd_sc_hd__mux4_2
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09886__A _13523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ _08358_/A _08358_/B _08360_/C vssd1 vssd1 vccd1 vccd1 _08359_/A sky130_fd_sc_hd__or3_1
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07309_ _07519_/A vssd1 vssd1 vccd1 vccd1 _07490_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ _08289_/A vssd1 vssd1 vccd1 vccd1 _08289_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10320_ _10320_/A vssd1 vssd1 vccd1 vccd1 _12507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07837__C _08180_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10251_ _11028_/B _11412_/C _10693_/C vssd1 vssd1 vccd1 vccd1 _10293_/B sky130_fd_sc_hd__nor3_4
XFILLER_3_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ _10182_/A vssd1 vssd1 vccd1 vccd1 _12471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14032__A _14032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13941_ _13941_/A _06444_/X vssd1 vssd1 vccd1 vccd1 _14069_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07572__C _08089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09180__A1 _10670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13872_ _13872_/A _06635_/X vssd1 vssd1 vccd1 vccd1 _14064_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__08965__A _11388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12067__A1 _11160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ _12823_/CLK _12823_/D vssd1 vssd1 vccd1 vccd1 _12823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12754_ _12758_/CLK _12754_/D vssd1 vssd1 vccd1 vccd1 _13881_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11705_/A _11705_/B _11705_/C _11705_/D vssd1 vssd1 vccd1 vccd1 _11709_/A
+ sky130_fd_sc_hd__or4_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12687_/CLK _12685_/D vssd1 vssd1 vccd1 vccd1 _13814_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11636_ _11634_/X _11682_/B _11636_/C vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__and3b_1
XFILLER_128_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11567_ _11565_/X _11604_/B _11567_/C vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__and3b_1
XFILLER_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10518_ _13681_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _10518_/X sky130_fd_sc_hd__or2_1
X_11498_ _13979_/A _11459_/A _11496_/X _11497_/X vssd1 vssd1 vccd1 vccd1 _12805_/D
+ sky130_fd_sc_hd__o211a_1
X_10449_ _10449_/A vssd1 vssd1 vccd1 vccd1 _12539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12119_ _12132_/A _12119_/B vssd1 vssd1 vccd1 vccd1 _12120_/A sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_41_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11285__B _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09171__A1 _10662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07660_ _07660_/A vssd1 vssd1 vccd1 vccd1 _07660_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_56_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06611_ _06611_/A vssd1 vssd1 vccd1 vccd1 _06611_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__12058__A1 _13376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07591_ _07601_/A _07598_/B _07593_/C vssd1 vssd1 vccd1 vccd1 _07592_/A sky130_fd_sc_hd__or3_1
XFILLER_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _09330_/A _09330_/B _09330_/C _09330_/D vssd1 vssd1 vccd1 vccd1 _09331_/D
+ sky130_fd_sc_hd__and4_1
X_06542_ _06694_/A vssd1 vssd1 vccd1 vccd1 _06604_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10629__B _13747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09261_ _09370_/A _09334_/C vssd1 vssd1 vccd1 vccd1 _09332_/B sky130_fd_sc_hd__and2_1
X_06473_ _06473_/A vssd1 vssd1 vccd1 vccd1 _06473_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08212_ _08212_/A _08222_/B _08212_/C vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__or3_1
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09192_ _12155_/A vssd1 vssd1 vccd1 vccd1 _09192_/X sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_114_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ _08143_/A vssd1 vssd1 vccd1 vccd1 _08143_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10645__A _10645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08074_ _08074_/A vssd1 vssd1 vccd1 vccd1 _08074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08115__A _11026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10364__B _13755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07025_ _07031_/A _07031_/B vssd1 vssd1 vccd1 vccd1 _07026_/A sky130_fd_sc_hd__or2_1
XFILLER_115_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09934__A0 _14034_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10380__A _11156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ _11641_/D _12830_/Q _12831_/Q _12832_/Q _08928_/X _08929_/X vssd1 vssd1 vccd1
+ vccd1 _08976_/X sky130_fd_sc_hd__mux4_2
XFILLER_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07927_ _07936_/A _07931_/B _07931_/C vssd1 vssd1 vccd1 vccd1 _07928_/A sky130_fd_sc_hd__or3_1
XFILLER_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07858_ _07858_/A vssd1 vssd1 vccd1 vccd1 _07858_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08785__A _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06809_ _06809_/A vssd1 vssd1 vccd1 vccd1 _07947_/B sky130_fd_sc_hd__clkbuf_2
X_07789_ _07817_/A vssd1 vssd1 vccd1 vccd1 _07801_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13041__197 vssd1 vssd1 vccd1 vccd1 _13041__197/HI _13484_/A sky130_fd_sc_hd__conb_1
X_09528_ _09846_/A vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__clkbuf_2
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09459_ _12279_/Q _13555_/A vssd1 vssd1 vccd1 vccd1 _09459_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12470_ _12470_/CLK _12470_/D vssd1 vssd1 vccd1 vccd1 _12470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11421_ _13906_/A _11423_/B vssd1 vssd1 vccd1 vccd1 _11421_/X sky130_fd_sc_hd__or2_1
XANTENNA__07848__B _07854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10555__A _13785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11352_ _11352_/A vssd1 vssd1 vccd1 vccd1 _12766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10303_ _10303_/A vssd1 vssd1 vccd1 vccd1 _12502_/D sky130_fd_sc_hd__clkbuf_1
X_14071_ _14071_/A _08015_/X vssd1 vssd1 vccd1 vccd1 _14103_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11283_ _11410_/A _11283_/B _11410_/C vssd1 vssd1 vccd1 vccd1 _11312_/A sky130_fd_sc_hd__or3_4
XFILLER_153_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10234_ _12480_/Q _13755_/A vssd1 vssd1 vccd1 vccd1 _10237_/B sky130_fd_sc_hd__xor2_1
XFILLER_105_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11386__A _12773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10165_ _10165_/A _10165_/B _10165_/C _10165_/D vssd1 vssd1 vccd1 vccd1 _10166_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_121_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10096_ _10096_/A vssd1 vssd1 vccd1 vccd1 _12451_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09153__A1 _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ _13924_/A _06491_/X vssd1 vssd1 vccd1 vccd1 _13988_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13855_ _13855_/A _06683_/X vssd1 vssd1 vccd1 vccd1 _13983_/Z sky130_fd_sc_hd__ebufn_8
X_12806_ _12806_/CLK _12806_/D vssd1 vssd1 vccd1 vccd1 _13980_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_34_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10998_ _10998_/A vssd1 vssd1 vccd1 vccd1 _12676_/D sky130_fd_sc_hd__clkbuf_1
X_13786_ _13786_/A _06876_/X vssd1 vssd1 vccd1 vccd1 _13978_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_43_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12753_/CLK _12737_/D vssd1 vssd1 vccd1 vccd1 _12737_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _12853_/CLK _12668_/D vssd1 vssd1 vccd1 vccd1 _12668_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06943__A _06955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ _11619_/A vssd1 vssd1 vccd1 vccd1 _12834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12599_ _12599_/CLK _12599_/D vssd1 vssd1 vccd1 vccd1 _13726_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11971__A0 _14108_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13776__A _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _10163_/D vssd1 vssd1 vccd1 vccd1 _13746_/A sky130_fd_sc_hd__buf_4
XFILLER_111_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08761_ _08750_/X _08759_/X _08863_/S vssd1 vssd1 vccd1 vccd1 _10163_/A sky130_fd_sc_hd__mux2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07712_ _09614_/A vssd1 vssd1 vccd1 vccd1 _07892_/A sky130_fd_sc_hd__buf_4
X_08692_ _08689_/X _08691_/X _08712_/S vssd1 vssd1 vccd1 vccd1 _09398_/C sky130_fd_sc_hd__mux2_1
XFILLER_38_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07643_ _08022_/A vssd1 vssd1 vccd1 vccd1 _07654_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07574_ _07615_/A vssd1 vssd1 vccd1 vccd1 _07585_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__10359__B _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ _09380_/A _09313_/B _09313_/C vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__and3_1
X_06525_ _06525_/A vssd1 vssd1 vccd1 vccd1 _06525_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_60_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _12821_/CLK sky130_fd_sc_hd__clkbuf_16
X_09244_ _09317_/B _09242_/C _09317_/A vssd1 vssd1 vccd1 vccd1 _09245_/C sky130_fd_sc_hd__a21o_1
X_06456_ _06548_/A _09102_/A _06548_/C _09096_/C vssd1 vssd1 vccd1 vccd1 _08210_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA__07949__A _08064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ input27/X vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12203__A1 _10665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06387_ _06391_/A _08349_/A vssd1 vssd1 vccd1 vccd1 _06388_/A sky130_fd_sc_hd__or2_1
XFILLER_147_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10375__A _11151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08502__S0 _08368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ _08135_/A _08128_/B _08138_/C vssd1 vssd1 vccd1 vccd1 _08127_/A sky130_fd_sc_hd__or3_1
XFILLER_135_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08057_ _08065_/A _08110_/B _08057_/C vssd1 vssd1 vccd1 vccd1 _08058_/A sky130_fd_sc_hd__or3_1
XFILLER_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07008_ _07008_/A vssd1 vssd1 vccd1 vccd1 _07008_/X sky130_fd_sc_hd__clkbuf_1
Xoutput37 _13404_/A vssd1 vssd1 vccd1 vccd1 pwm_en[3] sky130_fd_sc_hd__buf_2
XFILLER_134_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput48 _13952_/A vssd1 vssd1 vccd1 vccd1 pwm_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__11918__B _13363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10517__A1 _10385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput59 _13760_/A vssd1 vssd1 vccd1 vccd1 pwm_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__08805__S1 _08735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08959_ _12832_/Q _11641_/B _12834_/Q _12835_/Q _08928_/X _08929_/X vssd1 vssd1 vccd1
+ vccd1 _08959_/X sky130_fd_sc_hd__mux4_2
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11970_ _11970_/A vssd1 vssd1 vccd1 vccd1 _12916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09404__A _09404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10921_ _10921_/A _10921_/B _10921_/C vssd1 vssd1 vccd1 vccd1 _10922_/D sky130_fd_sc_hd__and3_1
XFILLER_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13640_ _13640_/A _07254_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
X_10852_ _10868_/D _10854_/C _10803_/X vssd1 vssd1 vccd1 vccd1 _10852_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13571_ _13571_/A _07441_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10790_/C _10783_/B vssd1 vssd1 vccd1 vccd1 _12623_/D sky130_fd_sc_hd__nor2_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _12699_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07859__A _07861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ _12522_/CLK _12522_/D vssd1 vssd1 vccd1 vccd1 _13651_/A sky130_fd_sc_hd__dfxtp_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12453_ _12461_/CLK _12453_/D vssd1 vssd1 vccd1 vccd1 _12453_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10285__A _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ _12764_/Q _13939_/A vssd1 vssd1 vccd1 vccd1 _11405_/D sky130_fd_sc_hd__xor2_1
XFILLER_138_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12384_ _12386_/CLK _12384_/D vssd1 vssd1 vccd1 vccd1 _12384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11335_ _11335_/A vssd1 vssd1 vccd1 vccd1 _12761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13596__A _13596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14123_ _14123_/A _08271_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
XFILLER_4_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11266_ _12733_/Q _13941_/A vssd1 vssd1 vccd1 vccd1 _11268_/C sky130_fd_sc_hd__xor2_1
X_14054_ _14054_/A _07926_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[23] sky130_fd_sc_hd__ebufn_8
XFILLER_98_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10732__B _10732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10217_ _13629_/A _12482_/Q _10220_/S vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__mux2_1
XFILLER_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11197_ _13853_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11197_/X sky130_fd_sc_hd__or2_1
XANTENNA__11181__A1 _10665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08202__B _08208_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10148_ _10148_/A _10148_/B _10148_/C vssd1 vssd1 vccd1 vccd1 _10149_/C sky130_fd_sc_hd__and3_1
XFILLER_79_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11844__A _11852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10079_ _10083_/B _10135_/B _10079_/C vssd1 vssd1 vccd1 vccd1 _10080_/A sky130_fd_sc_hd__and3b_1
XFILLER_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13907_ _13907_/A _06535_/X vssd1 vssd1 vccd1 vccd1 _14067_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13838_ _13838_/A _06730_/X vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__ebufn_8
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13769_ _13769_/A _06920_/X vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__ebufn_8
Xclkbuf_leaf_42_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _12565_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06310_ _11457_/B vssd1 vssd1 vccd1 vccd1 _06688_/A sky130_fd_sc_hd__buf_2
X_07290_ _07290_/A vssd1 vssd1 vccd1 vccd1 _07290_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07488__B _08180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11944__A0 peripheralBus_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09931_ _14033_/Z _08709_/X _09934_/S vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__mux2_1
XFILLER_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _12381_/Q _13558_/A vssd1 vssd1 vccd1 vccd1 _09863_/D sky130_fd_sc_hd__xor2_1
XFILLER_86_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater85_A _14065_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ _08800_/X _08802_/X _08805_/X _08809_/X _08810_/X _08812_/X vssd1 vssd1 vccd1
+ vccd1 _08813_/X sky130_fd_sc_hd__mux4_1
XANTENNA__07009__A _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _13519_/A _12374_/Q _09871_/B vssd1 vssd1 vccd1 vccd1 _09794_/B sky130_fd_sc_hd__mux2_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater120 peripheralBus_data[15] vssd1 vssd1 vccd1 vccd1 _14078_/Z sky130_fd_sc_hd__buf_12
Xrepeater131 _14106_/Z vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__buf_12
X_13304__460 vssd1 vssd1 vccd1 vccd1 _13304__460/HI _14025_/A sky130_fd_sc_hd__conb_1
XFILLER_85_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08744_ _12622_/Q _12623_/Q _12624_/Q _12625_/Q _08742_/X _08743_/X vssd1 vssd1 vccd1
+ vccd1 _08744_/X sky130_fd_sc_hd__mux4_2
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08675_ _08640_/X _08643_/X _08646_/X _08674_/X _08632_/X _08634_/X vssd1 vssd1 vccd1
+ vccd1 _08675_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _07630_/A _07626_/B _07635_/C vssd1 vssd1 vccd1 vccd1 _07627_/A sky130_fd_sc_hd__or3_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07557_ _07557_/A vssd1 vssd1 vccd1 vccd1 _07557_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_33_clk _12759_/CLK vssd1 vssd1 vccd1 vccd1 _12776_/CLK sky130_fd_sc_hd__clkbuf_16
X_06508_ _06508_/A vssd1 vssd1 vccd1 vccd1 _06508_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07488_ _07739_/A _08180_/B _08089_/B vssd1 vssd1 vccd1 vccd1 _07489_/A sky130_fd_sc_hd__or3_1
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06439_ _06913_/A vssd1 vssd1 vccd1 vccd1 _06449_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09227_ _09316_/C _09316_/D _09315_/C _09315_/D vssd1 vssd1 vccd1 vccd1 _09260_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09158_ _10652_/A _09145_/X _09157_/X _09148_/X vssd1 vssd1 vccd1 vccd1 _12218_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_135_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08109_ _08109_/A vssd1 vssd1 vccd1 vccd1 _08109_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11929__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ _09086_/X _09088_/X _09089_/S vssd1 vssd1 vccd1 vccd1 _10941_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11120_ _11120_/A vssd1 vssd1 vccd1 vccd1 _12707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _13816_/A _11051_/B vssd1 vssd1 vccd1 vccd1 _11051_/X sky130_fd_sc_hd__or2_1
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10002_ _10029_/D _10008_/D vssd1 vssd1 vccd1 vccd1 _10004_/A sky130_fd_sc_hd__and2_1
XFILLER_1_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10910__A1 _10872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07861__B _07962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input14_A peripheralBus_address[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _11953_/A vssd1 vssd1 vccd1 vccd1 _12911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10904_ _10936_/A _10904_/B _10904_/C vssd1 vssd1 vccd1 vccd1 _10905_/A sky130_fd_sc_hd__and3_1
XFILLER_60_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13353__509 vssd1 vssd1 vccd1 vccd1 _13353__509/HI _14122_/A sky130_fd_sc_hd__conb_1
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11884_ _11884_/A vssd1 vssd1 vccd1 vccd1 _12897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13623_ _13623_/A _07299_/X vssd1 vssd1 vccd1 vccd1 _13623_/Z sky130_fd_sc_hd__ebufn_8
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_10835_ _10833_/X _10917_/B _10835_/C vssd1 vssd1 vccd1 vccd1 _10836_/A sky130_fd_sc_hd__and3b_1
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_24_clk _12881_/CLK vssd1 vssd1 vccd1 vccd1 _12886_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _13554_/A _07483_/X vssd1 vssd1 vccd1 vccd1 _14034_/Z sky130_fd_sc_hd__ebufn_8
X_10766_ _10864_/D _10767_/C _10765_/Y vssd1 vssd1 vccd1 vccd1 _12620_/D sky130_fd_sc_hd__a21oi_1
Xrepeater67 _14070_/Z vssd1 vssd1 vccd1 vccd1 _14102_/Z sky130_fd_sc_hd__buf_12
Xrepeater78 _14098_/Z vssd1 vssd1 vccd1 vccd1 _14066_/Z sky130_fd_sc_hd__buf_12
Xrepeater89 peripheralBus_data[29] vssd1 vssd1 vccd1 vccd1 _14028_/Z sky130_fd_sc_hd__buf_12
X_12505_ _12505_/CLK _12505_/D vssd1 vssd1 vccd1 vccd1 _12505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13485_ _13485_/A _07660_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
X_10697_ _10697_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10697_/X sky130_fd_sc_hd__or2_1
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12436_ _12443_/CLK _12436_/D vssd1 vssd1 vccd1 vccd1 _12436_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11926__A0 _14063_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__A1 _10414_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12367_ _12367_/CLK _12367_/D vssd1 vssd1 vccd1 vccd1 _13496_/A sky130_fd_sc_hd__dfxtp_1
X_13247__403 vssd1 vssd1 vccd1 vccd1 _13247__403/HI _13902_/A sky130_fd_sc_hd__conb_1
XFILLER_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14106_ _14106_/A _08226_/X vssd1 vssd1 vccd1 vccd1 _14106_/Z sky130_fd_sc_hd__ebufn_8
X_11318_ _13883_/A _11323_/B vssd1 vssd1 vccd1 vccd1 _11318_/X sky130_fd_sc_hd__or2_1
XFILLER_141_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12298_ _12301_/CLK _12298_/D vssd1 vssd1 vccd1 vccd1 _13429_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11249_ _11255_/A _11249_/B vssd1 vssd1 vccd1 vccd1 _11250_/A sky130_fd_sc_hd__and2_1
X_14037_ _14037_/A _07878_/X vssd1 vssd1 vccd1 vccd1 _14037_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06790_ _06803_/A vssd1 vssd1 vccd1 vccd1 _06801_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__06668__A _06722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07490__C _07496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08460_ _12262_/Q vssd1 vssd1 vccd1 vccd1 _09352_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08883__A _10613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07411_ _09873_/B vssd1 vssd1 vccd1 vccd1 _08131_/C sky130_fd_sc_hd__buf_2
XANTENNA__08873__A3 _08872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08391_ _08386_/X _08388_/X _08389_/X _08390_/X _08382_/X _08383_/X vssd1 vssd1 vccd1
+ vccd1 _08391_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_15_clk _12217_/CLK vssd1 vssd1 vccd1 vccd1 _12980_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__07499__A _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07342_ _07342_/A _07351_/B _07347_/C vssd1 vssd1 vccd1 vccd1 _07343_/A sky130_fd_sc_hd__or3_1
XFILLER_148_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10637__B _10637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ _07279_/A _07276_/B _07273_/C vssd1 vssd1 vccd1 vccd1 _07274_/A sky130_fd_sc_hd__or3_1
XFILLER_148_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09012_ _13970_/A vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14125__A _14125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09914_ _09116_/X _09902_/X _09913_/X _09905_/X vssd1 vssd1 vccd1 vccd1 _12405_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09845_ _09845_/A vssd1 vssd1 vccd1 vccd1 _12389_/D sky130_fd_sc_hd__clkbuf_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A peripheralBus_address[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11484__A _11490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09776_ _09776_/A vssd1 vssd1 vccd1 vccd1 _09776_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06988_ _06988_/A vssd1 vssd1 vccd1 vccd1 _06988_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06578__A _08035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08727_ _08646_/X _08674_/X _08699_/X _08726_/X _08694_/X _08695_/X vssd1 vssd1 vccd1
+ vccd1 _08727_/X sky130_fd_sc_hd__mux4_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09889__A _09915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _08577_/X _08582_/X _08580_/X _08588_/X _08695_/A _08652_/X vssd1 vssd1 vccd1
+ vccd1 _08658_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _07609_/A vssd1 vssd1 vccd1 vccd1 _07609_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _12442_/Q vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10620_ _12570_/Q _13746_/A vssd1 vssd1 vccd1 vccd1 _10622_/C sky130_fd_sc_hd__xor2_1
XANTENNA__09274__B1 _09206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ _10548_/X _10538_/X _10549_/X _10550_/X vssd1 vssd1 vccd1 vccd1 _12565_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10482_ _10482_/A vssd1 vssd1 vccd1 vccd1 _12549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ _12903_/CLK _12221_/D vssd1 vssd1 vccd1 vccd1 _13398_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12152_ _12155_/A _12152_/B vssd1 vssd1 vccd1 vccd1 _12153_/A sky130_fd_sc_hd__and2_1
XFILLER_78_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11103_ _11103_/A vssd1 vssd1 vccd1 vccd1 _12702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13874__A _13874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12083_ _14071_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12083_/X sky130_fd_sc_hd__or2_1
XFILLER_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11034_ _13809_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11034_/X sky130_fd_sc_hd__or2_1
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11936_ _11936_/A vssd1 vssd1 vccd1 vccd1 _12906_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11867_ _11867_/A vssd1 vssd1 vccd1 vccd1 _12892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13606_ _13606_/A _07348_/X vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_8
X_10818_ _10840_/C vssd1 vssd1 vccd1 vccd1 _10833_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11798_ _09620_/A _14001_/A _11805_/S vssd1 vssd1 vccd1 vccd1 _11799_/B sky130_fd_sc_hd__mux2_1
X_13537_ _13537_/A _07525_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
X_10749_ _10803_/A vssd1 vssd1 vccd1 vccd1 _10749_/X sky130_fd_sc_hd__buf_2
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13468_ _13468_/A _07705_/X vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11569__A _11582_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12419_ _12420_/CLK _12419_/D vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__dfxtp_4
X_13399_ _13399_/A _07841_/X vssd1 vssd1 vccd1 vccd1 _13623_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07960_ _07983_/A _07971_/B _07962_/C vssd1 vssd1 vccd1 vccd1 _07961_/A sky130_fd_sc_hd__or3_1
XFILLER_114_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_4_clk _12917_/CLK vssd1 vssd1 vccd1 vccd1 _12914_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06911_ _08168_/A _06916_/B vssd1 vssd1 vccd1 vccd1 _06912_/A sky130_fd_sc_hd__or2_1
X_07891_ _07891_/A vssd1 vssd1 vccd1 vccd1 _07891_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09630_ _13460_/A _09627_/X _09629_/X _09621_/X vssd1 vssd1 vccd1 vccd1 _12330_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06842_ _06842_/A vssd1 vssd1 vccd1 vccd1 _06842_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09561_ _09582_/S vssd1 vssd1 vccd1 vccd1 _09575_/S sky130_fd_sc_hd__clkbuf_2
X_06773_ _06775_/A _06780_/B _06780_/C vssd1 vssd1 vccd1 vccd1 _06774_/A sky130_fd_sc_hd__or3_1
X_08512_ _08517_/A vssd1 vssd1 vccd1 vccd1 _09157_/A sky130_fd_sc_hd__buf_2
XFILLER_36_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09492_ _09623_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _09492_/X sky130_fd_sc_hd__or2_1
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09502__A _11170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ _09317_/A _12240_/Q _09315_/A _09316_/B _08368_/X _08370_/X vssd1 vssd1 vccd1
+ vccd1 _08443_/X sky130_fd_sc_hd__mux4_2
XANTENNA__10648__A _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ _08525_/A vssd1 vssd1 vccd1 vccd1 _08374_/X sky130_fd_sc_hd__buf_2
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08118__A _08122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07325_ _09918_/B vssd1 vssd1 vccd1 vccd1 _09875_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__07022__A _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07256_ _07266_/A _07263_/B _07260_/C vssd1 vssd1 vccd1 vccd1 _07257_/A sky130_fd_sc_hd__or3_1
XANTENNA__09875__C _11156_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07187_ _07193_/A _07190_/B _07187_/C vssd1 vssd1 vccd1 vccd1 _07188_/A sky130_fd_sc_hd__or3_1
XFILLER_145_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09828_ _09834_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__and2_1
XANTENNA__12103__A _13401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09759_ _09776_/A vssd1 vssd1 vccd1 vccd1 _09759_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12782_/CLK _12770_/D vssd1 vssd1 vccd1 vccd1 _12770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11721_/A vssd1 vssd1 vccd1 vccd1 _12856_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11652_/A _11652_/B _11515_/X vssd1 vssd1 vccd1 vccd1 _12839_/D sky130_fd_sc_hd__nor3b_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10603_ _10603_/A vssd1 vssd1 vccd1 vccd1 _12580_/D sky130_fd_sc_hd__clkbuf_1
X_11583_ _11583_/A vssd1 vssd1 vccd1 vccd1 _12824_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07867__A _07920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10534_ _09770_/X _10525_/X _10533_/X _10523_/X vssd1 vssd1 vccd1 vccd1 _12559_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10465_ _10477_/A _10465_/B vssd1 vssd1 vccd1 vccd1 _10466_/A sky130_fd_sc_hd__and2_1
XFILLER_108_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12204_ _14104_/A _12206_/B vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__or2_1
XFILLER_142_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10396_ _10423_/B vssd1 vssd1 vccd1 vccd1 _10406_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_108_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ _12962_/Q _14104_/A _12135_/S vssd1 vssd1 vccd1 vccd1 _12136_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater116_A peripheralBus_data[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12066_ _14064_/A _12073_/B vssd1 vssd1 vccd1 vccd1 _12066_/X sky130_fd_sc_hd__or2_1
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10740__B _10895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _12666_/Q _13940_/A vssd1 vssd1 vccd1 vccd1 _11021_/A sky130_fd_sc_hd__xor2_1
XFILLER_65_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output45_A _13761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11852__A _11852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12968_ _12968_/CLK _12968_/D vssd1 vssd1 vccd1 vccd1 _12968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_0_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11919_ _12887_/Q _13359_/A vssd1 vssd1 vccd1 vccd1 _11920_/D sky130_fd_sc_hd__xor2_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _12918_/CLK _12899_/D vssd1 vssd1 vccd1 vccd1 _12899_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07110_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07121_/A sky130_fd_sc_hd__clkbuf_1
X_08090_ _08090_/A vssd1 vssd1 vccd1 vccd1 _08090_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_158_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06681__A _06722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11299__A _11312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07041_ _07043_/A _07043_/B vssd1 vssd1 vccd1 vccd1 _07042_/A sky130_fd_sc_hd__or2_1
XFILLER_134_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08992_ _12824_/Q vssd1 vssd1 vccd1 vccd1 _11639_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07943_ _07951_/A _07945_/B _07945_/C vssd1 vssd1 vccd1 vccd1 _07944_/A sky130_fd_sc_hd__or3_1
XFILLER_96_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07874_ _07874_/A vssd1 vssd1 vccd1 vccd1 _07874_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08120__B _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09613_ _09640_/A vssd1 vssd1 vccd1 vccd1 _09613_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06825_ _06879_/A vssd1 vssd1 vccd1 vccd1 _06836_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _09582_/S vssd1 vssd1 vccd1 vccd1 _09558_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_70_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06756_ _06760_/A _06765_/B _06765_/C vssd1 vssd1 vccd1 vccd1 _06757_/A sky130_fd_sc_hd__or3_1
XFILLER_83_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08375__S1 _08374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09475_ _12277_/Q _13553_/A vssd1 vssd1 vccd1 vccd1 _09478_/B sky130_fd_sc_hd__xnor2_1
X_06687_ _06687_/A vssd1 vssd1 vccd1 vccd1 _06687_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10378__A _11156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08426_ _12249_/Q vssd1 vssd1 vccd1 vccd1 _09322_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13152__308 vssd1 vssd1 vccd1 vccd1 _13152__308/HI _13709_/A sky130_fd_sc_hd__conb_1
XFILLER_149_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08357_ _08357_/A vssd1 vssd1 vccd1 vccd1 _08357_/X sky130_fd_sc_hd__clkbuf_1
X_07308_ _07308_/A vssd1 vssd1 vccd1 vccd1 _07308_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08288_ _08288_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08289_/A sky130_fd_sc_hd__or2_1
XFILLER_109_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07239_ _07239_/A _07250_/B _07246_/C vssd1 vssd1 vccd1 vccd1 _07240_/A sky130_fd_sc_hd__or3_1
XFILLER_152_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10250_ _10250_/A vssd1 vssd1 vccd1 vccd1 _11412_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10181_ _10191_/A _10181_/B vssd1 vssd1 vccd1 vccd1 _10182_/A sky130_fd_sc_hd__and2_1
X_13046__202 vssd1 vssd1 vccd1 vccd1 _13046__202/HI _13505_/A sky130_fd_sc_hd__conb_1
XFILLER_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09407__A _11408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08311__A _08335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _13940_/A _06446_/X vssd1 vssd1 vccd1 vccd1 _14068_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__09126__B input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13871_ _13871_/A _07858_/X vssd1 vssd1 vccd1 vccd1 _14063_/Z sky130_fd_sc_hd__ebufn_8
X_12822_ _12823_/CLK _12822_/D vssd1 vssd1 vccd1 vccd1 _12822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11391__B _13945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12753_ _12753_/CLK _12753_/D vssd1 vssd1 vccd1 vccd1 _13880_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10288__A _11064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11704_/A vssd1 vssd1 vccd1 vccd1 _12853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12806_/CLK _12684_/D vssd1 vssd1 vccd1 vccd1 _13813_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ _11640_/A _11622_/B _11639_/A vssd1 vssd1 vccd1 vccd1 _11636_/C sky130_fd_sc_hd__a21o_1
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11566_ _11563_/A _11572_/C _11626_/B vssd1 vssd1 vccd1 vccd1 _11567_/C sky130_fd_sc_hd__a21o_1
XFILLER_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10517_ _10385_/X _10511_/X _10516_/X _10425_/X vssd1 vssd1 vccd1 vccd1 _12552_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11497_ _12084_/A vssd1 vssd1 vccd1 vccd1 _11497_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10448_ _10461_/A _10448_/B vssd1 vssd1 vccd1 vccd1 _10449_/A sky130_fd_sc_hd__and2_1
XFILLER_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11847__A _11898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10379_ _10409_/A vssd1 vssd1 vccd1 vccd1 _10379_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12118_ _12957_/Q _14099_/A _12118_/S vssd1 vssd1 vccd1 vccd1 _12119_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11285__C _11412_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12049_ _12932_/Q _13371_/A vssd1 vssd1 vccd1 vccd1 _12050_/D sky130_fd_sc_hd__xor2_1
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06610_ _06610_/A _06616_/B _06616_/C vssd1 vssd1 vccd1 vccd1 _06611_/A sky130_fd_sc_hd__or3_1
X_07590_ _07590_/A vssd1 vssd1 vccd1 vccd1 _07601_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__06676__A _06686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12058__A2 _12057_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06541_ _06541_/A vssd1 vssd1 vccd1 vccd1 _06541_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09260_ _09318_/A _09260_/B _09260_/C _09260_/D vssd1 vssd1 vccd1 vccd1 _09334_/C
+ sky130_fd_sc_hd__and4_2
X_06472_ _06481_/A _07827_/B _06472_/C vssd1 vssd1 vccd1 vccd1 _06473_/A sky130_fd_sc_hd__or3_1
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08211_ _08263_/A vssd1 vssd1 vccd1 vccd1 _08222_/B sky130_fd_sc_hd__clkbuf_1
X_09191_ _13404_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _09191_/X sky130_fd_sc_hd__or2_1
XFILLER_159_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08142_ _08148_/A _08151_/B _08151_/C vssd1 vssd1 vccd1 vccd1 _08143_/A sky130_fd_sc_hd__or3_1
X_08073_ _08081_/A _08077_/B _08087_/C vssd1 vssd1 vccd1 vccd1 _08074_/A sky130_fd_sc_hd__or3_1
XFILLER_162_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07024_ _07024_/A vssd1 vssd1 vccd1 vccd1 _07024_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08131__A _08135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _12825_/Q _12826_/Q _12827_/Q _11632_/A _08915_/X _08916_/X vssd1 vssd1 vccd1
+ vccd1 _08975_/X sky130_fd_sc_hd__mux4_2
XANTENNA__10380__B _11412_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07926_ _07926_/A vssd1 vssd1 vccd1 vccd1 _07926_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07857_ _07857_/A _07962_/B _07995_/B vssd1 vssd1 vccd1 vccd1 _07858_/A sky130_fd_sc_hd__or3_1
XANTENNA__11492__A _14009_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06808_ _06832_/A vssd1 vssd1 vccd1 vccd1 _06830_/B sky130_fd_sc_hd__clkbuf_1
X_07788_ _07788_/A vssd1 vssd1 vccd1 vccd1 _07788_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09527_ _13438_/A _09513_/A _09526_/X _09522_/X vssd1 vssd1 vccd1 vccd1 _12307_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06739_ _06739_/A vssd1 vssd1 vccd1 vccd1 _06739_/X sky130_fd_sc_hd__clkbuf_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09458_ _12276_/Q _13552_/A vssd1 vssd1 vccd1 vccd1 _09468_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09870__B1 _13567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08409_ _12253_/Q _09320_/D _12255_/Q _12256_/Q _08379_/X _08380_/X vssd1 vssd1 vccd1
+ vccd1 _08409_/X sky130_fd_sc_hd__mux4_2
X_09389_ _09389_/A _09389_/B _09391_/B vssd1 vssd1 vccd1 vccd1 _09390_/A sky130_fd_sc_hd__and3_1
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11420_ _10645_/X _11411_/X _11419_/X _11417_/X vssd1 vssd1 vccd1 vccd1 _12779_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11351_ _11361_/A _11351_/B vssd1 vssd1 vccd1 vccd1 _11352_/A sky130_fd_sc_hd__and2_1
XFILLER_152_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10302_ _10315_/A _10302_/B vssd1 vssd1 vccd1 vccd1 _10303_/A sky130_fd_sc_hd__and2_1
X_14070_ _14070_/A _08011_/X vssd1 vssd1 vccd1 vccd1 _14070_/Z sky130_fd_sc_hd__ebufn_8
X_11282_ _11282_/A vssd1 vssd1 vccd1 vccd1 _12743_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09386__C1 _09263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ _12483_/Q _13758_/A vssd1 vssd1 vccd1 vccd1 _10237_/A sky130_fd_sc_hd__xor2_1
XFILLER_161_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10164_ _10164_/A _10164_/B _10164_/C _10613_/B vssd1 vssd1 vccd1 vccd1 _10166_/C
+ sky130_fd_sc_hd__or4_1
XANTENNA__08041__A _08067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13280__436 vssd1 vssd1 vccd1 vccd1 _13280__436/HI _13985_/A sky130_fd_sc_hd__conb_1
XFILLER_94_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10095_ _10146_/A _10095_/B _10095_/C vssd1 vssd1 vccd1 vccd1 _10096_/A sky130_fd_sc_hd__and3_1
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07880__A _07920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13923_ _13923_/A _06493_/X vssd1 vssd1 vccd1 vccd1 _13987_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13321__477 vssd1 vssd1 vccd1 vccd1 _13321__477/HI _14058_/A sky130_fd_sc_hd__conb_1
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13854_ _13854_/A _06685_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
X_12805_ _12806_/CLK _12805_/D vssd1 vssd1 vccd1 vccd1 _13979_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13785_ _13785_/A _06878_/X vssd1 vssd1 vccd1 vccd1 _14105_/Z sky130_fd_sc_hd__ebufn_8
X_10997_ _11078_/A _10997_/B vssd1 vssd1 vccd1 vccd1 _10998_/A sky130_fd_sc_hd__and2_1
XFILLER_43_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12736_ _12753_/CLK _12736_/D vssd1 vssd1 vccd1 vccd1 _12736_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13174__330 vssd1 vssd1 vccd1 vccd1 _13174__330/HI _13767_/A sky130_fd_sc_hd__conb_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _12853_/CLK _12667_/D vssd1 vssd1 vccd1 vccd1 _12667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11618_ _11622_/B _11682_/B _11618_/C vssd1 vssd1 vccd1 vccd1 _11619_/A sky130_fd_sc_hd__and3b_1
X_12598_ _12598_/CLK _12598_/D vssd1 vssd1 vccd1 vccd1 _13725_/A sky130_fd_sc_hd__dfxtp_1
X_13215__371 vssd1 vssd1 vccd1 vccd1 _13215__371/HI _13838_/A sky130_fd_sc_hd__conb_1
XFILLER_144_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11549_ _11627_/B _11563_/A vssd1 vssd1 vccd1 vccd1 _11550_/C sky130_fd_sc_hd__or2_1
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08760_ _13780_/A vssd1 vssd1 vccd1 vccd1 _08863_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_112_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ _07711_/A vssd1 vssd1 vccd1 vccd1 _07711_/X sky130_fd_sc_hd__clkbuf_1
X_08691_ _08617_/X _08619_/X _08666_/X _08690_/X _08678_/X _08647_/X vssd1 vssd1 vccd1
+ vccd1 _08691_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07642_ _07642_/A vssd1 vssd1 vccd1 vccd1 _07642_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07573_ _07573_/A vssd1 vssd1 vccd1 vccd1 _07573_/X sky130_fd_sc_hd__clkbuf_1
X_09312_ _09329_/A _09312_/B vssd1 vssd1 vccd1 vccd1 _09313_/C sky130_fd_sc_hd__nand2_1
X_06524_ _06534_/A _06526_/B _06526_/C vssd1 vssd1 vccd1 vccd1 _06525_/A sky130_fd_sc_hd__or3_1
XFILLER_34_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09243_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09389_/A sky130_fd_sc_hd__buf_2
X_06455_ input18/X vssd1 vssd1 vccd1 vccd1 _06548_/A sky130_fd_sc_hd__inv_2
XANTENNA__10656__A _10686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11251__S _11254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06386_ _06386_/A vssd1 vssd1 vccd1 vccd1 _06386_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09174_ _13399_/A _09179_/B vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__and2_1
XANTENNA__08126__A _08135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08502__S1 _08370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ _08153_/A vssd1 vssd1 vccd1 vccd1 _08138_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__13967__A _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07965__A _08084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _08056_/A vssd1 vssd1 vccd1 vccd1 _08056_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07007_ _07007_/A _07007_/B vssd1 vssd1 vccd1 vccd1 _07008_/A sky130_fd_sc_hd__or2_1
XANTENNA__11487__A _11490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput38 _13593_/A vssd1 vssd1 vccd1 vccd1 pwm_en[4] sky130_fd_sc_hd__buf_2
Xoutput49 _13953_/A vssd1 vssd1 vccd1 vccd1 pwm_out[14] sky130_fd_sc_hd__buf_2
XFILLER_115_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08958_ _12833_/Q vssd1 vssd1 vccd1 vccd1 _11641_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07909_ _07909_/A vssd1 vssd1 vccd1 vccd1 _07909_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08889_ _08757_/X _08833_/X _08861_/X _08888_/X _08810_/X _08812_/X vssd1 vssd1 vccd1
+ vccd1 _08889_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10920_ _10921_/B _10915_/X _10919_/Y vssd1 vssd1 vccd1 vccd1 _12655_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__07205__A _07205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158__314 vssd1 vssd1 vccd1 vccd1 _13158__314/HI _13731_/A sky130_fd_sc_hd__conb_1
XFILLER_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ _10876_/B vssd1 vssd1 vccd1 vccd1 _10868_/D sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _13570_/A _07443_/X vssd1 vssd1 vccd1 vccd1 _13666_/Z sky130_fd_sc_hd__ebufn_8
X_10782_ _10865_/C _10780_/B _10781_/X vssd1 vssd1 vccd1 vccd1 _10783_/B sky130_fd_sc_hd__o21ai_1
XFILLER_52_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12522_/CLK _12521_/D vssd1 vssd1 vccd1 vccd1 _13650_/A sky130_fd_sc_hd__dfxtp_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07859__B _07962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _12457_/CLK _12452_/D vssd1 vssd1 vccd1 vccd1 _12452_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08036__A _11283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ _12768_/Q _13943_/A vssd1 vssd1 vccd1 vccd1 _11405_/C sky130_fd_sc_hd__xor2_1
XFILLER_126_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12383_ _12400_/CLK _12383_/D vssd1 vssd1 vccd1 vccd1 _12383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14122_ _14122_/A _08269_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
X_11334_ _11344_/A _11334_/B vssd1 vssd1 vccd1 vccd1 _11335_/A sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_55_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14053_ _14053_/A _07922_/X vssd1 vssd1 vccd1 vccd1 _14117_/Z sky130_fd_sc_hd__ebufn_8
X_11265_ _12741_/Q _13949_/A vssd1 vssd1 vccd1 vccd1 _11268_/B sky130_fd_sc_hd__xor2_1
XFILLER_106_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10216_ _10216_/A vssd1 vssd1 vccd1 vccd1 _12481_/D sky130_fd_sc_hd__clkbuf_1
X_11196_ _11064_/X _11185_/X _11194_/X _11195_/X vssd1 vssd1 vccd1 vccd1 _12724_/D
+ sky130_fd_sc_hd__o211a_1
X_10147_ _10147_/A vssd1 vssd1 vccd1 vccd1 _12463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_113_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ _10099_/B _10086_/B _10076_/D _10099_/A vssd1 vssd1 vccd1 vccd1 _10079_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13906_ _13906_/A _06539_/X vssd1 vssd1 vccd1 vccd1 _14066_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10141__B1 _09978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ _13837_/A _06732_/X vssd1 vssd1 vccd1 vccd1 _14125_/Z sky130_fd_sc_hd__ebufn_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13768_ _13768_/A _06922_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_43_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12719_ _12722_/CLK _12719_/D vssd1 vssd1 vccd1 vccd1 _13847_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_13699_ _13699_/A _07095_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07488__C _08089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13787__A _13787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09930_ _09139_/X _09921_/X _09929_/X _09916_/X vssd1 vssd1 vccd1 vccd1 _12408_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _12389_/Q _13566_/A vssd1 vssd1 vccd1 vccd1 _09863_/C sky130_fd_sc_hd__xor2_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _08876_/A vssd1 vssd1 vccd1 vccd1 _08812_/X sky130_fd_sc_hd__clkbuf_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _09843_/S vssd1 vssd1 vccd1 vccd1 _09871_/B sky130_fd_sc_hd__buf_2
Xrepeater110 peripheralBus_data[1] vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__buf_12
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater121 peripheralBus_data[15] vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__buf_12
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater132 peripheralBus_data[11] vssd1 vssd1 vccd1 vccd1 _14106_/Z sky130_fd_sc_hd__buf_12
XFILLER_85_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater78_A _14098_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08743_ _13777_/A vssd1 vssd1 vccd1 vccd1 _08743_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07951__C _07962_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _10130_/D _12457_/Q _10130_/B _10130_/A _08602_/X _08603_/X vssd1 vssd1 vccd1
+ vccd1 _08674_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08420__S0 _08373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07625_ _07625_/A vssd1 vssd1 vccd1 vccd1 _07625_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10683__A1 _10288_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07556_ _07558_/A _07558_/B _07564_/C vssd1 vssd1 vccd1 vccd1 _07557_/A sky130_fd_sc_hd__or3_1
X_06507_ _06507_/A _06512_/B _06512_/C vssd1 vssd1 vccd1 vccd1 _06508_/A sky130_fd_sc_hd__or3_1
X_07487_ _07487_/A vssd1 vssd1 vccd1 vccd1 _07487_/X sky130_fd_sc_hd__clkbuf_1
X_09226_ _09226_/A _09226_/B vssd1 vssd1 vccd1 vccd1 _12234_/D sky130_fd_sc_hd__nor2_1
XFILLER_42_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06438_ _06438_/A vssd1 vssd1 vccd1 vccd1 _06438_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12188__A1 _10645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09157_ _09157_/A _09179_/B vssd1 vssd1 vccd1 vccd1 _09157_/X sky130_fd_sc_hd__and2_1
XFILLER_108_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06369_ _06822_/A _07822_/B _07822_/C vssd1 vssd1 vccd1 vccd1 _06370_/A sky130_fd_sc_hd__or3_1
XFILLER_108_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08108_ _08110_/A _08113_/B _08122_/C vssd1 vssd1 vccd1 vccd1 _08109_/A sky130_fd_sc_hd__or3_1
XFILLER_135_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09088_ _09008_/X _09036_/X _09061_/X _09087_/X _09056_/X _09057_/X vssd1 vssd1 vccd1
+ vccd1 _09088_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08039_ _08039_/A _08047_/B _08044_/C vssd1 vssd1 vccd1 vccd1 _08040_/A sky130_fd_sc_hd__or3_1
XFILLER_123_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11050_ _10665_/X _11041_/X _11049_/X _11039_/X vssd1 vssd1 vccd1 vccd1 _12686_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10001_ _12429_/Q vssd1 vssd1 vccd1 vccd1 _10029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07861__C _07947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09134__B _11460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11952_ _11962_/A _11952_/B vssd1 vssd1 vccd1 vccd1 _11953_/A sky130_fd_sc_hd__and2_1
XANTENNA__11320__C1 _11319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _10907_/B _10903_/B vssd1 vssd1 vccd1 vccd1 _10904_/C sky130_fd_sc_hd__nand2_1
XFILLER_45_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11883_ _11886_/A _11883_/B vssd1 vssd1 vccd1 vccd1 _11884_/A sky130_fd_sc_hd__and2_1
XANTENNA__11680__A _11680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13622_ _13622_/A _07301_/X vssd1 vssd1 vccd1 vccd1 _13974_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10834_ _10870_/B _10828_/A _10870_/A vssd1 vssd1 vccd1 vccd1 _10835_/C sky130_fd_sc_hd__a21o_1
XFILLER_25_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09150__A _14066_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10426__A1 _09120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13553_ _13553_/A _07485_/X vssd1 vssd1 vccd1 vccd1 _14033_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10765_ _10864_/D _10767_/C _10757_/X vssd1 vssd1 vccd1 vccd1 _10765_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater68 peripheralBus_data[7] vssd1 vssd1 vccd1 vccd1 _14070_/Z sky130_fd_sc_hd__buf_12
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ _12505_/CLK _12504_/D vssd1 vssd1 vccd1 vccd1 _12504_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater79 _14034_/Z vssd1 vssd1 vccd1 vccd1 _14098_/Z sky130_fd_sc_hd__buf_12
XFILLER_40_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13484_ _13484_/A _07663_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_40_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10696_ _10377_/X _10690_/X _10695_/X _10682_/X vssd1 vssd1 vccd1 vccd1 _12600_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12179__A1 _13375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12435_ _12443_/CLK _12435_/D vssd1 vssd1 vccd1 vccd1 _12435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12366_ _12367_/CLK _12366_/D vssd1 vssd1 vccd1 vccd1 _13495_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13286__442 vssd1 vssd1 vccd1 vccd1 _13286__442/HI _13991_/A sky130_fd_sc_hd__conb_1
XFILLER_114_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14105_ _14105_/A _08223_/X vssd1 vssd1 vccd1 vccd1 _14105_/Z sky130_fd_sc_hd__ebufn_8
X_11317_ _11189_/X _11312_/X _11316_/X _11306_/X vssd1 vssd1 vccd1 vccd1 _12755_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12297_ _12301_/CLK _12297_/D vssd1 vssd1 vccd1 vccd1 _13428_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12016__A _12033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14036_ _14036_/A _07876_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[5] sky130_fd_sc_hd__ebufn_8
X_11248_ _13884_/A _12740_/Q _11248_/S vssd1 vssd1 vccd1 vccd1 _11249_/B sky130_fd_sc_hd__mux2_1
X_13327__483 vssd1 vssd1 vccd1 vccd1 _13327__483/HI _14080_/A sky130_fd_sc_hd__conb_1
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11179_ _13847_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11179_/X sky130_fd_sc_hd__or2_1
XFILLER_121_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07410_ _09918_/B vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__buf_2
XANTENNA__09807__A0 _13523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08390_ _12256_/Q _12257_/Q _12258_/Q _12259_/Q _08379_/X _08380_/X vssd1 vssd1 vccd1
+ vccd1 _08390_/X sky130_fd_sc_hd__mux4_2
XANTENNA__06684__A _06686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11614__B1 _11505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07341_ _07341_/A vssd1 vssd1 vccd1 vccd1 _07341_/X sky130_fd_sc_hd__clkbuf_1
X_07272_ _07272_/A vssd1 vssd1 vccd1 vccd1 _07272_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09011_ _10939_/D vssd1 vssd1 vccd1 vccd1 _13938_/A sky130_fd_sc_hd__buf_4
XFILLER_117_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09913_ _13533_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09913_/X sky130_fd_sc_hd__or2_1
XFILLER_59_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09844_ _10173_/A _09844_/B vssd1 vssd1 vccd1 vccd1 _09845_/A sky130_fd_sc_hd__and2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07962__B _07962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06859__A _06900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _09773_/X _09759_/X _09774_/X _09765_/X vssd1 vssd1 vccd1 vccd1 _12367_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06987_ _06995_/A _06995_/B vssd1 vssd1 vccd1 vccd1 _06988_/A sky130_fd_sc_hd__or2_1
XANTENNA__13980__A _13980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ _10149_/A _10155_/B _12466_/Q _12467_/Q _09929_/A _08709_/X vssd1 vssd1 vccd1
+ vccd1 _08726_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _09867_/B vssd1 vssd1 vccd1 vccd1 _13555_/A sky130_fd_sc_hd__buf_4
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _07616_/A _07613_/B _07608_/C vssd1 vssd1 vccd1 vccd1 _07609_/A sky130_fd_sc_hd__or3_1
X_13120__276 vssd1 vssd1 vccd1 vccd1 _13120__276/HI _13645_/A sky130_fd_sc_hd__conb_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _10097_/B _12439_/Q _10052_/C _12441_/Q _08578_/X _08579_/X vssd1 vssd1 vccd1
+ vccd1 _08588_/X sky130_fd_sc_hd__mux4_2
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07539_ _07539_/A vssd1 vssd1 vccd1 vccd1 _07539_/X sky130_fd_sc_hd__clkbuf_1
X_10550_ _10650_/A vssd1 vssd1 vccd1 vccd1 _10550_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _09370_/A vssd1 vssd1 vccd1 vccd1 _09347_/A sky130_fd_sc_hd__buf_2
X_10481_ _10567_/A _10481_/B vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__and2_1
XFILLER_136_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12220_ _12903_/CLK _12220_/D vssd1 vssd1 vccd1 vccd1 _13397_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13014__170 vssd1 vssd1 vccd1 vccd1 _13014__170/HI _13441_/A sky130_fd_sc_hd__conb_1
XFILLER_163_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12151_ _12967_/Q _14109_/A _12151_/S vssd1 vssd1 vccd1 vccd1 _12152_/B sky130_fd_sc_hd__mux2_1
XFILLER_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11102_ _11112_/A _11102_/B vssd1 vssd1 vccd1 vccd1 _11103_/A sky130_fd_sc_hd__and2_1
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12082_ _10662_/A _12075_/X _12081_/X _12071_/X vssd1 vssd1 vccd1 vccd1 _12944_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11033_ _10385_/X _11027_/X _11032_/X _11024_/X vssd1 vssd1 vccd1 vccd1 _12679_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11394__B _13938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10647__A1 _10645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11935_ _11945_/A _11935_/B vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__and2_1
XFILLER_91_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11866_ _11869_/A _11866_/B vssd1 vssd1 vccd1 vccd1 _11867_/A sky130_fd_sc_hd__and2_1
XFILLER_72_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13605_ _13605_/A _07352_/X vssd1 vssd1 vccd1 vccd1 _13765_/Z sky130_fd_sc_hd__ebufn_8
X_10817_ _13775_/A _10874_/B _10870_/D _10880_/C vssd1 vssd1 vccd1 vccd1 _10840_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__08699__S0 _08602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11797_ _11797_/A vssd1 vssd1 vccd1 vccd1 _12872_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08208__B _08208_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13536_ _13536_/A _07528_/X vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__ebufn_8
X_10748_ _10768_/A vssd1 vssd1 vccd1 vccd1 _10803_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13467_ _13467_/A _07709_/X vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__ebufn_8
X_10679_ _13723_/A _10684_/B vssd1 vssd1 vccd1 vccd1 _10679_/X sky130_fd_sc_hd__or2_1
XFILLER_145_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12418_ _12418_/CLK _12418_/D vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_126_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13398_ _13398_/A _08361_/X vssd1 vssd1 vccd1 vccd1 _14102_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__08224__A _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _12349_/CLK _12349_/D vssd1 vssd1 vccd1 vccd1 _12349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14019_ _14019_/A _08069_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
X_06910_ _06910_/A vssd1 vssd1 vccd1 vccd1 _06910_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07890_ _07894_/A _07890_/B _07890_/C vssd1 vssd1 vccd1 vccd1 _07891_/A sky130_fd_sc_hd__or3_1
X_13063__219 vssd1 vssd1 vccd1 vccd1 _13063__219/HI _13538_/A sky130_fd_sc_hd__conb_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06841_ _06850_/A _06843_/B _06843_/C vssd1 vssd1 vccd1 vccd1 _06842_/A sky130_fd_sc_hd__or3_1
XFILLER_95_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09560_ _09560_/A vssd1 vssd1 vccd1 vccd1 _12316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06772_ _06772_/A vssd1 vssd1 vccd1 vccd1 _06772_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08511_ _13394_/A vssd1 vssd1 vccd1 vccd1 _08511_/X sky130_fd_sc_hd__buf_2
X_09491_ _13425_/A _09483_/X _09490_/X _09192_/X vssd1 vssd1 vccd1 vccd1 _12294_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08442_ _12242_/Q vssd1 vssd1 vccd1 vccd1 _09316_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08373_ _08524_/A vssd1 vssd1 vccd1 vccd1 _08373_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11063__A1 _11061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07324_ _07324_/A vssd1 vssd1 vccd1 vccd1 _07324_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07255_ _07281_/A vssd1 vssd1 vccd1 vccd1 _07266_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_117_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07186_ _07186_/A vssd1 vssd1 vccd1 vccd1 _07186_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10023__C1 _09987_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__C1 _09959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09827_ _13529_/A _12384_/Q _09837_/S vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__mux2_1
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09758_ _09756_/X _09741_/X _09757_/X _09748_/X vssd1 vssd1 vccd1 vccd1 _12362_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ _08709_/A vssd1 vssd1 vccd1 vccd1 _08709_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _10988_/A vssd1 vssd1 vccd1 vccd1 _09836_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11723_/A _11720_/B vssd1 vssd1 vccd1 vccd1 _11721_/A sky130_fd_sc_hd__and2_1
XFILLER_70_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11658_/A _11657_/C _11688_/B vssd1 vssd1 vccd1 vccd1 _11652_/B sky130_fd_sc_hd__and3_1
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11054__A1 _10670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ _10602_/A _10602_/B vssd1 vssd1 vccd1 vccd1 _10603_/A sky130_fd_sc_hd__and2_1
XFILLER_23_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11582_ _11595_/A _11582_/B _11582_/C vssd1 vssd1 vccd1 vccd1 _11583_/A sky130_fd_sc_hd__and3b_1
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10533_ _13687_/A _10535_/B vssd1 vssd1 vccd1 vccd1 _10533_/X sky130_fd_sc_hd__or2_1
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11389__B _13946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ _13689_/A _12544_/Q _10473_/S vssd1 vssd1 vccd1 vccd1 _10465_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10293__B _10293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12203_ _10665_/A _12195_/X _12202_/X _12200_/X vssd1 vssd1 vccd1 vccd1 _12978_/D
+ sky130_fd_sc_hd__o211a_1
X_10395_ _10409_/A vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07883__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ _12134_/A vssd1 vssd1 vccd1 vccd1 _12149_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12065_ _11153_/X _12061_/X _12064_/X _11497_/X vssd1 vssd1 vccd1 vccd1 _12937_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater109_A _13616_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11016_ _11016_/A _11016_/B _11016_/C _11016_/D vssd1 vssd1 vccd1 vccd1 _11022_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output38_A _13593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12967_ _12968_/CLK _12967_/D vssd1 vssd1 vccd1 vccd1 _12967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11918_ _12891_/Q _13363_/A vssd1 vssd1 vccd1 vccd1 _11920_/C sky130_fd_sc_hd__xor2_1
XFILLER_73_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ _12914_/CLK _12898_/D vssd1 vssd1 vccd1 vccd1 _12898_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11849_ _11852_/A _11849_/B vssd1 vssd1 vccd1 vccd1 _11850_/A sky130_fd_sc_hd__and2_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13519_ _13519_/A _08104_/X vssd1 vssd1 vccd1 vccd1 _13775_/Z sky130_fd_sc_hd__ebufn_8
X_07040_ _07040_/A vssd1 vssd1 vccd1 vccd1 _07040_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__07496__C _07496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08991_ _11562_/C _11625_/B _11625_/A _11626_/B _08911_/X _08913_/X vssd1 vssd1 vccd1
+ vccd1 _08991_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07942_ _07942_/A vssd1 vssd1 vccd1 vccd1 _07942_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07873_ _07881_/A _07877_/B _07877_/C vssd1 vssd1 vccd1 vccd1 _07874_/A sky130_fd_sc_hd__or3_1
X_09612_ _11154_/B _09873_/B _10637_/B vssd1 vssd1 vccd1 vccd1 _09640_/A sky130_fd_sc_hd__nor3_4
XANTENNA__08120__C _08131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06824_ _09125_/A vssd1 vssd1 vccd1 vccd1 _06879_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater60_A _14072_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__A _09513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ _09543_/A vssd1 vssd1 vccd1 vccd1 _12311_/D sky130_fd_sc_hd__clkbuf_1
X_06755_ _06809_/A vssd1 vssd1 vccd1 vccd1 _06765_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__10659__A _10659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11254__S _11254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ _12285_/Q _13561_/A vssd1 vssd1 vccd1 vccd1 _09478_/A sky130_fd_sc_hd__xnor2_1
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06686_ _06686_/A _06692_/B _06692_/C vssd1 vssd1 vccd1 vccd1 _06687_/A sky130_fd_sc_hd__or3_1
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07033__A _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08425_ _08419_/X _08420_/X _08421_/X _08423_/X _08382_/X _08424_/X vssd1 vssd1 vccd1
+ vccd1 _08425_/X sky130_fd_sc_hd__mux4_1
X_13191__347 vssd1 vssd1 vccd1 vccd1 _13191__347/HI _13798_/A sky130_fd_sc_hd__conb_1
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08356_ _08358_/A _08358_/B _08360_/C vssd1 vssd1 vccd1 vccd1 _08357_/A sky130_fd_sc_hd__or3_1
XANTENNA__06872__A _06900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07307_ _07307_/A _07317_/B _07314_/C vssd1 vssd1 vccd1 vccd1 _07308_/A sky130_fd_sc_hd__or3_1
X_08287_ _08364_/C vssd1 vssd1 vccd1 vccd1 _08297_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__10394__A _11170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07238_ _07291_/A vssd1 vssd1 vccd1 vccd1 _07250_/B sky130_fd_sc_hd__clkbuf_1
X_13232__388 vssd1 vssd1 vccd1 vccd1 _13232__388/HI _13887_/A sky130_fd_sc_hd__conb_1
XFILLER_118_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11002__B _13948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07169_ _07180_/A _07177_/B _07173_/C vssd1 vssd1 vccd1 vccd1 _07170_/A sky130_fd_sc_hd__or3_1
XFILLER_133_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10180_ _13618_/A _12471_/Q _10180_/S vssd1 vssd1 vccd1 vccd1 _10181_/B sky130_fd_sc_hd__mux2_1
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13085__241 vssd1 vssd1 vccd1 vccd1 _13085__241/HI _13580_/A sky130_fd_sc_hd__conb_1
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13126__282 vssd1 vssd1 vccd1 vccd1 _13126__282/HI _13667_/A sky130_fd_sc_hd__conb_1
X_13870_ _13870_/A _06643_/X vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12821_ _12821_/CLK _12821_/D vssd1 vssd1 vccd1 vccd1 _12821_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10569__A _10988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ _12753_/CLK _12752_/D vssd1 vssd1 vccd1 vccd1 _13879_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11703_/A _11703_/B _11703_/C vssd1 vssd1 vccd1 vccd1 _11704_/A sky130_fd_sc_hd__and3_1
XFILLER_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12806_/CLK _12683_/D vssd1 vssd1 vccd1 vccd1 _13812_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11634_/A _11645_/C _11645_/D vssd1 vssd1 vccd1 vccd1 _11634_/X sky130_fd_sc_hd__and3_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11565_ _11626_/B _11625_/A _11565_/C vssd1 vssd1 vccd1 vccd1 _11565_/X sky130_fd_sc_hd__and3_1
XFILLER_11_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10516_ _13680_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _10516_/X sky130_fd_sc_hd__or2_1
XFILLER_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11496_ _13979_/Z _11499_/B vssd1 vssd1 vccd1 vccd1 _11496_/X sky130_fd_sc_hd__or2_1
XFILLER_143_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10447_ _13684_/A _12539_/Q _10456_/S vssd1 vssd1 vccd1 vccd1 _10448_/B sky130_fd_sc_hd__mux2_1
X_10378_ _11156_/B _12060_/A _10693_/C vssd1 vssd1 vccd1 vccd1 _10409_/A sky130_fd_sc_hd__or3_4
XFILLER_97_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12117_ _12134_/A vssd1 vssd1 vccd1 vccd1 _12132_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12048_ _12927_/Q _13366_/A vssd1 vssd1 vccd1 vccd1 _12050_/C sky130_fd_sc_hd__xor2_1
XFILLER_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10479__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13999_ _13999_/A _08190_/X vssd1 vssd1 vccd1 vccd1 _14063_/Z sky130_fd_sc_hd__ebufn_8
X_06540_ _06556_/A _06540_/B _06540_/C vssd1 vssd1 vccd1 vccd1 _06541_/A sky130_fd_sc_hd__or3_1
XFILLER_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06471_ _06471_/A vssd1 vssd1 vccd1 vccd1 _06471_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08210_ _08210_/A vssd1 vssd1 vccd1 vccd1 _08263_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_33_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09190_ _09092_/X _09152_/B _09189_/X _09141_/X vssd1 vssd1 vccd1 vccd1 _12226_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08141_ _08153_/A vssd1 vssd1 vccd1 vccd1 _08151_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_119_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ _08072_/A vssd1 vssd1 vccd1 vccd1 _08087_/C sky130_fd_sc_hd__clkbuf_1
X_07023_ _07031_/A _07031_/B vssd1 vssd1 vccd1 vccd1 _07024_/A sky130_fd_sc_hd__or2_1
XFILLER_127_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13069__225 vssd1 vssd1 vccd1 vccd1 _13069__225/HI _13544_/A sky130_fd_sc_hd__conb_1
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09508__A _09636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07954__C _07962_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08974_ _12828_/Q vssd1 vssd1 vccd1 vccd1 _11632_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10380__C _10693_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08131__B _08189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07925_ _07936_/A _07931_/B _07931_/C vssd1 vssd1 vccd1 vccd1 _07926_/A sky130_fd_sc_hd__or3_1
XFILLER_130_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07856_ _08084_/A vssd1 vssd1 vccd1 vccd1 _07962_/B sky130_fd_sc_hd__buf_4
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06807_ _06807_/A vssd1 vssd1 vccd1 vccd1 _06807_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07787_ _07796_/A _07792_/B _07787_/C vssd1 vssd1 vccd1 vccd1 _07788_/A sky130_fd_sc_hd__or3_1
XFILLER_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09526_ _10552_/A _09526_/B vssd1 vssd1 vccd1 vccd1 _09526_/X sky130_fd_sc_hd__or2_1
X_06738_ _06746_/A _06738_/B _06738_/C vssd1 vssd1 vccd1 vccd1 _06739_/A sky130_fd_sc_hd__or3_1
XFILLER_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _12284_/Q _13560_/A vssd1 vssd1 vccd1 vccd1 _09468_/A sky130_fd_sc_hd__xnor2_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06669_ _06673_/A _06678_/B _06678_/C vssd1 vssd1 vccd1 vccd1 _06670_/A sky130_fd_sc_hd__or3_1
XFILLER_24_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08408_ _12254_/Q vssd1 vssd1 vccd1 vccd1 _09320_/D sky130_fd_sc_hd__clkbuf_2
X_09388_ _12273_/Q _09388_/B _09388_/C vssd1 vssd1 vccd1 vccd1 _09391_/B sky130_fd_sc_hd__nand3_1
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08339_ _08347_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08340_/A sky130_fd_sc_hd__or2_1
XFILLER_165_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11350_ _13909_/A _12766_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _11351_/B sky130_fd_sc_hd__mux2_1
XFILLER_138_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10301_ _13648_/A _12502_/Q _10375_/B vssd1 vssd1 vccd1 vccd1 _10302_/B sky130_fd_sc_hd__mux2_1
X_11281_ _11408_/A _11281_/B _11281_/C vssd1 vssd1 vccd1 vccd1 _11282_/A sky130_fd_sc_hd__and3_1
XFILLER_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10232_ _10232_/A _10232_/B _10232_/C _10232_/D vssd1 vssd1 vccd1 vccd1 _10243_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_126_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10163_ _10163_/A _10163_/B _10163_/C _10163_/D vssd1 vssd1 vccd1 vccd1 _10166_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_160_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10094_ _10101_/B _10094_/B vssd1 vssd1 vccd1 vccd1 _10095_/C sky130_fd_sc_hd__nand2_1
XFILLER_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13922_ _13922_/A _06495_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
XFILLER_74_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13853_ _13853_/A _06687_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[14] sky130_fd_sc_hd__ebufn_8
XFILLER_62_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11248__A1 _12740_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12804_ _12853_/CLK _12804_/D vssd1 vssd1 vccd1 vccd1 _13978_/A sky130_fd_sc_hd__dfxtp_2
X_10996_ _13822_/A _12676_/Q _10996_/S vssd1 vssd1 vccd1 vccd1 _10997_/B sky130_fd_sc_hd__mux2_1
XFILLER_90_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13784_ _13784_/A _06881_/X vssd1 vssd1 vccd1 vccd1 _13976_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_15_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12753_/CLK _12735_/D vssd1 vssd1 vccd1 vccd1 _12735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13403__A _13403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ _12853_/CLK _12666_/D vssd1 vssd1 vccd1 vccd1 _12666_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09600__B _13566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07401__A _07822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11617_ _11630_/D _11616_/C _11641_/A vssd1 vssd1 vccd1 vccd1 _11618_/C sky130_fd_sc_hd__a21o_1
X_12597_ _12597_/CLK _12597_/D vssd1 vssd1 vccd1 vccd1 _13724_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11420__A1 _10645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11548_ _11576_/A vssd1 vssd1 vccd1 vccd1 _11604_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_156_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11479_ _09089_/S _11459_/X _11478_/X _11464_/X vssd1 vssd1 vccd1 vccd1 _12798_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10931__B1 _10757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _07714_/A _07710_/B _07719_/C vssd1 vssd1 vccd1 vccd1 _07711_/A sky130_fd_sc_hd__or3_1
XFILLER_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08690_ _10130_/A _12460_/Q _12461_/Q _12462_/Q _08602_/X _08603_/X vssd1 vssd1 vccd1
+ vccd1 _08690_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07641_ _07644_/A _07641_/B _07649_/C vssd1 vssd1 vccd1 vccd1 _07642_/A sky130_fd_sc_hd__or3_1
XFILLER_26_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09998__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07572_ _07739_/A _07995_/B _08089_/B vssd1 vssd1 vccd1 vccd1 _07573_/A sky130_fd_sc_hd__or3_1
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09311_ _09329_/A _09312_/B vssd1 vssd1 vccd1 vccd1 _09313_/B sky130_fd_sc_hd__or2_1
XANTENNA__09301__B1 _09236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06523_ _06523_/A vssd1 vssd1 vccd1 vccd1 _06534_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08655__A2 _08568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ _09317_/A _09317_/B _09242_/C vssd1 vssd1 vccd1 vccd1 _09253_/C sky130_fd_sc_hd__and3_1
X_06454_ _06454_/A vssd1 vssd1 vccd1 vccd1 _06454_/X sky130_fd_sc_hd__clkbuf_1
X_09173_ _09636_/A vssd1 vssd1 vccd1 vccd1 _10665_/A sky130_fd_sc_hd__buf_4
X_06385_ _06391_/A _08349_/A vssd1 vssd1 vccd1 vccd1 _06386_/A sky130_fd_sc_hd__or2_1
X_08124_ _08150_/A vssd1 vssd1 vccd1 vccd1 _08135_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08055_ _08065_/A _08110_/B _08057_/C vssd1 vssd1 vccd1 vccd1 _08056_/A sky130_fd_sc_hd__or3_1
XFILLER_162_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07006_ _07006_/A vssd1 vssd1 vccd1 vccd1 _07006_/X sky130_fd_sc_hd__clkbuf_1
Xoutput28 _13401_/A vssd1 vssd1 vccd1 vccd1 pwm_en[0] sky130_fd_sc_hd__buf_2
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput39 _13594_/A vssd1 vssd1 vccd1 vccd1 pwm_en[5] sky130_fd_sc_hd__buf_2
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07981__A _08064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _12828_/Q _11641_/D _12830_/Q _12831_/Q _08918_/X _08919_/X vssd1 vssd1 vccd1
+ vccd1 _08957_/X sky130_fd_sc_hd__mux4_2
XFILLER_57_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07908_ _07908_/A _07917_/B _07917_/C vssd1 vssd1 vccd1 vccd1 _07909_/A sky130_fd_sc_hd__or3_1
X_08888_ _10921_/C _12655_/Q _10921_/A _12657_/Q _10697_/A _08887_/X vssd1 vssd1 vccd1
+ vccd1 _08888_/X sky130_fd_sc_hd__mux4_2
XFILLER_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07839_ _08335_/A vssd1 vssd1 vccd1 vccd1 _07852_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10850_ _10854_/C _10850_/B vssd1 vssd1 vccd1 vccd1 _12639_/D sky130_fd_sc_hd__nor2_1
X_13197__353 vssd1 vssd1 vccd1 vccd1 _13197__353/HI _13804_/A sky130_fd_sc_hd__conb_1
XFILLER_71_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09509_ _09634_/A vssd1 vssd1 vccd1 vccd1 _09509_/X sky130_fd_sc_hd__clkbuf_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _10820_/C vssd1 vssd1 vccd1 vccd1 _10781_/X sky130_fd_sc_hd__buf_2
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12520_ _12522_/CLK _12520_/D vssd1 vssd1 vccd1 vccd1 _13649_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11650__A1 _11689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13238__394 vssd1 vssd1 vccd1 vccd1 _13238__394/HI _13893_/A sky130_fd_sc_hd__conb_1
XANTENNA__08317__A _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12451_ _12451_/CLK _12451_/D vssd1 vssd1 vccd1 vccd1 _12451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11402_ _12760_/Q _13935_/A vssd1 vssd1 vccd1 vccd1 _11405_/B sky130_fd_sc_hd__xor2_1
XFILLER_165_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12382_ _12386_/CLK _12382_/D vssd1 vssd1 vccd1 vccd1 _12382_/Q sky130_fd_sc_hd__dfxtp_1
X_14121_ _14121_/A _08265_/X vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__ebufn_8
X_11333_ _13904_/A _12761_/Q _11408_/B vssd1 vssd1 vccd1 vccd1 _11334_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09148__A _11490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ _14052_/A _07918_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[21] sky130_fd_sc_hd__ebufn_8
X_11264_ _12737_/Q _13945_/A vssd1 vssd1 vccd1 vccd1 _11268_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11397__B _13950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10215_ _10298_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__and2_1
X_11195_ _11195_/A vssd1 vssd1 vccd1 vccd1 _11195_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09582__S _09582_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ _10146_/A _10146_/B _10146_/C vssd1 vssd1 vccd1 vccd1 _10147_/A sky130_fd_sc_hd__and3_1
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10077_ _10077_/A vssd1 vssd1 vccd1 vccd1 _10135_/B sky130_fd_sc_hd__clkbuf_2
X_13905_ _13905_/A _06541_/X vssd1 vssd1 vccd1 vccd1 _14065_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13836_ _13836_/A _06734_/X vssd1 vssd1 vccd1 vccd1 _14028_/Z sky130_fd_sc_hd__ebufn_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10979_ _13817_/A _12671_/Q _10990_/S vssd1 vssd1 vccd1 vccd1 _10980_/B sky130_fd_sc_hd__mux2_1
X_13767_ _13767_/A _06924_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12718_ _12722_/CLK _12718_/D vssd1 vssd1 vccd1 vccd1 _13846_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08227__A _08240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13698_ _13698_/A _07098_/X vssd1 vssd1 vccd1 vccd1 _14082_/Z sky130_fd_sc_hd__ebufn_8
X_12649_ _12652_/CLK _12649_/D vssd1 vssd1 vccd1 vccd1 _12649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09984__C _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13031__187 vssd1 vssd1 vccd1 vccd1 _13031__187/HI _13474_/A sky130_fd_sc_hd__conb_1
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09860_ _12386_/Q _13563_/A vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__xor2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _13779_/A vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__buf_2
X_09791_ _13593_/A _09791_/B vssd1 vssd1 vccd1 vccd1 _09843_/S sky130_fd_sc_hd__and2_2
XFILLER_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater100 _14086_/Z vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__buf_12
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater111 _14082_/Z vssd1 vssd1 vccd1 vccd1 _13666_/Z sky130_fd_sc_hd__buf_12
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08742_ _13776_/A vssd1 vssd1 vccd1 vccd1 _08742_/X sky130_fd_sc_hd__clkbuf_4
Xrepeater122 peripheralBus_data[14] vssd1 vssd1 vccd1 vccd1 _14077_/Z sky130_fd_sc_hd__buf_12
Xrepeater133 _13625_/Z vssd1 vssd1 vccd1 vccd1 _14105_/Z sky130_fd_sc_hd__buf_12
XFILLER_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08673_ _12459_/Q vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08420__S1 _08374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07624_ _07630_/A _07626_/B _07635_/C vssd1 vssd1 vccd1 vccd1 _07625_/A sky130_fd_sc_hd__or3_1
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09521__A _11064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07555_ _07555_/A vssd1 vssd1 vccd1 vccd1 _07555_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10667__A _10667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06506_ _06506_/A vssd1 vssd1 vccd1 vccd1 _06506_/X sky130_fd_sc_hd__clkbuf_1
X_07486_ _08089_/A _08089_/B vssd1 vssd1 vccd1 vccd1 _07487_/A sky130_fd_sc_hd__or2_1
XFILLER_22_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09225_ _09316_/D _09223_/A _09217_/X vssd1 vssd1 vccd1 vccd1 _09226_/B sky130_fd_sc_hd__o21ai_1
X_06437_ _06440_/A _06437_/B vssd1 vssd1 vccd1 vccd1 _06438_/A sky130_fd_sc_hd__or2_1
XANTENNA__13978__A _13978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09156_ _09156_/A vssd1 vssd1 vccd1 vccd1 _09179_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06368_ _06368_/A vssd1 vssd1 vccd1 vccd1 _06368_/X sky130_fd_sc_hd__clkbuf_1
X_08107_ _08153_/A vssd1 vssd1 vccd1 vccd1 _08122_/C sky130_fd_sc_hd__clkbuf_1
X_09087_ _11695_/B _12851_/Q _12852_/Q _12853_/Q _09067_/X _09068_/X vssd1 vssd1 vccd1
+ vccd1 _09087_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_110_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _12313_/CLK sky130_fd_sc_hd__clkbuf_16
X_06299_ _06303_/A _06308_/B _06308_/C vssd1 vssd1 vccd1 vccd1 _06300_/A sky130_fd_sc_hd__or3_1
XFILLER_123_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08038_ _08038_/A vssd1 vssd1 vccd1 vccd1 _08038_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11010__B _13938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10000_ _10008_/D _10000_/B vssd1 vssd1 vccd1 vccd1 _12428_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08600__A _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ _09993_/C _09989_/B vssd1 vssd1 vccd1 vccd1 _12425_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11951_ _09633_/A _14038_/A _11957_/S vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__mux2_1
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10902_ _10907_/B _10903_/B vssd1 vssd1 vccd1 vccd1 _10904_/B sky130_fd_sc_hd__or2_1
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11882_ _12897_/Q _14041_/A _11895_/S vssd1 vssd1 vccd1 vccd1 _11883_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13621_ _13621_/A _07304_/X vssd1 vssd1 vccd1 vccd1 _13973_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10833_ _10833_/A _10877_/A vssd1 vssd1 vccd1 vccd1 _10833_/X sky130_fd_sc_hd__and2_1
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10426__A2 _10409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13552_ _13552_/A _07487_/X vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10764_ _10773_/B vssd1 vssd1 vccd1 vccd1 _10864_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12503_ _12515_/CLK _12503_/D vssd1 vssd1 vccd1 vccd1 _12503_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater69 peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 _13973_/Z sky130_fd_sc_hd__buf_12
X_13483_ _13483_/A _07665_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
X_10695_ _10872_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10695_/X sky130_fd_sc_hd__or2_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12434_ _12617_/CLK _12434_/D vssd1 vssd1 vccd1 vccd1 _12434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12365_ _12369_/CLK _12365_/D vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_101_clk _12555_/CLK vssd1 vssd1 vccd1 vccd1 _12420_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11201__A _13978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11316_ _13882_/A _11323_/B vssd1 vssd1 vccd1 vccd1 _11316_/X sky130_fd_sc_hd__or2_1
X_14104_ _14104_/A _08221_/X vssd1 vssd1 vccd1 vccd1 _14104_/Z sky130_fd_sc_hd__ebufn_8
X_12296_ _12301_/CLK _12296_/D vssd1 vssd1 vccd1 vccd1 _13427_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_153_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14035_ _14035_/A _07874_/X vssd1 vssd1 vccd1 vccd1 _14035_/Z sky130_fd_sc_hd__ebufn_8
X_11247_ _11247_/A vssd1 vssd1 vccd1 vccd1 _12739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11178_ _10662_/X _11171_/X _11177_/X _11166_/X vssd1 vssd1 vccd1 vccd1 _12718_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10129_ _10130_/A vssd1 vssd1 vccd1 vccd1 _10129_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12032__A _12134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13819_ _13819_/A _06781_/X vssd1 vssd1 vccd1 vccd1 _13979_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07340_ _07342_/A _07351_/B _07347_/C vssd1 vssd1 vccd1 vccd1 _07341_/A sky130_fd_sc_hd__or3_1
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07271_ _07279_/A _07276_/B _07273_/C vssd1 vssd1 vccd1 vccd1 _07272_/A sky130_fd_sc_hd__or3_1
XFILLER_148_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09010_ _08997_/X _09009_/X _09071_/S vssd1 vssd1 vccd1 vccd1 _10939_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10050__B1 _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09991__B1 _09987_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09912_ _09112_/X _09902_/X _09911_/X _09905_/X vssd1 vssd1 vccd1 vccd1 _12404_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater90_A _13995_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _13534_/A _12389_/Q _09843_/S vssd1 vssd1 vccd1 vccd1 _09844_/B sky130_fd_sc_hd__mux2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07962__C _07962_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _07979_/B vssd1 vssd1 vccd1 vccd1 _06995_/B sky130_fd_sc_hd__clkbuf_1
X_09774_ _13496_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09774_/X sky130_fd_sc_hd__or2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08725_ _12465_/Q vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _08653_/X _08655_/X _13588_/A vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__mux2_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_54_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _07607_/A vssd1 vssd1 vccd1 vccd1 _07607_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _12440_/Q vssd1 vssd1 vccd1 vccd1 _10052_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ _07545_/A _07545_/B _07538_/C vssd1 vssd1 vccd1 vccd1 _07539_/A sky130_fd_sc_hd__or3_1
XFILLER_50_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11005__B _13946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ _07478_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07470_/A sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_69_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ _09210_/B _09201_/X _09207_/Y vssd1 vssd1 vccd1 vccd1 _12230_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__13501__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10480_ _13694_/A _12549_/Q _10480_/S vssd1 vssd1 vccd1 vccd1 _10481_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_112_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ _11160_/A vssd1 vssd1 vccd1 vccd1 _09139_/X sky130_fd_sc_hd__buf_4
XANTENNA__12117__A _12134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12150_ _12150_/A vssd1 vssd1 vccd1 vccd1 _12966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11101_ _13847_/A _12702_/Q _11101_/S vssd1 vssd1 vccd1 vccd1 _11102_/B sky130_fd_sc_hd__mux2_1
XFILLER_135_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12081_ _14070_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12081_/X sky130_fd_sc_hd__or2_1
XANTENNA__10860__A _10936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ _13808_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11032_/X sky130_fd_sc_hd__or2_1
XFILLER_1_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11541__B1 _11540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11934_ _09620_/A _14033_/A _11940_/S vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__mux2_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11865_ _12892_/Q _14036_/A _11878_/S vssd1 vssd1 vccd1 vccd1 _11866_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13604_ _13604_/A _07355_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10816_ _10870_/D _10878_/B _10815_/Y vssd1 vssd1 vccd1 vccd1 _12630_/D sky130_fd_sc_hd__a21oi_1
X_11796_ _11799_/A _11796_/B vssd1 vssd1 vccd1 vccd1 _11797_/A sky130_fd_sc_hd__and2_1
XANTENNA__08699__S1 _08603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13535_ _13535_/A _07530_/X vssd1 vssd1 vccd1 vccd1 _14111_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10747_ _13775_/A _10806_/B _10806_/C _10806_/D vssd1 vssd1 vccd1 vccd1 _10760_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13466_ _13466_/A _07711_/X vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_8
X_10678_ _10414_/X _10673_/X _10677_/X _10668_/X vssd1 vssd1 vccd1 vccd1 _12595_/D
+ sky130_fd_sc_hd__o211a_1
X_12417_ _12418_/CLK _12417_/D vssd1 vssd1 vccd1 vccd1 _13593_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_64_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13397_ _13397_/A _08363_/X vssd1 vssd1 vccd1 vccd1 _14037_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12348_ _12349_/CLK _12348_/D vssd1 vssd1 vccd1 vccd1 _12348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12279_ _12289_/CLK _12279_/D vssd1 vssd1 vccd1 vccd1 _12279_/Q sky130_fd_sc_hd__dfxtp_1
X_14018_ _14018_/A _08117_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08240__A _08240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ _06840_/A vssd1 vssd1 vccd1 vccd1 _06840_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06771_ _06775_/A _06780_/B _06780_/C vssd1 vssd1 vccd1 vccd1 _06772_/A sky130_fd_sc_hd__or3_1
XANTENNA__09489__C1 _09192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08510_ _11707_/C vssd1 vssd1 vccd1 vccd1 _13369_/A sky130_fd_sc_hd__buf_4
XFILLER_76_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13143__299 vssd1 vssd1 vccd1 vccd1 _13143__299/HI _13700_/A sky130_fd_sc_hd__conb_1
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09490_ _09620_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _09490_/X sky130_fd_sc_hd__or2_1
XFILLER_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08441_ _12241_/Q vssd1 vssd1 vccd1 vccd1 _09315_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08372_ _12235_/Q vssd1 vssd1 vccd1 vccd1 _09316_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07323_ _07827_/A _07323_/B _08089_/B vssd1 vssd1 vccd1 vccd1 _07324_/A sky130_fd_sc_hd__or3_1
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07254_ _07254_/A vssd1 vssd1 vccd1 vccd1 _07254_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08415__A _11706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13037__193 vssd1 vssd1 vccd1 vccd1 _13037__193/HI _13480_/A sky130_fd_sc_hd__conb_1
X_07185_ _07193_/A _07190_/B _07187_/C vssd1 vssd1 vccd1 vccd1 _07186_/A sky130_fd_sc_hd__or3_1
XFILLER_117_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09826_ _09826_/A vssd1 vssd1 vccd1 vccd1 _12383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09757_ _13491_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09757_/X sky130_fd_sc_hd__or2_1
XFILLER_27_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06969_ _06969_/A vssd1 vssd1 vccd1 vccd1 _06969_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _08708_/A vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__buf_2
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09967_/B vssd1 vssd1 vccd1 vccd1 _10988_/A sky130_fd_sc_hd__buf_6
XFILLER_104_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _12445_/Q vssd1 vssd1 vccd1 vccd1 _10098_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11689_/A _11688_/B _11657_/C vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__a21oi_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ _13724_/A _12580_/Q _10601_/S vssd1 vssd1 vccd1 vccd1 _10602_/B sky130_fd_sc_hd__mux2_1
X_11581_ _11634_/A _11632_/D _11649_/C _11639_/B vssd1 vssd1 vccd1 vccd1 _11582_/B
+ sky130_fd_sc_hd__a31o_1
X_10532_ _09767_/X _10525_/X _10531_/X _10523_/X vssd1 vssd1 vccd1 vccd1 _12558_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10463_ _10479_/A vssd1 vssd1 vccd1 vccd1 _10477_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_108_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12202_ _14103_/A _12206_/B vssd1 vssd1 vccd1 vccd1 _12202_/X sky130_fd_sc_hd__or2_1
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10394_ _11170_/A vssd1 vssd1 vccd1 vccd1 _10394_/X sky130_fd_sc_hd__buf_6
XFILLER_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12133_ _12133_/A vssd1 vssd1 vccd1 vccd1 _12961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12064_ _14063_/A _12073_/B vssd1 vssd1 vccd1 vccd1 _12064_/X sky130_fd_sc_hd__or2_1
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11015_ _12663_/Q _13937_/A vssd1 vssd1 vccd1 vccd1 _11016_/D sky130_fd_sc_hd__xor2_1
XFILLER_38_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09603__B _13551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ _12968_/CLK _12966_/D vssd1 vssd1 vccd1 vccd1 _12966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07404__A _07822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11917_ _12895_/Q _13367_/A vssd1 vssd1 vccd1 vccd1 _11920_/B sky130_fd_sc_hd__xor2_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12914_/CLK _12897_/D vssd1 vssd1 vccd1 vccd1 _12897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11848_ _12887_/Q _14031_/A _11861_/S vssd1 vssd1 vccd1 vccd1 _11849_/B sky130_fd_sc_hd__mux2_1
XFILLER_159_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11779_ _12866_/Q _13371_/A vssd1 vssd1 vccd1 vccd1 _11780_/D sky130_fd_sc_hd__xor2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13518_ _13518_/A _07573_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10484__B _13754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13449_ _13449_/A _07754_/X vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_161_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08990_ _12821_/Q vssd1 vssd1 vccd1 vccd1 _11626_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07941_ _07951_/A _07945_/B _07945_/C vssd1 vssd1 vccd1 vccd1 _07942_/A sky130_fd_sc_hd__or3_1
XFILLER_130_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12759__CLK _12759_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _07872_/A vssd1 vssd1 vccd1 vccd1 _07872_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09611_ _09611_/A vssd1 vssd1 vccd1 vccd1 _12324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06823_ _06823_/A vssd1 vssd1 vccd1 vccd1 _06823_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09542_ _09546_/A _09542_/B vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__and2_1
X_06754_ _11028_/B vssd1 vssd1 vccd1 vccd1 _06809_/A sky130_fd_sc_hd__buf_2
XFILLER_64_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09473_ _09473_/A _09473_/B _09473_/C _09473_/D vssd1 vssd1 vccd1 vccd1 _09479_/B
+ sky130_fd_sc_hd__and4_1
X_06685_ _06685_/A vssd1 vssd1 vccd1 vccd1 _06685_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_90_clk _12438_/CLK vssd1 vssd1 vccd1 vccd1 _12467_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10378__C _10693_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ _13395_/A vssd1 vssd1 vccd1 vccd1 _08424_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08355_ _08355_/A vssd1 vssd1 vccd1 vccd1 _08355_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08532__S0 _09140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07317_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_149_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08286_ _08286_/A vssd1 vssd1 vccd1 vccd1 _08286_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07237_ _09484_/A vssd1 vssd1 vccd1 vccd1 _07291_/A sky130_fd_sc_hd__buf_2
XFILLER_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07168_ _07208_/A vssd1 vssd1 vccd1 vccd1 _07180_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10547__A1 _10288_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07099_ _07108_/A _07105_/B _07101_/C vssd1 vssd1 vccd1 vccd1 _07100_/A sky130_fd_sc_hd__or3_1
XFILLER_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09809_ _09809_/A vssd1 vssd1 vccd1 vccd1 _12378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12820_ _12820_/CLK _12820_/D vssd1 vssd1 vccd1 vccd1 _12820_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12751_ _12753_/CLK _12751_/D vssd1 vssd1 vccd1 vccd1 _13878_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _12660_/CLK sky130_fd_sc_hd__clkbuf_16
X_11702_ _12853_/Q _11702_/B vssd1 vssd1 vccd1 vccd1 _11703_/C sky130_fd_sc_hd__nand2_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12682_/CLK _12682_/D vssd1 vssd1 vccd1 vccd1 _13811_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11633_ _11633_/A _11633_/B _11633_/C _11633_/D vssd1 vssd1 vccd1 vccd1 _11645_/D
+ sky130_fd_sc_hd__and4_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11564_ _11625_/A _11565_/C _11563_/Y _11515_/X vssd1 vssd1 vccd1 vccd1 _12820_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10515_ _10377_/X _10511_/X _10514_/X _10425_/X vssd1 vssd1 vccd1 vccd1 _12551_/D
+ sky130_fd_sc_hd__o211a_1
X_11495_ _13978_/A _11459_/X _11494_/X _11464_/X vssd1 vssd1 vccd1 vccd1 _12804_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10446_ _10479_/A vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10377_ _11153_/A vssd1 vssd1 vccd1 vccd1 _10377_/X sky130_fd_sc_hd__buf_6
XANTENNA_repeater121_A peripheralBus_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12116_ _12116_/A vssd1 vssd1 vccd1 vccd1 _12956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12047_ _12935_/Q _13374_/A vssd1 vssd1 vccd1 vccd1 _12050_/B sky130_fd_sc_hd__xor2_1
XFILLER_49_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output50_A _13954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11582__C _11582_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13998_ _13998_/A _06287_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07134__A _07615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ _12952_/CLK _12949_/D vssd1 vssd1 vccd1 vccd1 _14075_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_72_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _12550_/CLK sky130_fd_sc_hd__clkbuf_16
X_06470_ _06481_/A _07827_/B _06472_/C vssd1 vssd1 vccd1 vccd1 _06471_/A sky130_fd_sc_hd__or3_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08140_ _11283_/B vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_147_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11974__A0 _14109_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08071_ _08071_/A vssd1 vssd1 vccd1 vccd1 _08071_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07022_ _10637_/A vssd1 vssd1 vccd1 vccd1 _07031_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_161_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08973_ _08966_/X _08969_/X _08970_/X _08972_/X _08924_/X _08925_/X vssd1 vssd1 vccd1
+ vccd1 _08973_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08131__C _08131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07924_ _07999_/A vssd1 vssd1 vccd1 vccd1 _07936_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09524__A _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__B _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ _07855_/A vssd1 vssd1 vccd1 vccd1 _07855_/X sky130_fd_sc_hd__clkbuf_1
X_06806_ _07857_/A _06806_/B _06806_/C vssd1 vssd1 vccd1 vccd1 _06807_/A sky130_fd_sc_hd__or3_1
XFILLER_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07786_ _07786_/A vssd1 vssd1 vccd1 vccd1 _07786_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ _13437_/A _09513_/X _09524_/X _09522_/X vssd1 vssd1 vccd1 vccd1 _12306_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06737_ _06737_/A vssd1 vssd1 vccd1 vccd1 _06737_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_63_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _12813_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09456_/A vssd1 vssd1 vccd1 vccd1 _12290_/D sky130_fd_sc_hd__clkbuf_1
X_06668_ _06722_/A vssd1 vssd1 vccd1 vccd1 _06678_/C sky130_fd_sc_hd__clkbuf_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08407_ _12249_/Q _12250_/Q _12251_/Q _12252_/Q _08379_/X _08380_/X vssd1 vssd1 vccd1
+ vccd1 _08407_/X sky130_fd_sc_hd__mux4_2
XFILLER_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09387_ _09388_/B _09388_/C _12273_/Q vssd1 vssd1 vccd1 vccd1 _09389_/B sky130_fd_sc_hd__a21o_1
X_06599_ _06599_/A vssd1 vssd1 vccd1 vccd1 _06610_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08338_ _08338_/A vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__08425__A3 _08423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__A0 _14106_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11013__B _13950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13349__505 vssd1 vssd1 vccd1 vccd1 _13349__505/HI _14118_/A sky130_fd_sc_hd__conb_1
X_08269_ _08269_/A vssd1 vssd1 vccd1 vccd1 _08269_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ _10317_/A vssd1 vssd1 vccd1 vccd1 _10315_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11280_ _11257_/Y _11263_/X _11279_/Y _13952_/A vssd1 vssd1 vccd1 vccd1 _11281_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10231_ _12482_/Q _13757_/A vssd1 vssd1 vccd1 vccd1 _10232_/D sky130_fd_sc_hd__xor2_1
XANTENNA__11193__A1 _11061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10162_ _10162_/A _10162_/B _10162_/C _10162_/D vssd1 vssd1 vccd1 vccd1 _10166_/A
+ sky130_fd_sc_hd__or4_1
XANTENNA__11964__A _11998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10093_ _10101_/B _10094_/B vssd1 vssd1 vccd1 vccd1 _10095_/B sky130_fd_sc_hd__or2_1
XANTENNA__09434__A _09454_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ _13921_/A _06498_/X vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13852_ _13852_/A _06691_/X vssd1 vssd1 vccd1 vccd1 _14012_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ _12806_/CLK _12803_/D vssd1 vssd1 vccd1 vccd1 _13977_/A sky130_fd_sc_hd__dfxtp_2
X_13783_ _13783_/A _06883_/X vssd1 vssd1 vccd1 vccd1 _14103_/Z sky130_fd_sc_hd__ebufn_8
X_10995_ _10995_/A vssd1 vssd1 vccd1 vccd1 _12675_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_54_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _12806_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _12753_/CLK _12734_/D vssd1 vssd1 vccd1 vccd1 _12734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12853_/CLK _12665_/D vssd1 vssd1 vccd1 vccd1 _12665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11616_ _11641_/A _11630_/D _11616_/C vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__and3_1
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12596_ _12597_/CLK _12596_/D vssd1 vssd1 vccd1 vccd1 _13723_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11547_ _11627_/B _11627_/C _11627_/D _11547_/D vssd1 vssd1 vccd1 vccd1 _11558_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_129_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11478_ _14068_/Z _11494_/B vssd1 vssd1 vccd1 vccd1 _11478_/X sky130_fd_sc_hd__or2_1
X_10429_ _10480_/S vssd1 vssd1 vccd1 vccd1 _10507_/B sky130_fd_sc_hd__clkbuf_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07640_ _07640_/A vssd1 vssd1 vccd1 vccd1 _07640_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07571_ _07571_/A vssd1 vssd1 vccd1 vccd1 _07571_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _12598_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09310_ _12256_/Q vssd1 vssd1 vccd1 vccd1 _09329_/A sky130_fd_sc_hd__clkbuf_1
X_06522_ _06522_/A vssd1 vssd1 vccd1 vccd1 _06522_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11644__C1 _11515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09241_ _09317_/B _09242_/C _09240_/Y vssd1 vssd1 vccd1 vccd1 _12238_/D sky130_fd_sc_hd__a21oi_1
X_06453_ _07845_/A _07845_/B vssd1 vssd1 vccd1 vccd1 _06454_/A sky130_fd_sc_hd__or2_1
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11114__A _11206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09172_ _14007_/Z vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__buf_4
X_06384_ _06384_/A vssd1 vssd1 vccd1 vccd1 _06384_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _08123_/A vssd1 vssd1 vccd1 vccd1 _08123_/X sky130_fd_sc_hd__clkbuf_1
X_08054_ _08067_/A vssd1 vssd1 vccd1 vccd1 _08065_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__09519__A _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11768__B _13372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07005_ _07007_/A _07007_/B vssd1 vssd1 vccd1 vccd1 _07006_/A sky130_fd_sc_hd__or2_1
Xoutput29 _13787_/A vssd1 vssd1 vccd1 vccd1 pwm_en[10] sky130_fd_sc_hd__buf_2
XFILLER_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08956_ _12829_/Q vssd1 vssd1 vccd1 vccd1 _11641_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07907_ _07920_/A vssd1 vssd1 vccd1 vccd1 _07917_/C sky130_fd_sc_hd__clkbuf_1
X_08887_ _08887_/A vssd1 vssd1 vccd1 vccd1 _08887_/X sky130_fd_sc_hd__buf_2
XFILLER_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07838_ _07838_/A vssd1 vssd1 vccd1 vccd1 _07838_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11008__B _13949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ _07769_/A _07779_/B _07774_/C vssd1 vssd1 vccd1 vccd1 _07770_/A sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_36_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _12704_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09508_ _09636_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09508_/X sky130_fd_sc_hd__or2_1
XANTENNA__08726__S0 _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ _10865_/C _10780_/B vssd1 vssd1 vccd1 vccd1 _10790_/C sky130_fd_sc_hd__and2_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09439_ _09439_/A _09439_/B vssd1 vssd1 vccd1 vccd1 _09440_/A sky130_fd_sc_hd__and2_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11024__A _11039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12450_ _12457_/CLK _12450_/D vssd1 vssd1 vccd1 vccd1 _12450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11401_ _12765_/Q _13940_/A vssd1 vssd1 vccd1 vccd1 _11405_/A sky130_fd_sc_hd__xor2_1
X_12381_ _12386_/CLK _12381_/D vssd1 vssd1 vccd1 vccd1 _12381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14120_ _14120_/A _08262_/X vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__ebufn_8
X_11332_ _11332_/A vssd1 vssd1 vccd1 vccd1 _12760_/D sky130_fd_sc_hd__clkbuf_1
X_14051_ _14051_/A _07916_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[20] sky130_fd_sc_hd__ebufn_8
X_11263_ _11258_/Y _11259_/X _11260_/Y _11261_/X _11262_/Y vssd1 vssd1 vccd1 vccd1
+ _11263_/X sky130_fd_sc_hd__o221a_1
XFILLER_141_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08052__B _08110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ _13628_/A _12481_/Q _10214_/S vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__mux2_1
X_11194_ _13852_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11194_/X sky130_fd_sc_hd__or2_1
XFILLER_79_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10145_ _10148_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _10146_/C sky130_fd_sc_hd__nand2_1
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09164__A peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ _10099_/A _10099_/B _10086_/B _10076_/D vssd1 vssd1 vccd1 vccd1 _10083_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13904_ _13904_/A _06546_/X vssd1 vssd1 vccd1 vccd1 _14064_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_63_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13835_ _13835_/A _06737_/X vssd1 vssd1 vccd1 vccd1 _13995_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ _13766_/A _06928_/X vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_8
X_10978_ _10978_/A vssd1 vssd1 vccd1 vccd1 _12670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07412__A _08131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12717_ _12722_/CLK _12717_/D vssd1 vssd1 vccd1 vccd1 _13845_/A sky130_fd_sc_hd__dfxtp_1
X_13697_ _13697_/A _07100_/X vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _12652_/CLK _12648_/D vssd1 vssd1 vccd1 vccd1 _12648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12579_ _12597_/CLK _12579_/D vssd1 vssd1 vccd1 vccd1 _12579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10492__B _13746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _13778_/A vssd1 vssd1 vccd1 vccd1 _08810_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_140_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09120_/X _09776_/A _09789_/X _09781_/X vssd1 vssd1 vccd1 vccd1 _12373_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater101 peripheralBus_data[23] vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__buf_12
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater112 peripheralBus_data[19] vssd1 vssd1 vccd1 vccd1 _14082_/Z sky130_fd_sc_hd__buf_12
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater123 peripheralBus_data[14] vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__buf_12
X_08741_ _10773_/D _12619_/Q _10773_/B _12621_/Q _08739_/X _08740_/X vssd1 vssd1 vccd1
+ vccd1 _08741_/X sky130_fd_sc_hd__mux4_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater134 peripheralBus_data[10] vssd1 vssd1 vccd1 vccd1 _13625_/Z sky130_fd_sc_hd__buf_12
XFILLER_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08672_ _12458_/Q vssd1 vssd1 vccd1 vccd1 _10130_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09802__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07623_ _07623_/A vssd1 vssd1 vccd1 vccd1 _07635_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_18_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _12946_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07554_ _07558_/A _07558_/B _07564_/C vssd1 vssd1 vccd1 vccd1 _07555_/A sky130_fd_sc_hd__or3_1
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06505_ _06507_/A _06512_/B _06512_/C vssd1 vssd1 vccd1 vccd1 _06506_/A sky130_fd_sc_hd__or3_1
X_07485_ _07485_/A vssd1 vssd1 vccd1 vccd1 _07485_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13270__426 vssd1 vssd1 vccd1 vccd1 _13270__426/HI _13961_/A sky130_fd_sc_hd__conb_1
XFILLER_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09224_ _09316_/D _09315_/C _09224_/C vssd1 vssd1 vccd1 vccd1 _09226_/A sky130_fd_sc_hd__and3_1
X_06436_ _06436_/A vssd1 vssd1 vccd1 vccd1 _06436_/X sky130_fd_sc_hd__clkbuf_1
X_09155_ _09625_/A vssd1 vssd1 vccd1 vccd1 _10652_/A sky130_fd_sc_hd__buf_4
X_06367_ _06822_/A _07822_/B _07822_/C vssd1 vssd1 vccd1 vccd1 _06368_/A sky130_fd_sc_hd__or3_1
XFILLER_108_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13311__467 vssd1 vssd1 vccd1 vccd1 _13311__467/HI _14048_/A sky130_fd_sc_hd__conb_1
X_08106_ _08106_/A vssd1 vssd1 vccd1 vccd1 _08106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09086_ _08993_/X _09002_/X _08999_/X _09004_/X _08934_/X _09030_/X vssd1 vssd1 vccd1
+ vccd1 _09086_/X sky130_fd_sc_hd__mux4_1
X_06298_ _06298_/A vssd1 vssd1 vccd1 vccd1 _06298_/X sky130_fd_sc_hd__clkbuf_1
X_08037_ _08039_/A _08047_/B _08044_/C vssd1 vssd1 vccd1 vccd1 _08038_/A sky130_fd_sc_hd__or3_1
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164__320 vssd1 vssd1 vccd1 vccd1 _13164__320/HI _13737_/A sky130_fd_sc_hd__conb_1
XFILLER_89_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09988_ _09997_/D _09982_/X _09987_/X vssd1 vssd1 vccd1 vccd1 _09989_/B sky130_fd_sc_hd__o21ai_1
XFILLER_89_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08939_ _12809_/Q vssd1 vssd1 vccd1 vccd1 _11518_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13205__361 vssd1 vssd1 vccd1 vccd1 _13205__361/HI _13828_/A sky130_fd_sc_hd__conb_1
X_11950_ _11950_/A vssd1 vssd1 vccd1 vccd1 _12910_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11320__A1 _11061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08867__A3 _08866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ _10901_/A _10903_/B vssd1 vssd1 vccd1 vccd1 _12650_/D sky130_fd_sc_hd__nor2_1
XFILLER_84_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11881_ _11898_/S vssd1 vssd1 vccd1 vccd1 _11895_/S sky130_fd_sc_hd__buf_2
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13620_ _13620_/A _07308_/X vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_8
X_10832_ _10870_/A _10870_/B _10869_/C _10869_/D vssd1 vssd1 vccd1 vccd1 _10877_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_25_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13551_ _13551_/A _08090_/X vssd1 vssd1 vccd1 vccd1 _13775_/Z sky130_fd_sc_hd__ebufn_8
X_10763_ _10763_/A vssd1 vssd1 vccd1 vccd1 _12619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12502_ _12505_/CLK _12502_/D vssd1 vssd1 vccd1 vccd1 _12502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13482_ _13482_/A _07668_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_139_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10694_ _10732_/B vssd1 vssd1 vccd1 vccd1 _10728_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11689__A _11689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ _12617_/CLK _12433_/D vssd1 vssd1 vccd1 vccd1 _12433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09159__A _14100_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ _12367_/CLK _12364_/D vssd1 vssd1 vccd1 vccd1 _13493_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14103_ _14103_/A _08219_/X vssd1 vssd1 vccd1 vccd1 _14103_/Z sky130_fd_sc_hd__ebufn_8
X_11315_ _11184_/X _11312_/X _11314_/X _11306_/X vssd1 vssd1 vccd1 vccd1 _12754_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12295_ _12295_/CLK _12295_/D vssd1 vssd1 vccd1 vccd1 _13426_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_153_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14034_ _14034_/A _07872_/X vssd1 vssd1 vccd1 vccd1 _14034_/Z sky130_fd_sc_hd__ebufn_8
X_11246_ _11255_/A _11246_/B vssd1 vssd1 vccd1 vccd1 _11247_/A sky130_fd_sc_hd__and2_1
XFILLER_106_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09752__A1 _09750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ _13846_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11177_/X sky130_fd_sc_hd__or2_1
XANTENNA__09606__B _13555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07407__A _08084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ _10128_/A vssd1 vssd1 vccd1 vccd1 _12458_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__06311__A _06688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10059_ _10088_/C _10060_/C _10058_/Y vssd1 vssd1 vccd1 vccd1 _12443_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__11311__A1 _10670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13818_ _13818_/A _06785_/X vssd1 vssd1 vccd1 vccd1 _13978_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10487__B _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ _13749_/A _06969_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[6] sky130_fd_sc_hd__ebufn_8
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07270_ _07270_/A vssd1 vssd1 vccd1 vccd1 _07270_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06981__A _08266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13148__304 vssd1 vssd1 vccd1 vccd1 _13148__304/HI _13705_/A sky130_fd_sc_hd__conb_1
X_09911_ _13532_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09911_/X sky130_fd_sc_hd__or2_1
XFILLER_144_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09842_ _09842_/A vssd1 vssd1 vccd1 vccd1 _12388_/D sky130_fd_sc_hd__clkbuf_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater83_A _14125_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _10670_/A vssd1 vssd1 vccd1 vccd1 _09773_/X sky130_fd_sc_hd__buf_6
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _10637_/A vssd1 vssd1 vccd1 vccd1 _07979_/B sky130_fd_sc_hd__clkbuf_4
X_08724_ _08631_/X _08640_/X _08637_/X _08643_/X _08563_/X _08670_/X vssd1 vssd1 vccd1
+ vccd1 _08724_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11302__A1 _11170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11781__B _13364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _08566_/X _08567_/X _08568_/X _08654_/X _08670_/A _08563_/X vssd1 vssd1 vccd1
+ vccd1 _08655_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07606_ _07616_/A _07613_/B _07608_/C vssd1 vssd1 vccd1 vccd1 _07607_/A sky130_fd_sc_hd__or3_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _12438_/Q vssd1 vssd1 vccd1 vccd1 _10097_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07537_ _07537_/A vssd1 vssd1 vccd1 vccd1 _07537_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07468_ _07468_/A vssd1 vssd1 vccd1 vccd1 _07478_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ _09210_/B _09201_/X _09206_/X vssd1 vssd1 vccd1 vccd1 _09207_/Y sky130_fd_sc_hd__o21ai_1
X_06419_ _06428_/A _06425_/B vssd1 vssd1 vccd1 vccd1 _06420_/A sky130_fd_sc_hd__or2_1
XFILLER_148_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07399_ _07822_/A _07404_/B _07401_/C vssd1 vssd1 vccd1 vccd1 _07400_/A sky130_fd_sc_hd__or3_1
XFILLER_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09138_ _14096_/Z vssd1 vssd1 vccd1 vccd1 _11160_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_151_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09069_ _11687_/C _12848_/Q _12849_/Q _12850_/Q _09067_/X _09068_/X vssd1 vssd1 vccd1
+ vccd1 _09069_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11100_ _11100_/A vssd1 vssd1 vccd1 vccd1 _12701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09707__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _10659_/A _12075_/X _12079_/X _12071_/X vssd1 vssd1 vccd1 vccd1 _12943_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11031_ _10377_/X _11027_/X _11030_/X _11024_/X vssd1 vssd1 vccd1 vccd1 _12678_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input12_A peripheralBus_address[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11933_ _11933_/A vssd1 vssd1 vccd1 vccd1 _12905_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11864_ _11898_/S vssd1 vssd1 vccd1 vccd1 _11878_/S sky130_fd_sc_hd__buf_2
X_13603_ _13603_/A _07357_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
X_10815_ _10870_/D _10878_/B _10803_/X vssd1 vssd1 vccd1 vccd1 _10815_/Y sky130_fd_sc_hd__o21ai_1
X_11795_ _14064_/Z _14000_/A _11805_/S vssd1 vssd1 vccd1 vccd1 _11796_/B sky130_fd_sc_hd__mux2_1
XFILLER_158_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13534_ _13534_/A _07532_/X vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10804__B1 _10803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10746_ _10746_/A vssd1 vssd1 vccd1 vccd1 _12615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13465_ _13465_/A _07715_/X vssd1 vssd1 vccd1 vccd1 _13625_/Z sky130_fd_sc_hd__ebufn_8
X_10677_ _13722_/A _10684_/B vssd1 vssd1 vccd1 vccd1 _10677_/X sky130_fd_sc_hd__or2_1
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12416_ _12470_/CLK _12416_/D vssd1 vssd1 vccd1 vccd1 _13592_/A sky130_fd_sc_hd__dfxtp_1
X_13396_ _13396_/A _08353_/X vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06306__A _09125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09973__A1 _09982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12347_ _12349_/CLK _12347_/D vssd1 vssd1 vccd1 vccd1 _12347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12278_ _12289_/CLK _12278_/D vssd1 vssd1 vccd1 vccd1 _12278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10770__B _10936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14017_ _14017_/A _08114_/X vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__ebufn_8
X_11229_ _11239_/A _11229_/B vssd1 vssd1 vccd1 vccd1 _11230_/A sky130_fd_sc_hd__and2_1
XFILLER_67_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06770_ _06809_/A vssd1 vssd1 vccd1 vccd1 _06780_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_64_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08440_ _12239_/Q vssd1 vssd1 vccd1 vccd1 _09317_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08371_ _12228_/Q _12229_/Q _12230_/Q _09210_/A _08368_/X _08370_/X vssd1 vssd1 vccd1
+ vccd1 _08371_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07322_ _07817_/A vssd1 vssd1 vccd1 vccd1 _08089_/B sky130_fd_sc_hd__buf_4
XANTENNA__07600__A _07615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10271__A1 _09763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07253_ _07253_/A _07263_/B _07260_/C vssd1 vssd1 vccd1 vccd1 _07254_/A sky130_fd_sc_hd__or3_1
X_07184_ _07184_/A vssd1 vssd1 vccd1 vccd1 _07184_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09964__A1 _09112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11776__B _13361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07973__C _07977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09825_ _09834_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__and2_1
XANTENNA_input4_A peripheralBus_address[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09756_ _10652_/A vssd1 vssd1 vccd1 vccd1 _09756_/X sky130_fd_sc_hd__buf_6
XFILLER_104_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06968_ _06972_/A _06977_/B vssd1 vssd1 vccd1 vccd1 _06969_/A sky130_fd_sc_hd__or2_1
XFILLER_101_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06886__A _06900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08707_ _12464_/Q vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _09687_/A vssd1 vssd1 vccd1 vccd1 _12349_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ _06899_/A vssd1 vssd1 vccd1 vccd1 _06899_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13276__432 vssd1 vssd1 vccd1 vccd1 _13276__432/HI _13981_/A sky130_fd_sc_hd__conb_1
XFILLER_161_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08638_ _12444_/Q vssd1 vssd1 vccd1 vccd1 _10099_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _08565_/X _08566_/X _08567_/X _08568_/X _08670_/A _08563_/X vssd1 vssd1 vccd1
+ vccd1 _08569_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10600_ _10600_/A vssd1 vssd1 vccd1 vccd1 _12579_/D sky130_fd_sc_hd__clkbuf_1
X_11580_ _11602_/C vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13317__473 vssd1 vssd1 vccd1 vccd1 _13317__473/HI _14054_/A sky130_fd_sc_hd__conb_1
X_10531_ _13686_/A _10535_/B vssd1 vssd1 vccd1 vccd1 _10531_/X sky130_fd_sc_hd__or2_1
XFILLER_155_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12990__146 vssd1 vssd1 vccd1 vccd1 _12990__146/HI _13387_/A sky130_fd_sc_hd__conb_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10462_ _10462_/A vssd1 vssd1 vccd1 vccd1 _12543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12201_ _10662_/A _12195_/X _12199_/X _12200_/X vssd1 vssd1 vccd1 vccd1 _12977_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10393_ _09756_/X _10379_/X _10392_/X _10383_/X vssd1 vssd1 vccd1 vccd1 _12522_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12132_ _12132_/A _12132_/B vssd1 vssd1 vccd1 vccd1 _12133_/A sky130_fd_sc_hd__and2_1
XFILLER_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12063_ _12101_/B vssd1 vssd1 vccd1 vccd1 _12073_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08060__B _08062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11014_ _12673_/Q _13947_/A vssd1 vssd1 vccd1 vccd1 _11016_/C sky130_fd_sc_hd__xor2_1
XFILLER_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06796__A _06809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09172__A _14007_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12965_ _12968_/CLK _12965_/D vssd1 vssd1 vccd1 vccd1 _12965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11916_ _12892_/Q _13364_/A vssd1 vssd1 vccd1 vccd1 _11920_/A sky130_fd_sc_hd__xor2_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12896_ _12914_/CLK _12896_/D vssd1 vssd1 vccd1 vccd1 _12896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _11898_/S vssd1 vssd1 vccd1 vccd1 _11861_/S sky130_fd_sc_hd__buf_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _12861_/Q _13366_/A vssd1 vssd1 vccd1 vccd1 _11780_/C sky130_fd_sc_hd__xor2_1
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07420__A _07468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13517_ _13517_/A _07576_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
X_10729_ _10414_/X _10690_/X _10728_/X _10711_/X vssd1 vssd1 vccd1 vccd1 _12611_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13448_ _13448_/A _07757_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10781__A _10820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ _13379_/A _08325_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[20] sky130_fd_sc_hd__ebufn_8
XFILLER_115_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_53_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__A _09347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13110__266 vssd1 vssd1 vccd1 vccd1 _13110__266/HI _13635_/A sky130_fd_sc_hd__conb_1
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07940_ _07940_/A vssd1 vssd1 vccd1 vccd1 _07940_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07871_ _07881_/A _07877_/B _07877_/C vssd1 vssd1 vccd1 vccd1 _07872_/A sky130_fd_sc_hd__or3_1
XFILLER_68_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09610_ _12200_/A _09610_/B _09610_/C vssd1 vssd1 vccd1 vccd1 _09611_/A sky130_fd_sc_hd__and3_1
XFILLER_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_68_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ _06822_/A _06830_/B _07234_/C vssd1 vssd1 vccd1 vccd1 _06823_/A sky130_fd_sc_hd__or3_1
XFILLER_56_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09541_ _13458_/A _12311_/Q _09610_/B vssd1 vssd1 vccd1 vccd1 _09542_/B sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_111_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06753_ _06753_/A vssd1 vssd1 vccd1 vccd1 _06765_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09472_ _12283_/Q _13559_/A vssd1 vssd1 vccd1 vccd1 _09473_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__07314__B _07317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004__160 vssd1 vssd1 vccd1 vccd1 _13004__160/HI _13415_/A sky130_fd_sc_hd__conb_1
X_06684_ _06686_/A _06692_/B _06692_/C vssd1 vssd1 vccd1 vccd1 _06685_/A sky130_fd_sc_hd__or3_1
XFILLER_64_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08423_ _12242_/Q _09316_/A _09322_/D _12245_/Q _08404_/X _08405_/X vssd1 vssd1 vccd1
+ vccd1 _08423_/X sky130_fd_sc_hd__mux4_2
XFILLER_11_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08354_ _08358_/A _08358_/B _08360_/C vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__or3_1
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07305_ _09484_/A vssd1 vssd1 vccd1 vccd1 _07781_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__07330__A _07371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08532__S1 _09146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08285_ _08288_/A _08285_/B vssd1 vssd1 vccd1 vccd1 _08286_/A sky130_fd_sc_hd__or2_1
XFILLER_149_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07236_ _11790_/A vssd1 vssd1 vccd1 vccd1 _09484_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10691__A _13775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07167_ _07167_/A vssd1 vssd1 vccd1 vccd1 _07167_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08161__A _08161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07098_ _07098_/A vssd1 vssd1 vccd1 vccd1 _07098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09808_ _09817_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09809_/A sky130_fd_sc_hd__and2_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09739_ _09739_/A vssd1 vssd1 vccd1 vccd1 _12357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11027__A _11055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _12768_/CLK _12750_/D vssd1 vssd1 vccd1 vccd1 _13877_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07224__B _07231_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _12853_/Q _11702_/B vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__or2_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12681_ _12682_/CLK _12681_/D vssd1 vssd1 vccd1 vccd1 _13810_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11632_/A _11632_/B _11639_/B _11632_/D vssd1 vssd1 vccd1 vccd1 _11633_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13053__209 vssd1 vssd1 vccd1 vccd1 _13053__209/HI _13512_/A sky130_fd_sc_hd__conb_1
X_11563_ _11563_/A _11572_/C vssd1 vssd1 vccd1 vccd1 _11563_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08055__B _08110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10514_ _13679_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _10514_/X sky130_fd_sc_hd__or2_1
X_11494_ _13978_/Z _11494_/B vssd1 vssd1 vccd1 vccd1 _11494_/X sky130_fd_sc_hd__or2_1
XANTENNA__09928__A1 _09124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ _10445_/A vssd1 vssd1 vccd1 vccd1 _12538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10376_ _10376_/A vssd1 vssd1 vccd1 vccd1 _12517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12115_ _12115_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _12116_/A sky130_fd_sc_hd__and2_1
XFILLER_112_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater114_A peripheralBus_data[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12046_ _12922_/Q _13361_/A vssd1 vssd1 vccd1 vccd1 _12050_/A sky130_fd_sc_hd__xor2_1
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09614__B _09918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output43_A _13786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07415__A _07417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13997_ _13997_/A _06289_/X vssd1 vssd1 vccd1 vccd1 _14125_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_1_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12948_ _12952_/CLK _12948_/D vssd1 vssd1 vccd1 vccd1 _14074_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12879_ _12904_/CLK _12879_/D vssd1 vssd1 vccd1 vccd1 _14007_/A sky130_fd_sc_hd__dfxtp_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10495__B _13758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08070_ _08081_/A _08077_/B _08070_/C vssd1 vssd1 vccd1 vccd1 _08071_/A sky130_fd_sc_hd__or3_1
X_07021_ _07033_/A vssd1 vssd1 vccd1 vccd1 _07031_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ _12821_/Q _11626_/A _11639_/C _12824_/Q _08918_/X _08919_/X vssd1 vssd1 vccd1
+ vccd1 _08972_/X sky130_fd_sc_hd__mux4_2
XFILLER_114_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07923_ _07923_/A vssd1 vssd1 vccd1 vccd1 _07999_/A sky130_fd_sc_hd__buf_2
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07854_ _07857_/A _07854_/B _08180_/B vssd1 vssd1 vccd1 vccd1 _07855_/A sky130_fd_sc_hd__or3_1
XANTENNA__07325__A _09918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06805_ _06805_/A vssd1 vssd1 vccd1 vccd1 _06805_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07785_ _07796_/A _07792_/B _07787_/C vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__or3_1
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09524_ _10548_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09524_/X sky130_fd_sc_hd__or2_1
X_06736_ _06746_/A _06738_/B _06738_/C vssd1 vssd1 vccd1 vccd1 _06737_/A sky130_fd_sc_hd__or3_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09455_/A _09455_/B vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__and2_1
XFILLER_101_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07979__B _07979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06667_ _11156_/B vssd1 vssd1 vccd1 vccd1 _06722_/A sky130_fd_sc_hd__clkbuf_4
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ _12245_/Q _09321_/D _12247_/Q _12248_/Q _08404_/X _08405_/X vssd1 vssd1 vccd1
+ vccd1 _08406_/X sky130_fd_sc_hd__mux4_2
X_09386_ _09388_/B _09388_/C _09385_/Y _09263_/X vssd1 vssd1 vccd1 vccd1 _12272_/D
+ sky130_fd_sc_hd__o211a_1
X_06598_ _06598_/A vssd1 vssd1 vccd1 vccd1 _06598_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07060__A _08364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13997__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ _08337_/A vssd1 vssd1 vccd1 vccd1 _08337_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08268_ _08276_/A _08274_/B _08276_/C vssd1 vssd1 vccd1 vccd1 _08269_/A sky130_fd_sc_hd__or3_1
XFILLER_20_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07219_ _07698_/A vssd1 vssd1 vccd1 vccd1 _07231_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08199_ _08199_/A vssd1 vssd1 vccd1 vccd1 _08199_/X sky130_fd_sc_hd__clkbuf_1
X_10230_ _12471_/Q _13746_/A vssd1 vssd1 vccd1 vccd1 _10232_/C sky130_fd_sc_hd__xor2_1
XFILLER_106_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10161_ _10161_/A vssd1 vssd1 vccd1 vccd1 _12467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10092_ _10092_/A vssd1 vssd1 vccd1 vccd1 _12450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13920_ _13920_/A _06500_/X vssd1 vssd1 vccd1 vccd1 _14112_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13851_ _13851_/A _06693_/X vssd1 vssd1 vccd1 vccd1 _13979_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11980__A _11998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ _12802_/CLK _12802_/D vssd1 vssd1 vccd1 vccd1 _13976_/A sky130_fd_sc_hd__dfxtp_1
X_13782_ _13782_/A _06885_/X vssd1 vssd1 vccd1 vccd1 _13974_/Z sky130_fd_sc_hd__ebufn_8
X_10994_ _11078_/A _10994_/B vssd1 vssd1 vccd1 vccd1 _10995_/A sky130_fd_sc_hd__and2_1
XFILLER_27_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12733_ _12753_/CLK _12733_/D vssd1 vssd1 vccd1 vccd1 _12733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11653__B1 _11569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996__152 vssd1 vssd1 vccd1 vccd1 _12996__152/HI _13407_/A sky130_fd_sc_hd__conb_1
X_12664_ _12853_/CLK _12664_/D vssd1 vssd1 vccd1 vccd1 _12664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _11630_/D _11616_/C _11614_/Y vssd1 vssd1 vccd1 vccd1 _12833_/D sky130_fd_sc_hd__a21oi_1
XFILLER_156_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12595_ _12800_/CLK _12595_/D vssd1 vssd1 vccd1 vccd1 _13722_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11546_ _11563_/A _11546_/B vssd1 vssd1 vccd1 vccd1 _12816_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11477_ _11477_/A vssd1 vssd1 vccd1 vccd1 _12797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10762__C _10820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10428_ _13786_/A _10555_/B vssd1 vssd1 vccd1 vccd1 _10480_/S sky130_fd_sc_hd__and2_2
XFILLER_98_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _12507_/Q _13749_/A vssd1 vssd1 vccd1 vccd1 _10362_/B sky130_fd_sc_hd__xor2_1
XFILLER_97_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13181__337 vssd1 vssd1 vccd1 vccd1 _13181__337/HI _13774_/A sky130_fd_sc_hd__conb_1
X_12029_ _12934_/Q _14077_/A _12029_/S vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__mux2_1
XFILLER_120_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13222__378 vssd1 vssd1 vccd1 vccd1 _13222__378/HI _13861_/A sky130_fd_sc_hd__conb_1
XFILLER_66_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07570_ _07575_/A _08103_/B _07580_/C vssd1 vssd1 vccd1 vccd1 _07571_/A sky130_fd_sc_hd__or3_1
XFILLER_19_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06521_ _06521_/A _06526_/B _06526_/C vssd1 vssd1 vccd1 vccd1 _06522_/A sky130_fd_sc_hd__or3_1
X_09240_ _09317_/B _09242_/C _09206_/X vssd1 vssd1 vccd1 vccd1 _09240_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06452_ _06452_/A vssd1 vssd1 vccd1 vccd1 _06452_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13075__231 vssd1 vssd1 vccd1 vccd1 _13075__231/HI _13550_/A sky130_fd_sc_hd__conb_1
X_09171_ _10662_/A _09145_/X _09170_/X _09148_/X vssd1 vssd1 vccd1 vccd1 _12221_/D
+ sky130_fd_sc_hd__a211o_1
X_06383_ _06391_/A _08349_/A vssd1 vssd1 vccd1 vccd1 _06384_/A sky130_fd_sc_hd__or2_1
XFILLER_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08122_ _08122_/A _08128_/B _08122_/C vssd1 vssd1 vccd1 vccd1 _08123_/A sky130_fd_sc_hd__or3_1
XFILLER_147_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116__272 vssd1 vssd1 vccd1 vccd1 _13116__272/HI _13641_/A sky130_fd_sc_hd__conb_1
XFILLER_162_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08053_ _08053_/A vssd1 vssd1 vccd1 vccd1 _08053_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07004_ _07004_/A vssd1 vssd1 vccd1 vccd1 _07004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11784__B _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ _12824_/Q _12825_/Q _12826_/Q _12827_/Q _08928_/X _08929_/X vssd1 vssd1 vccd1
+ vccd1 _08955_/X sky130_fd_sc_hd__mux4_2
XFILLER_102_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07906_ _11154_/B vssd1 vssd1 vccd1 vccd1 _07917_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08886_ _08886_/A vssd1 vssd1 vccd1 vccd1 _10697_/A sky130_fd_sc_hd__buf_4
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07837_ _07843_/A _07840_/B _08180_/C vssd1 vssd1 vccd1 vccd1 _07838_/A sky130_fd_sc_hd__or3_1
X_07768_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07779_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__06894__A _07328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ _13430_/A _09500_/X _09506_/X _09496_/X vssd1 vssd1 vccd1 vccd1 _12299_/D
+ sky130_fd_sc_hd__o211a_1
X_06719_ _06733_/A _06719_/B _06719_/C vssd1 vssd1 vccd1 vccd1 _06720_/A sky130_fd_sc_hd__or3_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _07699_/A _07710_/B _07704_/C vssd1 vssd1 vccd1 vccd1 _07700_/A sky130_fd_sc_hd__or3_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _13433_/A _12285_/Q _09448_/S vssd1 vssd1 vccd1 vccd1 _09439_/B sky130_fd_sc_hd__mux2_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _09369_/A _09382_/B vssd1 vssd1 vccd1 vccd1 _12267_/D sky130_fd_sc_hd__nor2_1
X_11400_ _11400_/A _11400_/B _11400_/C _11400_/D vssd1 vssd1 vccd1 vccd1 _11406_/B
+ sky130_fd_sc_hd__or4_1
X_12380_ _12386_/CLK _12380_/D vssd1 vssd1 vccd1 vccd1 _12380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ _11344_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11332_/A sky130_fd_sc_hd__and2_1
XFILLER_126_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14050_ _14050_/A _07914_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
XFILLER_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11262_ _12738_/Q _13946_/A vssd1 vssd1 vccd1 vccd1 _11262_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10213_ _10213_/A vssd1 vssd1 vccd1 vccd1 _12480_/D sky130_fd_sc_hd__clkbuf_1
X_11193_ _11061_/X _11185_/X _11192_/X _11180_/X vssd1 vssd1 vccd1 vccd1 _12723_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10374__B1 _13761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10144_ _10148_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__or2_1
XFILLER_121_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10075_ _10073_/Y _10070_/C _10074_/Y vssd1 vssd1 vccd1 vccd1 _12447_/D sky130_fd_sc_hd__o21a_1
XFILLER_48_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13903_ _13903_/A _07855_/X vssd1 vssd1 vccd1 vccd1 _14063_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13834_ _13834_/A _06739_/X vssd1 vssd1 vccd1 vccd1 _13994_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13765_ _13765_/A _06930_/X vssd1 vssd1 vccd1 vccd1 _13765_/Z sky130_fd_sc_hd__ebufn_8
X_13059__215 vssd1 vssd1 vccd1 vccd1 _13059__215/HI _13518_/A sky130_fd_sc_hd__conb_1
X_10977_ _10986_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__and2_1
X_12716_ _12722_/CLK _12716_/D vssd1 vssd1 vccd1 vccd1 _13844_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_149_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13696_ _13696_/A _07102_/X vssd1 vssd1 vccd1 vccd1 _14112_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12647_ _12647_/CLK _12647_/D vssd1 vssd1 vccd1 vccd1 _12647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12578_ _12800_/CLK _12578_/D vssd1 vssd1 vccd1 vccd1 _12578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11529_ _11625_/C _11531_/C _11521_/X vssd1 vssd1 vccd1 vccd1 _11530_/B sky130_fd_sc_hd__o21ai_1
XFILLER_7_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06979__A _07417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _08887_/A vssd1 vssd1 vccd1 vccd1 _08740_/X sky130_fd_sc_hd__buf_2
XFILLER_100_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater102 _14117_/Z vssd1 vssd1 vccd1 vccd1 _13765_/Z sky130_fd_sc_hd__buf_12
XFILLER_112_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater113 peripheralBus_data[18] vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__buf_12
Xrepeater124 _14108_/Z vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__buf_12
Xrepeater135 peripheralBus_data[10] vssd1 vssd1 vccd1 vccd1 _14009_/Z sky130_fd_sc_hd__buf_12
X_08671_ _08626_/X _08631_/X _08628_/X _08637_/X _08663_/X _08670_/X vssd1 vssd1 vccd1
+ vccd1 _08671_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07622_ _07622_/A vssd1 vssd1 vccd1 vccd1 _07622_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07603__A _07603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07553_ _07553_/A vssd1 vssd1 vccd1 vccd1 _07564_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06504_ _06504_/A vssd1 vssd1 vccd1 vccd1 _06504_/X sky130_fd_sc_hd__clkbuf_1
X_07484_ _08089_/A _07484_/B vssd1 vssd1 vccd1 vccd1 _07485_/A sky130_fd_sc_hd__or2_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ _09223_/A _09223_/B vssd1 vssd1 vccd1 vccd1 _12233_/D sky130_fd_sc_hd__nor2_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06435_ _06440_/A _06437_/B vssd1 vssd1 vccd1 vccd1 _06436_/A sky130_fd_sc_hd__or2_1
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09154_ _14067_/Z vssd1 vssd1 vccd1 vccd1 _09625_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11779__B _13371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06366_ _06547_/A vssd1 vssd1 vccd1 vccd1 _07822_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_163_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08105_ _08110_/A _08113_/B _08105_/C vssd1 vssd1 vccd1 vccd1 _08106_/A sky130_fd_sc_hd__or3_1
XFILLER_162_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _10941_/C vssd1 vssd1 vccd1 vccd1 _13949_/A sky130_fd_sc_hd__buf_6
XFILLER_108_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06297_ _06303_/A _06308_/B _06308_/C vssd1 vssd1 vccd1 vccd1 _06298_/A sky130_fd_sc_hd__or3_1
X_08036_ _11283_/B vssd1 vssd1 vccd1 vccd1 _08047_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09987_ _10077_/A vssd1 vssd1 vccd1 vccd1 _09987_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08938_ _10939_/A vssd1 vssd1 vccd1 vccd1 _13935_/A sky130_fd_sc_hd__buf_6
XANTENNA__11019__B _13943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ _10164_/B vssd1 vssd1 vccd1 vccd1 _13752_/A sky130_fd_sc_hd__buf_4
XFILLER_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10900_ _10907_/C _10900_/B vssd1 vssd1 vccd1 vccd1 _10903_/B sky130_fd_sc_hd__and2_1
X_11880_ _11880_/A vssd1 vssd1 vccd1 vccd1 _12896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11608__B1 _11540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ _10870_/B _10828_/A _10830_/Y vssd1 vssd1 vccd1 vccd1 _12634_/D sky130_fd_sc_hd__a21oi_1
XFILLER_16_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ _13550_/A _07489_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10762_ _10767_/C _10762_/B _10820_/C vssd1 vssd1 vccd1 vccd1 _10763_/A sky130_fd_sc_hd__and3b_1
XFILLER_158_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12501_ _12505_/CLK _12501_/D vssd1 vssd1 vccd1 vccd1 _12501_/Q sky130_fd_sc_hd__dfxtp_1
X_13481_ _13481_/A _07670_/X vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_8
X_10693_ _10693_/A _11412_/C _10693_/C vssd1 vssd1 vccd1 vccd1 _10732_/B sky130_fd_sc_hd__nor3_4
X_12432_ _12617_/CLK _12432_/D vssd1 vssd1 vccd1 vccd1 _12432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08788__A0 _08781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12363_ _12369_/CLK _12363_/D vssd1 vssd1 vccd1 vccd1 _13492_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _14102_/A _08217_/X vssd1 vssd1 vccd1 vccd1 _14102_/Z sky130_fd_sc_hd__ebufn_8
X_11314_ _13881_/A _11323_/B vssd1 vssd1 vccd1 vccd1 _11314_/X sky130_fd_sc_hd__or2_1
X_12294_ _12295_/CLK _12294_/D vssd1 vssd1 vccd1 vccd1 _13425_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14033_ _14033_/A _07869_/X vssd1 vssd1 vccd1 vccd1 _14033_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_113_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11245_ _13883_/A _12739_/Q _11248_/S vssd1 vssd1 vccd1 vccd1 _11246_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09175__A input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _10659_/X _11171_/X _11175_/X _11166_/X vssd1 vssd1 vccd1 vccd1 _12717_/D
+ sky130_fd_sc_hd__o211a_1
X_10127_ _10146_/A _10127_/B _10127_/C vssd1 vssd1 vccd1 vccd1 _10128_/A sky130_fd_sc_hd__and3_1
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09903__A _09915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ _10088_/C _10060_/C _10123_/A vssd1 vssd1 vccd1 vccd1 _10058_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13817_ _13817_/A _06787_/X vssd1 vssd1 vccd1 vccd1 _14009_/Z sky130_fd_sc_hd__ebufn_8
X_13293__449 vssd1 vssd1 vccd1 vccd1 _13293__449/HI _13998_/A sky130_fd_sc_hd__conb_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08238__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13748_ _13748_/A _06971_/X vssd1 vssd1 vccd1 vccd1 _14100_/Z sky130_fd_sc_hd__ebufn_8
X_13679_ _13679_/A _07990_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[0] sky130_fd_sc_hd__ebufn_8
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08254__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13187__343 vssd1 vssd1 vccd1 vccd1 _13187__343/HI _13794_/A sky130_fd_sc_hd__conb_1
XFILLER_104_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09910_ _09092_/X _09902_/X _09909_/X _09905_/X vssd1 vssd1 vccd1 vccd1 _12403_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08626__S0 _08549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09841_ _10173_/A _09841_/B vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__and2_1
XFILLER_113_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06502__A _08276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13228__384 vssd1 vssd1 vccd1 vccd1 _13228__384/HI _13867_/A sky130_fd_sc_hd__conb_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09772_ _09770_/X _09759_/X _09771_/X _09765_/X vssd1 vssd1 vccd1 vccd1 _12366_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07317__B _07317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ _10639_/A vssd1 vssd1 vccd1 vccd1 _10637_/A sky130_fd_sc_hd__clkbuf_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08723_ _09399_/C vssd1 vssd1 vccd1 vccd1 _13565_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_repeater76_A _14035_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08654_ _12453_/Q _12454_/Q _12455_/Q _12456_/Q _08556_/X _08557_/X vssd1 vssd1 vccd1
+ vccd1 _08654_/X sky130_fd_sc_hd__mux4_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07605_ _07661_/A vssd1 vssd1 vccd1 vccd1 _07616_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08585_ _08573_/X _08577_/X _08580_/X _08582_/X _08583_/X _08584_/X vssd1 vssd1 vccd1
+ vccd1 _08585_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11066__A1 _11064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ _07545_/A _07545_/B _07538_/C vssd1 vssd1 vccd1 vccd1 _07537_/A sky130_fd_sc_hd__or3_1
XFILLER_149_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07467_ _07467_/A vssd1 vssd1 vccd1 vccd1 _07467_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10694__A _10732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09206_/X sky130_fd_sc_hd__clkbuf_4
X_06418_ _06442_/A vssd1 vssd1 vccd1 vccd1 _06428_/A sky130_fd_sc_hd__clkbuf_1
X_07398_ _07964_/A vssd1 vssd1 vccd1 vccd1 _07822_/A sky130_fd_sc_hd__clkbuf_4
X_09137_ _09124_/X _09130_/X _09136_/X _09109_/X vssd1 vssd1 vccd1 vccd1 _12214_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06349_ _06359_/A _06349_/B _06349_/C vssd1 vssd1 vccd1 vccd1 _06350_/A sky130_fd_sc_hd__or3_1
XFILLER_5_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09068_ _09068_/A vssd1 vssd1 vccd1 vccd1 _09068_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08019_ _08072_/A vssd1 vssd1 vccd1 vccd1 _08030_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11030_ _13807_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11030_/X sky130_fd_sc_hd__or2_1
XFILLER_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12981_ _12981_/CLK _12981_/D vssd1 vssd1 vccd1 vccd1 _14106_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11932_ _11945_/A _11932_/B vssd1 vssd1 vccd1 vccd1 _11933_/A sky130_fd_sc_hd__and2_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _11863_/A vssd1 vssd1 vccd1 vccd1 _12891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13602_ _13602_/A _07360_/X vssd1 vssd1 vccd1 vccd1 _13666_/Z sky130_fd_sc_hd__ebufn_8
X_13021__177 vssd1 vssd1 vccd1 vccd1 _13021__177/HI _13448_/A sky130_fd_sc_hd__conb_1
X_10814_ _10874_/C vssd1 vssd1 vccd1 vccd1 _10870_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_11794_ _11794_/A vssd1 vssd1 vccd1 vccd1 _12871_/D sky130_fd_sc_hd__clkbuf_1
X_13533_ _13533_/A _07537_/X vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__ebufn_8
X_10745_ _10742_/X _10745_/B _10917_/B vssd1 vssd1 vccd1 vccd1 _10746_/A sky130_fd_sc_hd__and3b_1
XFILLER_9_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13464_ _13464_/A _07718_/X vssd1 vssd1 vccd1 vccd1 _14104_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10676_ _10408_/X _10673_/X _10675_/X _10668_/X vssd1 vssd1 vccd1 vccd1 _12594_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12415_ _12470_/CLK _12415_/D vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__dfxtp_1
X_13395_ _13395_/A _08355_/X vssd1 vssd1 vccd1 vccd1 _14035_/Z sky130_fd_sc_hd__ebufn_8
X_12346_ _12349_/CLK _12346_/D vssd1 vssd1 vccd1 vccd1 _12346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12277_ _12289_/CLK _12277_/D vssd1 vssd1 vccd1 vccd1 _12277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14016_ _14016_/A _08119_/X vssd1 vssd1 vccd1 vccd1 _14112_/Z sky130_fd_sc_hd__ebufn_8
X_11228_ _13878_/A _12734_/Q _11231_/S vssd1 vssd1 vccd1 vccd1 _11229_/B sky130_fd_sc_hd__mux2_1
XFILLER_141_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12043__B _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11159_ _11153_/X _11155_/X _11158_/X _11068_/X vssd1 vssd1 vccd1 vccd1 _12711_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09633__A _09633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__A1 _10648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10498__B _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11048__A1 _10662_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08370_ _08525_/A vssd1 vssd1 vccd1 vccd1 _08370_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07321_ _09484_/B vssd1 vssd1 vccd1 vccd1 _07817_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07252_ _07291_/A vssd1 vssd1 vccd1 vccd1 _07263_/B sky130_fd_sc_hd__clkbuf_1
X_07183_ _07193_/A _07190_/B _07187_/C vssd1 vssd1 vccd1 vccd1 _07184_/A sky130_fd_sc_hd__or3_1
XFILLER_157_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07328__A _07328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09824_ _13528_/A _12383_/Q _09837_/S vssd1 vssd1 vccd1 vccd1 _09825_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09755_ _09753_/X _09741_/X _09754_/X _09748_/X vssd1 vssd1 vccd1 vccd1 _12361_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06967_ _06967_/A vssd1 vssd1 vccd1 vccd1 _06977_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_100_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10689__A _10706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08706_ _12463_/Q vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09686_ _09686_/A _09686_/B vssd1 vssd1 vccd1 vccd1 _09687_/A sky130_fd_sc_hd__and2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08159__A _08177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06898_ _07328_/A _06898_/B _06898_/C vssd1 vssd1 vccd1 vccd1 _06899_/A sky130_fd_sc_hd__or3_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07063__A _08177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _10052_/C _10052_/B _10052_/A _10099_/D _08629_/X _08630_/X vssd1 vssd1 vccd1
+ vccd1 _08637_/X sky130_fd_sc_hd__mux4_2
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08568_ _12449_/Q _12450_/Q _12451_/Q _12452_/Q _08559_/X _08560_/X vssd1 vssd1 vccd1
+ vccd1 _08568_/X sky130_fd_sc_hd__mux4_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07519_ _07519_/A vssd1 vssd1 vccd1 vccd1 _07531_/A sky130_fd_sc_hd__clkbuf_1
X_08499_ _11707_/A vssd1 vssd1 vccd1 vccd1 _13367_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11313__A _11325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10530_ _09763_/X _10525_/X _10529_/X _10523_/X vssd1 vssd1 vccd1 vccd1 _12557_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _10461_/A _10461_/B vssd1 vssd1 vccd1 vccd1 _10462_/A sky130_fd_sc_hd__and2_1
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12200_ _12200_/A vssd1 vssd1 vccd1 vccd1 _12200_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10392_ _13651_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__or2_1
XFILLER_163_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12131_ _12961_/Q _14103_/A _12135_/S vssd1 vssd1 vccd1 vccd1 _12132_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07238__A _07291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ _12062_/A _12062_/B _12059_/Y vssd1 vssd1 vccd1 vccd1 _12101_/B sky130_fd_sc_hd__nor3b_2
X_11013_ _12676_/Q _13950_/A vssd1 vssd1 vccd1 vccd1 _11016_/B sky130_fd_sc_hd__xor2_1
XFILLER_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12964_ _12968_/CLK _12964_/D vssd1 vssd1 vccd1 vccd1 _12964_/Q sky130_fd_sc_hd__dfxtp_1
X_11915_ _11915_/A _11915_/B _11915_/C _11915_/D vssd1 vssd1 vccd1 vccd1 _11921_/B
+ sky130_fd_sc_hd__or4_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07404__C _07496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12895_/CLK _12895_/D vssd1 vssd1 vccd1 vccd1 _12895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _13403_/A _12103_/B vssd1 vssd1 vccd1 vccd1 _11898_/S sky130_fd_sc_hd__nand2_2
XFILLER_159_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _12869_/Q _13374_/A vssd1 vssd1 vccd1 vccd1 _11780_/B sky130_fd_sc_hd__xor2_1
XFILLER_159_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11223__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13516_ _13516_/A _07579_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
X_10728_ _13786_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10728_/X sky130_fd_sc_hd__or2_1
XFILLER_158_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12038__B _13372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ _13447_/A _07760_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
X_10659_ _10659_/A vssd1 vssd1 vccd1 vccd1 _10659_/X sky130_fd_sc_hd__buf_6
XFILLER_127_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09628__A _09655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ _13378_/A _08322_/X vssd1 vssd1 vccd1 vccd1 _13666_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12329_ _12331_/CLK _12329_/D vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07870_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07881_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10713__A0 _13973_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06821_ _06967_/A vssd1 vssd1 vccd1 vccd1 _07234_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09096__D_N input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13299__455 vssd1 vssd1 vccd1 vccd1 _13299__455/HI _14020_/A sky130_fd_sc_hd__conb_1
X_09540_ _09540_/A vssd1 vssd1 vccd1 vccd1 _12310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06752_ _06752_/A vssd1 vssd1 vccd1 vccd1 _06752_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09471_ _12290_/Q _13566_/A vssd1 vssd1 vccd1 vccd1 _09473_/C sky130_fd_sc_hd__xnor2_1
X_06683_ _06683_/A vssd1 vssd1 vccd1 vccd1 _06683_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08422_ _12243_/Q vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08353_ _08353_/A vssd1 vssd1 vccd1 vccd1 _08353_/X sky130_fd_sc_hd__clkbuf_1
X_07304_ _07304_/A vssd1 vssd1 vccd1 vccd1 _07304_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11441__A1 _11184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08284_ _08284_/A vssd1 vssd1 vccd1 vccd1 _08284_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07235_ _07235_/A vssd1 vssd1 vccd1 vccd1 _07235_/X sky130_fd_sc_hd__clkbuf_1
X_07166_ _07166_/A _07177_/B _07173_/C vssd1 vssd1 vccd1 vccd1 _07167_/A sky130_fd_sc_hd__or3_1
X_07097_ _07108_/A _07105_/B _07101_/C vssd1 vssd1 vccd1 vccd1 _07098_/A sky130_fd_sc_hd__or3_1
XFILLER_160_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09807_ _13523_/A _12378_/Q _09820_/S vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__mux2_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07999_ _07999_/A vssd1 vssd1 vccd1 vccd1 _08010_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09738_ _12200_/A _09738_/B _09738_/C vssd1 vssd1 vccd1 vccd1 _09739_/A sky130_fd_sc_hd__and3_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09669_ _09669_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _09670_/A sky130_fd_sc_hd__and2_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11700_/A _11702_/B vssd1 vssd1 vccd1 vccd1 _12852_/D sky130_fd_sc_hd__nor2_1
XANTENNA__13523__A _13523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12680_ _12682_/CLK _12680_/D vssd1 vssd1 vccd1 vccd1 _13809_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11641_/C _11631_/B _11631_/C _11631_/D vssd1 vssd1 vccd1 vccd1 _11633_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__07521__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13092__248 vssd1 vssd1 vccd1 vccd1 _13092__248/HI _13601_/A sky130_fd_sc_hd__conb_1
X_11562_ _11625_/A _11625_/B _11562_/C _11627_/B vssd1 vssd1 vccd1 vccd1 _11572_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10513_ _10553_/B vssd1 vssd1 vccd1 vccd1 _10522_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11493_ _13977_/A _11459_/X _11492_/X _11464_/X vssd1 vssd1 vccd1 vccd1 _12803_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13133__289 vssd1 vssd1 vccd1 vccd1 _13133__289/HI _13674_/A sky130_fd_sc_hd__conb_1
X_10444_ _10444_/A _10444_/B vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__and2_1
XFILLER_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08352__A _08358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10375_ _11151_/A _10375_/B _10375_/C vssd1 vssd1 vccd1 vccd1 _10376_/A sky130_fd_sc_hd__and3_1
XFILLER_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12114_ _12956_/Q _14098_/A _12118_/S vssd1 vssd1 vccd1 vccd1 _12115_/B sky130_fd_sc_hd__mux2_1
XFILLER_151_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12045_ _12045_/A _12045_/B _12045_/C _12045_/D vssd1 vssd1 vccd1 vccd1 _12056_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_78_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater107_A peripheralBus_data[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09183__A _13401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09614__C _12062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13027__183 vssd1 vssd1 vccd1 vccd1 _13027__183/HI _13454_/A sky130_fd_sc_hd__conb_1
X_13996_ _13996_/A _06292_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA_output36_A _13403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12947_ _12952_/CLK _12947_/D vssd1 vssd1 vccd1 vccd1 _14073_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12904_/CLK _12878_/D vssd1 vssd1 vccd1 vccd1 _14006_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11829_ _11829_/A vssd1 vssd1 vccd1 vccd1 _12881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08246__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07020_ _07020_/A vssd1 vssd1 vccd1 vccd1 _07020_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08971_ _12822_/Q vssd1 vssd1 vccd1 vccd1 _11626_/A sky130_fd_sc_hd__clkbuf_2
X_07922_ _07922_/A vssd1 vssd1 vccd1 vccd1 _07922_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09093__A input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ _07853_/A vssd1 vssd1 vccd1 vccd1 _07853_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06804_ _07857_/A _06806_/B _06806_/C vssd1 vssd1 vccd1 vccd1 _06805_/A sky130_fd_sc_hd__or3_1
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07784_ _07798_/A vssd1 vssd1 vccd1 vccd1 _07796_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10032__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__B1 _09392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09523_ _13436_/A _09513_/X _09521_/X _09522_/X vssd1 vssd1 vccd1 vccd1 _12305_/D
+ sky130_fd_sc_hd__o211a_1
X_06735_ _06748_/A vssd1 vssd1 vccd1 vccd1 _06746_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09454_ _13438_/A _12290_/Q _09454_/S vssd1 vssd1 vccd1 vccd1 _09455_/B sky130_fd_sc_hd__mux2_1
X_06666_ _06680_/A vssd1 vssd1 vccd1 vccd1 _06678_/B sky130_fd_sc_hd__clkbuf_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10686__B _10686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08405_ _13393_/A vssd1 vssd1 vccd1 vccd1 _08405_/X sky130_fd_sc_hd__clkbuf_2
X_09385_ _09388_/B _09388_/C vssd1 vssd1 vccd1 vccd1 _09385_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06597_ _06597_/A _06602_/B _06602_/C vssd1 vssd1 vccd1 vccd1 _06598_/A sky130_fd_sc_hd__or3_1
XANTENNA__07060__B _07995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _08336_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08337_/A sky130_fd_sc_hd__or2_1
XFILLER_165_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07995__B _07995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ _08351_/A vssd1 vssd1 vccd1 vccd1 _08276_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_165_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07218_ _09614_/A vssd1 vssd1 vccd1 vccd1 _07698_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08198_ _08198_/A _08208_/B _08198_/C vssd1 vssd1 vccd1 vccd1 _08199_/A sky130_fd_sc_hd__or3_1
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07149_ _11924_/A vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__buf_2
XFILLER_133_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10160_ _10160_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__and2_1
XFILLER_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09715__B _09848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _10094_/B _10135_/B _10091_/C vssd1 vssd1 vccd1 vccd1 _10092_/A sky130_fd_sc_hd__and3b_1
XFILLER_75_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11038__A _13811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13850_ _13850_/A _06698_/X vssd1 vssd1 vccd1 vccd1 _13978_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12801_ _12811_/CLK _12801_/D vssd1 vssd1 vccd1 vccd1 _13975_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10993_ _13821_/A _12675_/Q _10996_/S vssd1 vssd1 vccd1 vccd1 _10994_/B sky130_fd_sc_hd__mux2_1
X_13781_ _13781_/A _06889_/X vssd1 vssd1 vccd1 vccd1 _13973_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_43_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12768_/CLK _12732_/D vssd1 vssd1 vccd1 vccd1 _12732_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_52_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12687_/CLK _12663_/D vssd1 vssd1 vccd1 vccd1 _12663_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _11630_/D _11616_/C _11505_/B vssd1 vssd1 vccd1 vccd1 _11614_/Y sky130_fd_sc_hd__o21ai_1
X_12594_ _12800_/CLK _12594_/D vssd1 vssd1 vccd1 vccd1 _13721_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11545_ _11627_/C _11542_/A _11540_/X vssd1 vssd1 vccd1 vccd1 _11546_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_67_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09178__A _09638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11476_ _11481_/A _11476_/B vssd1 vssd1 vccd1 vccd1 _11477_/A sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_110_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10427_ _10479_/A vssd1 vssd1 vccd1 vccd1 _10444_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10358_ _12511_/Q _13753_/A vssd1 vssd1 vccd1 vccd1 _10362_/A sky130_fd_sc_hd__xor2_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _13628_/A _10291_/B vssd1 vssd1 vccd1 vccd1 _10289_/X sky130_fd_sc_hd__or2_1
XFILLER_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12028_ _12028_/A vssd1 vssd1 vccd1 vccd1 _12933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12051__B _13364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09641__A _09655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13979_ _13979_/A _06343_/X vssd1 vssd1 vccd1 vccd1 _13979_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_81_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06520_ _06520_/A vssd1 vssd1 vccd1 vccd1 _06520_/X sky130_fd_sc_hd__clkbuf_1
X_06451_ _06451_/A _07845_/B vssd1 vssd1 vccd1 vccd1 _06452_/A sky130_fd_sc_hd__or2_1
XFILLER_61_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ _13398_/A _09179_/B vssd1 vssd1 vccd1 vccd1 _09170_/X sky130_fd_sc_hd__and2_1
X_06382_ _06382_/A vssd1 vssd1 vccd1 vccd1 _06382_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08121_ _08121_/A vssd1 vssd1 vccd1 vccd1 _08121_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ _08052_/A _08110_/B _08057_/C vssd1 vssd1 vccd1 vccd1 _08053_/A sky130_fd_sc_hd__or3_1
X_07003_ _07007_/A _07007_/B vssd1 vssd1 vccd1 vccd1 _07004_/A sky130_fd_sc_hd__or2_1
XANTENNA__11130__B _13936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08954_ _08943_/X _08948_/X _08950_/X _08951_/X _08952_/X _08953_/X vssd1 vssd1 vccd1
+ vccd1 _08954_/X sky130_fd_sc_hd__mux4_1
X_07905_ _09614_/A vssd1 vssd1 vccd1 vccd1 _11154_/B sky130_fd_sc_hd__buf_6
X_08885_ _12656_/Q vssd1 vssd1 vccd1 vccd1 _10921_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07836_ _07836_/A vssd1 vssd1 vccd1 vccd1 _07836_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07767_ _07767_/A vssd1 vssd1 vccd1 vccd1 _07767_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10697__A _10697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13355__511 vssd1 vssd1 vccd1 vccd1 _13355__511/HI _14124_/A sky130_fd_sc_hd__conb_1
X_09506_ _09633_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09506_/X sky130_fd_sc_hd__or2_1
X_06718_ _06718_/A vssd1 vssd1 vccd1 vccd1 _06718_/X sky130_fd_sc_hd__clkbuf_1
X_07698_ _07698_/A vssd1 vssd1 vccd1 vccd1 _07710_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09437_ _09437_/A vssd1 vssd1 vccd1 vccd1 _12284_/D sky130_fd_sc_hd__clkbuf_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06649_ _06659_/A _06651_/B _06651_/C vssd1 vssd1 vccd1 vccd1 _06650_/A sky130_fd_sc_hd__or3_1
XANTENNA__12373__CLK _12555_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09368_ _09368_/A _09368_/B _09368_/C _09368_/D vssd1 vssd1 vccd1 vccd1 _09382_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_165_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08319_ _08324_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08320_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_113_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _12301_/CLK sky130_fd_sc_hd__clkbuf_16
X_09299_ _09299_/A _09299_/B vssd1 vssd1 vccd1 vccd1 _12252_/D sky130_fd_sc_hd__nor2_1
X_11330_ _13903_/A _12760_/Q _11408_/B vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06415__A _06913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11261_ _12728_/Q _11388_/B vssd1 vssd1 vccd1 vccd1 _11261_/X sky130_fd_sc_hd__and2_1
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10212_ _10298_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10213_/A sky130_fd_sc_hd__and2_1
X_11192_ _13851_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11192_/X sky130_fd_sc_hd__or2_1
XFILLER_133_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10143_ _10143_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _12462_/D sky130_fd_sc_hd__nor2_1
XFILLER_153_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10074_ _10073_/Y _10070_/C _10160_/A vssd1 vssd1 vccd1 vccd1 _10074_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_75_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13902_ _13902_/A _06553_/X vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_75_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13833_ _13833_/A _06743_/X vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13098__254 vssd1 vssd1 vccd1 vccd1 _13098__254/HI _13607_/A sky130_fd_sc_hd__conb_1
X_13764_ _13764_/A _06933_/X vssd1 vssd1 vccd1 vccd1 _13988_/Z sky130_fd_sc_hd__ebufn_8
X_10976_ _13816_/A _12670_/Q _10990_/S vssd1 vssd1 vccd1 vccd1 _10977_/B sky130_fd_sc_hd__mux2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12715_ _12722_/CLK _12715_/D vssd1 vssd1 vccd1 vccd1 _13843_/A sky130_fd_sc_hd__dfxtp_1
X_13695_ _13695_/A _07106_/X vssd1 vssd1 vccd1 vccd1 _14079_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12646_ _12646_/CLK _12646_/D vssd1 vssd1 vccd1 vccd1 _12646_/Q sky130_fd_sc_hd__dfxtp_1
X_13139__295 vssd1 vssd1 vccd1 vccd1 _13139__295/HI _13696_/A sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_104_clk _12217_/CLK vssd1 vssd1 vccd1 vccd1 _12325_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12577_ _12597_/CLK _12577_/D vssd1 vssd1 vccd1 vccd1 _12577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ _11625_/C _11531_/C vssd1 vssd1 vccd1 vccd1 _11530_/A sky130_fd_sc_hd__and2_1
XFILLER_144_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06325__A _06462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12046__B _13361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11459_ _11459_/A vssd1 vssd1 vccd1 vccd1 _11459_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09636__A _09636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06979__B _07969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12062__A _12062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater103 peripheralBus_data[22] vssd1 vssd1 vccd1 vccd1 _14117_/Z sky130_fd_sc_hd__buf_12
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater114 peripheralBus_data[18] vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__buf_12
Xrepeater125 peripheralBus_data[13] vssd1 vssd1 vccd1 vccd1 _14108_/Z sky130_fd_sc_hd__buf_12
Xrepeater136 peripheralBus_data[0] vssd1 vssd1 vccd1 vccd1 _13775_/Z sky130_fd_sc_hd__buf_12
X_08670_ _08670_/A vssd1 vssd1 vccd1 vccd1 _08670_/X sky130_fd_sc_hd__buf_2
XFILLER_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07621_ _07630_/A _07626_/B _07621_/C vssd1 vssd1 vccd1 vccd1 _07622_/A sky130_fd_sc_hd__or3_1
XFILLER_66_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09093__B_N input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07552_ _07552_/A vssd1 vssd1 vccd1 vccd1 _07552_/X sky130_fd_sc_hd__clkbuf_1
X_06503_ _06507_/A _06512_/B _06512_/C vssd1 vssd1 vccd1 vccd1 _06504_/A sky130_fd_sc_hd__or3_1
X_07483_ _07483_/A vssd1 vssd1 vccd1 vccd1 _07483_/X sky130_fd_sc_hd__clkbuf_1
X_06434_ _06434_/A vssd1 vssd1 vccd1 vccd1 _06434_/X sky130_fd_sc_hd__clkbuf_1
X_09222_ _09315_/C _09224_/C _09217_/X vssd1 vssd1 vccd1 vccd1 _09223_/B sky130_fd_sc_hd__o21ai_1
X_09153_ _10648_/A _09145_/X _09152_/X _09148_/X vssd1 vssd1 vccd1 vccd1 _12217_/D
+ sky130_fd_sc_hd__a211o_1
X_06365_ _06803_/A vssd1 vssd1 vccd1 vccd1 _07822_/B sky130_fd_sc_hd__clkbuf_2
X_08104_ _08104_/A vssd1 vssd1 vccd1 vccd1 _08104_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09084_ _09081_/X _09083_/X _09089_/S vssd1 vssd1 vccd1 vccd1 _10941_/C sky130_fd_sc_hd__mux2_1
X_06296_ _07045_/A vssd1 vssd1 vccd1 vccd1 _06308_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_107_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08035_ _08035_/A vssd1 vssd1 vccd1 vccd1 _11283_/B sky130_fd_sc_hd__buf_4
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09986_ _10107_/A _09997_/D _10030_/A vssd1 vssd1 vccd1 vccd1 _09993_/C sky130_fd_sc_hd__and3_1
X_08937_ _08926_/X _08935_/X _09043_/S vssd1 vssd1 vccd1 vccd1 _10939_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08868_ _08865_/X _08867_/X _08890_/S vssd1 vssd1 vccd1 vccd1 _10164_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09281__A _09281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07819_ _07819_/A vssd1 vssd1 vccd1 vccd1 _07819_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08799_ _12619_/Q vssd1 vssd1 vccd1 vccd1 _10863_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10830_ _10870_/B _10828_/A _10803_/X vssd1 vssd1 vccd1 vccd1 _10830_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10761_ _10863_/D _10806_/A _10760_/D _10863_/C vssd1 vssd1 vccd1 vccd1 _10762_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _12522_/CLK _12500_/D vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13480_ _13480_/A _07673_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
X_10692_ _10915_/A vssd1 vssd1 vccd1 vccd1 _10872_/A sky130_fd_sc_hd__clkbuf_4
X_12431_ _12617_/CLK _12431_/D vssd1 vssd1 vccd1 vccd1 _12431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08788__A1 _08782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ _12367_/CLK _12362_/D vssd1 vssd1 vccd1 vccd1 _13491_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11792__A0 _14063_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14101_ _14101_/A _08213_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[6] sky130_fd_sc_hd__ebufn_8
XFILLER_138_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11313_ _11325_/B vssd1 vssd1 vccd1 vccd1 _11323_/B sky130_fd_sc_hd__clkbuf_1
X_12293_ _12969_/CLK _12293_/D vssd1 vssd1 vccd1 vccd1 _13424_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10890__A _13775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ _11244_/A vssd1 vssd1 vccd1 vccd1 _12738_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09737__B1 _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14032_ _14032_/A _07864_/X vssd1 vssd1 vccd1 vccd1 _14064_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08360__A _08364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11175_ _13845_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11175_/X sky130_fd_sc_hd__or2_1
XFILLER_79_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10126_ _10130_/B _10130_/C _10126_/C _10126_/D vssd1 vssd1 vccd1 vccd1 _10127_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10057_ _10099_/D vssd1 vssd1 vccd1 vccd1 _10088_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09191__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13816_ _13816_/A _06789_/X vssd1 vssd1 vccd1 vccd1 _13976_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13747_ _13747_/A _06973_/X vssd1 vssd1 vccd1 vccd1 _14099_/Z sky130_fd_sc_hd__ebufn_8
X_10959_ _13811_/A _12665_/Q _10972_/S vssd1 vssd1 vccd1 vccd1 _10960_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13678_ _13678_/A _07148_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12629_ _12634_/CLK _12629_/D vssd1 vssd1 vccd1 vccd1 _12629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10035__B1 _09978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08626__S1 _08551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09840_ _13533_/A _12388_/Q _09843_/S vssd1 vssd1 vccd1 vccd1 _09841_/B sky130_fd_sc_hd__mux2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09771_ _13495_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09771_/X sky130_fd_sc_hd__or2_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07317__C _07993_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06983_ _08210_/A _06983_/B vssd1 vssd1 vccd1 vccd1 _10639_/A sky130_fd_sc_hd__or2_1
XFILLER_140_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08722_ _08719_/X _08721_/X _09941_/A vssd1 vssd1 vccd1 vccd1 _09399_/C sky130_fd_sc_hd__mux2_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08653_ _08555_/X _08561_/X _08558_/X _08565_/X _08695_/A _08652_/X vssd1 vssd1 vccd1
+ vccd1 _08653_/X sky130_fd_sc_hd__mux4_1
XANTENNA_repeater69_A peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07604_ _07923_/A vssd1 vssd1 vccd1 vccd1 _07661_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07333__B _07336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _13587_/A vssd1 vssd1 vccd1 vccd1 _08584_/X sky130_fd_sc_hd__buf_2
XFILLER_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07535_ _08197_/A vssd1 vssd1 vccd1 vccd1 _07545_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07466_ _07466_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07467_/A sky130_fd_sc_hd__or2_1
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09205_ _09205_/A vssd1 vssd1 vccd1 vccd1 _12229_/D sky130_fd_sc_hd__clkbuf_1
X_06417_ _06417_/A vssd1 vssd1 vccd1 vccd1 _06417_/X sky130_fd_sc_hd__clkbuf_1
X_07397_ _07397_/A vssd1 vssd1 vccd1 vccd1 _07397_/X sky130_fd_sc_hd__clkbuf_1
X_09136_ _09379_/A _09145_/A vssd1 vssd1 vccd1 vccd1 _09136_/X sky130_fd_sc_hd__or2_1
X_06348_ _06361_/A vssd1 vssd1 vccd1 vccd1 _06359_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09067_ _09067_/A vssd1 vssd1 vccd1 vccd1 _09067_/X sky130_fd_sc_hd__buf_2
XFILLER_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06279_ _11412_/A vssd1 vssd1 vccd1 vccd1 _06442_/A sky130_fd_sc_hd__buf_2
XFILLER_162_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08018_ _08166_/A vssd1 vssd1 vccd1 vccd1 _08072_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06412__B _06412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _10077_/A vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__buf_4
XFILLER_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09723__B _13554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12980_ _12980_/CLK _12980_/D vssd1 vssd1 vccd1 vccd1 _14105_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11931_ _14096_/Z _14032_/A _11940_/S vssd1 vssd1 vccd1 vccd1 _11932_/B sky130_fd_sc_hd__mux2_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _11869_/A _11862_/B vssd1 vssd1 vccd1 vccd1 _11863_/A sky130_fd_sc_hd__and2_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ _13601_/A _07362_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
X_10813_ _10813_/A vssd1 vssd1 vccd1 vccd1 _12629_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10885__A _10885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ _11799_/A _11793_/B vssd1 vssd1 vccd1 vccd1 _11794_/A sky130_fd_sc_hd__and2_1
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13532_ _13532_/A _07539_/X vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10744_ _10768_/A vssd1 vssd1 vccd1 vccd1 _10917_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_43_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ _13463_/A _07720_/X vssd1 vssd1 vccd1 vccd1 _13623_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10675_ _13721_/A _10684_/B vssd1 vssd1 vccd1 vccd1 _10675_/X sky130_fd_sc_hd__or2_1
X_12414_ _12414_/CLK _12414_/D vssd1 vssd1 vccd1 vccd1 _13590_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13394_ _13394_/A _08359_/X vssd1 vssd1 vccd1 vccd1 _14034_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_138_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12345_ _12349_/CLK _12345_/D vssd1 vssd1 vccd1 vccd1 _12345_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_repeater137_A peripheralBus_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09186__A _11189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12276_ _12289_/CLK _12276_/D vssd1 vssd1 vccd1 vccd1 _12276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14015_ _14015_/A _08071_/X vssd1 vssd1 vccd1 vccd1 _14079_/Z sky130_fd_sc_hd__ebufn_8
X_11227_ _11227_/A vssd1 vssd1 vccd1 vccd1 _12733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13260__416 vssd1 vssd1 vccd1 vccd1 _13260__416/HI _13931_/A sky130_fd_sc_hd__conb_1
X_11158_ _13839_/A _11168_/B vssd1 vssd1 vccd1 vccd1 _11158_/X sky130_fd_sc_hd__or2_1
XFILLER_110_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10109_ _10111_/B _10108_/B _10123_/A vssd1 vssd1 vccd1 vccd1 _10109_/Y sky130_fd_sc_hd__o21ai_1
X_11089_ _11095_/A _11089_/B vssd1 vssd1 vccd1 vccd1 _11090_/A sky130_fd_sc_hd__and2_1
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13301__457 vssd1 vssd1 vccd1 vccd1 _13301__457/HI _14022_/A sky130_fd_sc_hd__conb_1
XFILLER_91_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09110__A1 _09092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07320_ _09918_/B vssd1 vssd1 vccd1 vccd1 _09484_/B sky130_fd_sc_hd__buf_2
X_13154__310 vssd1 vssd1 vccd1 vccd1 _13154__310/HI _13727_/A sky130_fd_sc_hd__conb_1
X_07251_ _07251_/A vssd1 vssd1 vccd1 vccd1 _07251_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11403__B _13943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07182_ _07208_/A vssd1 vssd1 vccd1 vccd1 _07193_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09096__A input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07328__B _07336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09823_ _09843_/S vssd1 vssd1 vccd1 vccd1 _09837_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10731__A1 _10285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09754_ _13490_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09754_/X sky130_fd_sc_hd__or2_1
XFILLER_86_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06966_ _06966_/A vssd1 vssd1 vccd1 vccd1 _06966_/X sky130_fd_sc_hd__clkbuf_1
X_08705_ _12462_/Q vssd1 vssd1 vccd1 vccd1 _10148_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__07344__A _07371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09685_ _13495_/A _12349_/Q _09685_/S vssd1 vssd1 vccd1 vccd1 _09686_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06897_ _06897_/A vssd1 vssd1 vccd1 vccd1 _06897_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_93_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _12400_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _12441_/Q vssd1 vssd1 vccd1 vccd1 _10052_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08567_ _12445_/Q _12446_/Q _12447_/Q _12448_/Q _08559_/X _08560_/X vssd1 vssd1 vccd1
+ vccd1 _08567_/X sky130_fd_sc_hd__mux4_2
XFILLER_154_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07518_ _07518_/A vssd1 vssd1 vccd1 vccd1 _07518_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08498_ _08493_/X _08497_/X _08498_/S vssd1 vssd1 vccd1 vccd1 _11707_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07449_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07459_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10460_ _13688_/A _12543_/Q _10473_/S vssd1 vssd1 vccd1 vccd1 _10461_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ peripheralBus_data[15] vssd1 vssd1 vccd1 vccd1 _10552_/A sky130_fd_sc_hd__clkbuf_4
X_10391_ _09753_/X _10379_/X _10390_/X _10383_/X vssd1 vssd1 vccd1 vccd1 _12521_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09718__B _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ _12130_/A vssd1 vssd1 vccd1 vccd1 _12960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ _12088_/A vssd1 vssd1 vccd1 vccd1 _12061_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ _12668_/Q _13942_/A vssd1 vssd1 vccd1 vccd1 _11016_/A sky130_fd_sc_hd__xor2_1
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12963_ _12981_/CLK _12963_/D vssd1 vssd1 vccd1 vccd1 _12963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_84_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _12470_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_161_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11914_ _12899_/Q _13371_/A vssd1 vssd1 vccd1 vccd1 _11915_/D sky130_fd_sc_hd__xor2_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12894_ _12918_/CLK _12894_/D vssd1 vssd1 vccd1 vccd1 _12894_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11845_ _11845_/A vssd1 vssd1 vccd1 vccd1 _12886_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08526__S0 _09140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _12856_/Q _13361_/A vssd1 vssd1 vccd1 vccd1 _11780_/A sky130_fd_sc_hd__xor2_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13515_ _13515_/A _07581_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
X_10727_ _10408_/X _10690_/X _10726_/X _10711_/X vssd1 vssd1 vccd1 vccd1 _12610_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13446_ _13446_/A _07762_/X vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10658_ _10394_/X _10655_/X _10657_/X _10650_/X vssd1 vssd1 vccd1 vccd1 _12589_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13377_ _13377_/A _08320_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
X_10589_ _13720_/A _12576_/Q _10601_/S vssd1 vssd1 vccd1 vccd1 _10590_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12328_ _12331_/CLK _12328_/D vssd1 vssd1 vccd1 vccd1 _13458_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12054__B _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12259_ _12264_/CLK _12259_/D vssd1 vssd1 vccd1 vccd1 _12259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09644__A _11189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06820_ _07248_/A vssd1 vssd1 vccd1 vccd1 _06967_/A sky130_fd_sc_hd__buf_2
XFILLER_96_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06751_ _06760_/A _06751_/B _06751_/C vssd1 vssd1 vccd1 vccd1 _06752_/A sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_75_clk _12555_/CLK vssd1 vssd1 vccd1 vccd1 _12492_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09470_ _12288_/Q _13564_/A vssd1 vssd1 vccd1 vccd1 _09473_/B sky130_fd_sc_hd__xnor2_1
X_06682_ _06686_/A _06692_/B _06692_/C vssd1 vssd1 vccd1 vccd1 _06683_/A sky130_fd_sc_hd__or3_1
XFILLER_64_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08421_ _09258_/D _12239_/Q _12240_/Q _12241_/Q _08373_/X _08374_/X vssd1 vssd1 vccd1
+ vccd1 _08421_/X sky130_fd_sc_hd__mux4_2
XFILLER_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08352_ _08358_/A _08358_/B _08360_/C vssd1 vssd1 vccd1 vccd1 _08353_/A sky130_fd_sc_hd__or3_1
XFILLER_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11977__A0 _14110_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07303_ _07307_/A _07303_/B _07314_/C vssd1 vssd1 vccd1 vccd1 _07304_/A sky130_fd_sc_hd__or3_1
XFILLER_165_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08283_ _08288_/A _08285_/B vssd1 vssd1 vccd1 vccd1 _08284_/A sky130_fd_sc_hd__or2_1
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09819__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07234_ _07739_/A _07947_/B _07234_/C vssd1 vssd1 vccd1 vccd1 _07235_/A sky130_fd_sc_hd__or3_1
X_07165_ _07205_/A vssd1 vssd1 vccd1 vccd1 _07177_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07339__A _07393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07096_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07108_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09806_ _09843_/S vssd1 vssd1 vccd1 vccd1 _09820_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07998_ _07998_/A vssd1 vssd1 vccd1 vccd1 _07998_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09737_ _09714_/Y _09720_/X _09736_/Y _13568_/A vssd1 vssd1 vccd1 vccd1 _09738_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_101_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06949_ _06949_/A vssd1 vssd1 vccd1 vccd1 _06949_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_66_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _12647_/CLK sky130_fd_sc_hd__clkbuf_16
X_09668_ _13490_/A _12344_/Q _09738_/B vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__mux2_1
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _12451_/Q _10101_/A _10111_/C _12454_/Q _08553_/X _08554_/X vssd1 vssd1 vccd1
+ vccd1 _08619_/X sky130_fd_sc_hd__mux4_2
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12209__A1 _11189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09599_ _12320_/Q _13563_/A vssd1 vssd1 vccd1 vccd1 _09602_/B sky130_fd_sc_hd__xor2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11639_/A _11640_/A _11641_/A _11630_/D vssd1 vssd1 vccd1 vccd1 _11633_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11968__A0 _14107_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06418__A _06442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ _11561_/A vssd1 vssd1 vccd1 vccd1 _12819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10512_ _11285_/B _10512_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _10553_/B sky130_fd_sc_hd__nor3_2
X_11492_ _14009_/Z _11494_/B vssd1 vssd1 vccd1 vccd1 _11492_/X sky130_fd_sc_hd__or2_1
XFILLER_109_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10443_ _13683_/A _12538_/Q _10456_/S vssd1 vssd1 vccd1 vccd1 _10444_/B sky130_fd_sc_hd__mux2_1
XFILLER_136_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11196__A1 _11064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08352__B _08358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10374_ _10351_/Y _10357_/X _10373_/Y _13761_/A vssd1 vssd1 vccd1 vccd1 _10375_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12113_ _12113_/A vssd1 vssd1 vccd1 vccd1 _12955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12044_ _12934_/Q _13373_/A vssd1 vssd1 vccd1 vccd1 _12045_/D sky130_fd_sc_hd__xor2_1
XFILLER_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13995_ _13995_/A _06298_/X vssd1 vssd1 vccd1 vccd1 _13995_/Z sky130_fd_sc_hd__ebufn_8
Xclkbuf_leaf_57_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _12842_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12946_ _12946_/CLK _12946_/D vssd1 vssd1 vccd1 vccd1 _14072_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output29_A _13787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ _12904_/CLK _12877_/D vssd1 vssd1 vccd1 vccd1 _14005_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11234__A _11254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _11834_/A _11828_/B vssd1 vssd1 vccd1 vccd1 _11829_/A sky130_fd_sc_hd__and2_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12049__B _13371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11759_ _11801_/A vssd1 vssd1 vccd1 vccd1 _11799_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13429_ _13429_/A _07807_/X vssd1 vssd1 vccd1 vccd1 _14037_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266__422 vssd1 vssd1 vccd1 vccd1 _13266__422/HI _13957_/A sky130_fd_sc_hd__conb_1
XFILLER_127_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08970_ _12817_/Q _11562_/C _12819_/Q _12820_/Q _08967_/X _08968_/X vssd1 vssd1 vccd1
+ vccd1 _08970_/X sky130_fd_sc_hd__mux4_2
XANTENNA__06998__A _07979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07921_ _07921_/A _07931_/B _07931_/C vssd1 vssd1 vccd1 vccd1 _07922_/A sky130_fd_sc_hd__or3_1
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13307__463 vssd1 vssd1 vccd1 vccd1 _13307__463/HI _14028_/A sky130_fd_sc_hd__conb_1
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07852_ _07962_/A _07854_/B _07852_/C vssd1 vssd1 vccd1 vccd1 _07853_/A sky130_fd_sc_hd__or3_1
XFILLER_96_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06803_ _06803_/A vssd1 vssd1 vccd1 vccd1 _07857_/A sky130_fd_sc_hd__buf_2
XANTENNA__11128__B _13948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 peripheralBus_address[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
X_07783_ _07783_/A vssd1 vssd1 vccd1 vccd1 _07783_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _12682_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09522_ _09634_/A vssd1 vssd1 vccd1 vccd1 _09522_/X sky130_fd_sc_hd__clkbuf_2
X_06734_ _06734_/A vssd1 vssd1 vccd1 vccd1 _06734_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09453_ _09453_/A vssd1 vssd1 vccd1 vccd1 _12289_/D sky130_fd_sc_hd__clkbuf_1
X_06665_ _06665_/A vssd1 vssd1 vccd1 vccd1 _06665_/X sky130_fd_sc_hd__clkbuf_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08404_ _13392_/A vssd1 vssd1 vccd1 vccd1 _08404_/X sky130_fd_sc_hd__buf_2
XFILLER_40_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09384_ _09388_/C _09384_/B vssd1 vssd1 vccd1 vccd1 _12271_/D sky130_fd_sc_hd__nor2_1
XFILLER_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06596_ _06596_/A vssd1 vssd1 vccd1 vccd1 _06596_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08335_ _08335_/A vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07060__C _07969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08266_ _08266_/A vssd1 vssd1 vccd1 vccd1 _08276_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__07995__C _08180_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07217_ _07217_/A vssd1 vssd1 vccd1 vccd1 _07217_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11178__A1 _10662_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ _08197_/A vssd1 vssd1 vccd1 vccd1 _08208_/B sky130_fd_sc_hd__clkbuf_2
X_07148_ _07148_/A vssd1 vssd1 vccd1 vccd1 _07148_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09240__B1 _09206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07079_ _07079_/A _07091_/B _07088_/C vssd1 vssd1 vccd1 vccd1 _07080_/A sky130_fd_sc_hd__or3_1
XFILLER_10_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10090_ _10098_/A _10083_/B _10097_/A vssd1 vssd1 vccd1 vccd1 _10091_/C sky130_fd_sc_hd__a21o_1
XFILLER_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _12780_/CLK sky130_fd_sc_hd__clkbuf_16
X_12800_ _12800_/CLK _12800_/D vssd1 vssd1 vccd1 vccd1 _13974_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09731__B _13551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13780_ _13780_/A _06891_/X vssd1 vssd1 vccd1 vccd1 _14100_/Z sky130_fd_sc_hd__ebufn_8
X_10992_ _10992_/A vssd1 vssd1 vccd1 vccd1 _12674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12731_ _12753_/CLK _12731_/D vssd1 vssd1 vccd1 vccd1 _12731_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08347__B _08349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13100__256 vssd1 vssd1 vccd1 vccd1 _13100__256/HI _13609_/A sky130_fd_sc_hd__conb_1
X_12662_ _12687_/CLK _12662_/D vssd1 vssd1 vccd1 vccd1 _12662_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11641_/B vssd1 vssd1 vccd1 vccd1 _11630_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _12593_/CLK _12593_/D vssd1 vssd1 vccd1 vccd1 _13720_/A sky130_fd_sc_hd__dfxtp_1
X_11544_ _11627_/C _11627_/D _11547_/D vssd1 vssd1 vccd1 vccd1 _11563_/A sky130_fd_sc_hd__and3_1
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11475_ _14099_/Z _09057_/X _11489_/S vssd1 vssd1 vccd1 vccd1 _11476_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11169__A1 _10652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10426_ _09120_/X _10409_/A _10423_/X _10425_/X vssd1 vssd1 vccd1 vccd1 _12533_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10916__A1 _10885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09782__A1 _09186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10357_ _10352_/Y _10353_/X _10354_/X _10355_/Y _10356_/Y vssd1 vssd1 vccd1 vccd1
+ _10357_/X sky130_fd_sc_hd__o221a_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10288_ _11064_/A vssd1 vssd1 vccd1 vccd1 _10288_/X sky130_fd_sc_hd__buf_4
XFILLER_25_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12027_ _12030_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _12028_/A sky130_fd_sc_hd__and2_1
XFILLER_66_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09922__A _13583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09298__B1 _09236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13978_ _13978_/A _06345_/X vssd1 vssd1 vccd1 vccd1 _13978_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_81_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12929_ _12929_/CLK _12929_/D vssd1 vssd1 vccd1 vccd1 _12929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10852__B1 _10803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06450_ _06450_/A vssd1 vssd1 vccd1 vccd1 _06450_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06381_ _06391_/A _08349_/A vssd1 vssd1 vccd1 vccd1 _06382_/A sky130_fd_sc_hd__or2_1
XFILLER_159_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08120_ _08122_/A _08184_/B _08131_/C vssd1 vssd1 vccd1 vccd1 _08121_/A sky130_fd_sc_hd__or3_2
X_08051_ _08051_/A vssd1 vssd1 vccd1 vccd1 _08051_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07002_ _07002_/A vssd1 vssd1 vccd1 vccd1 _07002_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08953_ _13971_/A vssd1 vssd1 vccd1 vccd1 _08953_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09525__A1 _13437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ _07904_/A vssd1 vssd1 vccd1 vccd1 _07904_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07336__B _07336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ _08747_/X _08754_/X _08752_/X _08756_/X _08837_/X _08838_/X vssd1 vssd1 vccd1
+ vccd1 _08884_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07835_ _07843_/A _07840_/B _08180_/C vssd1 vssd1 vccd1 vccd1 _07836_/A sky130_fd_sc_hd__or3_1
XFILLER_96_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07766_ _07769_/A _07766_/B _07774_/C vssd1 vssd1 vccd1 vccd1 _07767_/A sky130_fd_sc_hd__or3_1
XFILLER_72_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09505_ _13429_/A _09500_/X _09504_/X _09496_/X vssd1 vssd1 vccd1 vccd1 _12298_/D
+ sky130_fd_sc_hd__o211a_1
X_06717_ _06733_/A _06719_/B _06719_/C vssd1 vssd1 vccd1 vccd1 _06718_/A sky130_fd_sc_hd__or3_1
XFILLER_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07697_ _07697_/A vssd1 vssd1 vccd1 vccd1 _07697_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09436_ _09439_/A _09436_/B vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__and2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06648_ _06675_/A vssd1 vssd1 vccd1 vccd1 _06659_/A sky130_fd_sc_hd__clkbuf_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09367_ _09368_/A _09364_/B _09206_/X vssd1 vssd1 vccd1 vccd1 _09369_/A sky130_fd_sc_hd__o21ai_1
X_06579_ _06633_/A vssd1 vssd1 vccd1 vccd1 _06589_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08318_ _08318_/A vssd1 vssd1 vccd1 vccd1 _08318_/X sky130_fd_sc_hd__clkbuf_1
X_09298_ _09329_/C _09300_/C _09236_/X vssd1 vssd1 vccd1 vccd1 _09299_/B sky130_fd_sc_hd__o21ai_1
XFILLER_165_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08249_ _08249_/A vssd1 vssd1 vccd1 vccd1 _08249_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11260_ _12728_/Q _13936_/A vssd1 vssd1 vccd1 vccd1 _11260_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10211_ _13627_/A _12480_/Q _10214_/S vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__mux2_1
XFILLER_106_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11191_ _11189_/X _11185_/X _11190_/X _11180_/X vssd1 vssd1 vccd1 vccd1 _12722_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09726__B _13553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10142_ _10148_/B _10142_/B vssd1 vssd1 vccd1 vccd1 _10145_/B sky130_fd_sc_hd__and2_1
XFILLER_121_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10073_ _10099_/B vssd1 vssd1 vccd1 vccd1 _10073_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13901_ _13901_/A _06555_/X vssd1 vssd1 vccd1 vccd1 _14125_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_153_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13832_ _13832_/A _06745_/X vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__09461__B _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08358__A _08358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13763_ _13763_/A _06935_/X vssd1 vssd1 vccd1 vccd1 _13987_/Z sky130_fd_sc_hd__ebufn_8
X_10975_ _10996_/S vssd1 vssd1 vccd1 vccd1 _10990_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_43_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12714_ _12722_/CLK _12714_/D vssd1 vssd1 vccd1 vccd1 _13842_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13694_ _13694_/A _07109_/X vssd1 vssd1 vccd1 vccd1 _14078_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12645_ _12646_/CLK _12645_/D vssd1 vssd1 vccd1 vccd1 _12645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09189__A _13403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08093__A _09125_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ _12800_/CLK _12576_/D vssd1 vssd1 vccd1 vccd1 _12576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11527_ _12812_/Q vssd1 vssd1 vccd1 vccd1 _11625_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11458_ _11460_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _11459_/A sky130_fd_sc_hd__and2_1
XANTENNA__09755__A1 _09753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ _10409_/A vssd1 vssd1 vccd1 vccd1 _10409_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11389_ _12771_/Q _13946_/A vssd1 vssd1 vccd1 vccd1 _11389_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07437__A _08131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12062__B _12062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater104 peripheralBus_data[21] vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__buf_12
Xrepeater115 _14112_/Z vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__buf_12
Xrepeater126 peripheralBus_data[13] vssd1 vssd1 vccd1 vccd1 _14012_/Z sky130_fd_sc_hd__buf_12
Xrepeater137 peripheralBus_data[0] vssd1 vssd1 vccd1 vccd1 _14063_/Z sky130_fd_sc_hd__buf_12
XFILLER_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07620_ _07620_/A vssd1 vssd1 vccd1 vccd1 _07620_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07551_ _07558_/A _07558_/B _07551_/C vssd1 vssd1 vccd1 vccd1 _07552_/A sky130_fd_sc_hd__or3_1
X_06502_ _08276_/B vssd1 vssd1 vccd1 vccd1 _06512_/C sky130_fd_sc_hd__clkbuf_1
X_07482_ _08089_/A _07484_/B vssd1 vssd1 vccd1 vccd1 _07483_/A sky130_fd_sc_hd__or2_1
XFILLER_22_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09221_ _09315_/C _09224_/C vssd1 vssd1 vccd1 vccd1 _09223_/A sky130_fd_sc_hd__and2_1
X_06433_ _06440_/A _06437_/B vssd1 vssd1 vccd1 vccd1 _06434_/A sky130_fd_sc_hd__or2_1
X_09152_ _09152_/A _09152_/B vssd1 vssd1 vccd1 vccd1 _09152_/X sky130_fd_sc_hd__and2_1
X_06364_ _11457_/B vssd1 vssd1 vccd1 vccd1 _06803_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__06516__A _07507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08103_ _08110_/A _08103_/B _08110_/C vssd1 vssd1 vccd1 vccd1 _08104_/A sky130_fd_sc_hd__or3_1
XANTENNA__11141__B _13947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ _08980_/X _09026_/X _09052_/X _09082_/X _09056_/X _09057_/X vssd1 vssd1 vccd1
+ vccd1 _09083_/X sky130_fd_sc_hd__mux4_1
X_06295_ _08266_/A vssd1 vssd1 vccd1 vccd1 _07045_/A sky130_fd_sc_hd__buf_2
XANTENNA__10038__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ _08034_/A vssd1 vssd1 vccd1 vccd1 _08034_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09746__A1 _09124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_51_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09985_ _09985_/A vssd1 vssd1 vccd1 vccd1 _12424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12986__142 vssd1 vssd1 vccd1 vccd1 _12986__142/HI _13383_/A sky130_fd_sc_hd__conb_1
X_08936_ _13972_/A vssd1 vssd1 vccd1 vccd1 _09043_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08867_ _08773_/X _08774_/X _08840_/X _08866_/X _08826_/X _08859_/X vssd1 vssd1 vccd1
+ vccd1 _08867_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_66_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _07868_/A _07820_/B _08110_/C vssd1 vssd1 vccd1 vccd1 _07819_/A sky130_fd_sc_hd__or3_1
XFILLER_45_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08178__A _08358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08798_ _10163_/C vssd1 vssd1 vccd1 vccd1 _13745_/A sky130_fd_sc_hd__buf_4
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07082__A _07533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07749_ _07749_/A vssd1 vssd1 vccd1 vccd1 _07749_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09682__A0 _13494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ _10863_/C _10863_/D _10806_/A _10760_/D vssd1 vssd1 vccd1 vccd1 _10767_/C
+ sky130_fd_sc_hd__and4_1
X_09419_ _09422_/A _09419_/B vssd1 vssd1 vccd1 vccd1 _09420_/A sky130_fd_sc_hd__and2_1
XANTENNA__10292__A1 _09116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ _13775_/A vssd1 vssd1 vccd1 vccd1 _10915_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171__327 vssd1 vssd1 vccd1 vccd1 _13171__327/HI _13764_/A sky130_fd_sc_hd__conb_1
XFILLER_139_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12430_ _12617_/CLK _12430_/D vssd1 vssd1 vccd1 vccd1 _12430_/Q sky130_fd_sc_hd__dfxtp_1
X_12361_ _12367_/CLK _12361_/D vssd1 vssd1 vccd1 vccd1 _13490_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14100_ _14100_/A _08209_/X vssd1 vssd1 vccd1 vccd1 _14100_/Z sky130_fd_sc_hd__ebufn_8
X_11312_ _11312_/A vssd1 vssd1 vccd1 vccd1 _11312_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13212__368 vssd1 vssd1 vccd1 vccd1 _13212__368/HI _13835_/A sky130_fd_sc_hd__conb_1
XFILLER_165_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12292_ _12295_/CLK _12292_/D vssd1 vssd1 vccd1 vccd1 _13423_/A sky130_fd_sc_hd__dfxtp_1
X_14031_ _14031_/A _08185_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[0] sky130_fd_sc_hd__ebufn_8
XFILLER_141_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11243_ _11255_/A _11243_/B vssd1 vssd1 vccd1 vccd1 _11244_/A sky130_fd_sc_hd__and2_1
XFILLER_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08360__B _08364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_clk_A _12881_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ _11170_/X _11171_/X _11173_/X _11166_/X vssd1 vssd1 vccd1 vccd1 _12716_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13065__221 vssd1 vssd1 vccd1 vccd1 _13065__221/HI _13540_/A sky130_fd_sc_hd__conb_1
X_10125_ _10130_/C _10130_/D _10126_/D _10130_/B vssd1 vssd1 vccd1 vccd1 _10127_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10056_ _10056_/A vssd1 vssd1 vccd1 vccd1 _12442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13106__262 vssd1 vssd1 vccd1 vccd1 _13106__262/HI _13631_/A sky130_fd_sc_hd__conb_1
XANTENNA__11507__A _11634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13815_ _13815_/A _06792_/X vssd1 vssd1 vccd1 vccd1 _14007_/Z sky130_fd_sc_hd__ebufn_8
X_13746_ _13746_/A _06976_/X vssd1 vssd1 vccd1 vccd1 _14098_/Z sky130_fd_sc_hd__ebufn_8
X_10958_ _10996_/S vssd1 vssd1 vccd1 vccd1 _10972_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11480__A0 _13973_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13677_ _13677_/A _07153_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
X_10889_ _10908_/B vssd1 vssd1 vccd1 vccd1 _10897_/C sky130_fd_sc_hd__clkbuf_1
X_12628_ _12646_/CLK _12628_/D vssd1 vssd1 vccd1 vccd1 _12628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12559_ _12565_/CLK _12559_/D vssd1 vssd1 vccd1 vccd1 _13687_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09647__A _09846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _10665_/A vssd1 vssd1 vccd1 vccd1 _09770_/X sky130_fd_sc_hd__buf_6
X_06982_ _07033_/A vssd1 vssd1 vccd1 vccd1 _06995_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _08619_/X _08666_/X _08690_/X _08720_/X _08694_/X _08695_/X vssd1 vssd1 vccd1
+ vccd1 _08721_/X sky130_fd_sc_hd__mux4_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08652_ _08670_/A vssd1 vssd1 vccd1 vccd1 _08652_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07603_ _07603_/A vssd1 vssd1 vccd1 vccd1 _07923_/A sky130_fd_sc_hd__buf_4
XANTENNA__11136__B _13941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ _13586_/A vssd1 vssd1 vccd1 vccd1 _08583_/X sky130_fd_sc_hd__buf_2
XANTENNA__07333__C _07739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07534_ _07590_/A vssd1 vssd1 vccd1 vccd1 _07545_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11471__A0 _14066_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07465_ _07465_/A vssd1 vssd1 vccd1 vccd1 _07465_/X sky130_fd_sc_hd__clkbuf_1
X_09204_ _09201_/X _09204_/B _09372_/B vssd1 vssd1 vccd1 vccd1 _09205_/A sky130_fd_sc_hd__and3b_1
XFILLER_10_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06416_ _06416_/A _06425_/B vssd1 vssd1 vccd1 vccd1 _06417_/A sky130_fd_sc_hd__or2_1
XFILLER_148_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07396_ _07396_/A _07404_/B _07401_/C vssd1 vssd1 vccd1 vccd1 _07397_/A sky130_fd_sc_hd__or3_1
X_09135_ _09161_/A vssd1 vssd1 vccd1 vccd1 _09145_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06347_ _06347_/A vssd1 vssd1 vccd1 vccd1 _06347_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09066_ _08923_/X _08930_/X _08931_/X _08932_/X _08994_/X _08996_/X vssd1 vssd1 vccd1
+ vccd1 _09066_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06278_ _11457_/B vssd1 vssd1 vccd1 vccd1 _11412_/A sky130_fd_sc_hd__clkbuf_4
X_08017_ _08017_/A vssd1 vssd1 vccd1 vccd1 _08017_/X sky130_fd_sc_hd__clkbuf_1
X_13049__205 vssd1 vssd1 vccd1 vccd1 _13049__205/HI _13508_/A sky130_fd_sc_hd__conb_1
XANTENNA__08180__B _08180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09968_ _09977_/A vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08919_ _13969_/A vssd1 vssd1 vccd1 vccd1 _08919_/X sky130_fd_sc_hd__clkbuf_4
X_09899_ _09770_/X _09888_/X _09898_/X _09892_/X vssd1 vssd1 vccd1 vccd1 _12399_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11327__A _11363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ _11998_/A vssd1 vssd1 vccd1 vccd1 _11945_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11861_ _12891_/Q _14035_/A _11861_/S vssd1 vssd1 vccd1 vccd1 _11862_/B sky130_fd_sc_hd__mux2_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _13600_/A _07365_/X vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10812_ _10878_/B _10812_/B _10812_/C vssd1 vssd1 vccd1 vccd1 _10813_/A sky130_fd_sc_hd__and3b_1
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11792_ _14063_/Z _13999_/A _11805_/S vssd1 vssd1 vccd1 vccd1 _11793_/B sky130_fd_sc_hd__mux2_1
XFILLER_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13531_ _13531_/A _07542_/X vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__07540__A _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10743_ _10885_/A _10806_/D _10806_/C vssd1 vssd1 vccd1 vccd1 _10745_/B sky130_fd_sc_hd__a21o_1
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _13462_/A _07723_/X vssd1 vssd1 vccd1 vccd1 _14102_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10674_ _10686_/B vssd1 vssd1 vccd1 vccd1 _10684_/B sky130_fd_sc_hd__clkbuf_2
X_12413_ _12414_/CLK _12413_/D vssd1 vssd1 vccd1 vccd1 _13589_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13393_ _13393_/A _08357_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[2] sky130_fd_sc_hd__ebufn_8
XFILLER_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12344_ _12349_/CLK _12344_/D vssd1 vssd1 vccd1 vccd1 _12344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12275_ _12301_/CLK _12275_/D vssd1 vssd1 vccd1 vccd1 _12275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14014_ _14014_/A _08127_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
XFILLER_107_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11226_ _11239_/A _11226_/B vssd1 vssd1 vccd1 vccd1 _11227_/A sky130_fd_sc_hd__and2_1
XFILLER_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12190__A1 _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11157_ _11199_/B vssd1 vssd1 vccd1 vccd1 _11168_/B sky130_fd_sc_hd__clkbuf_1
X_10108_ _10108_/A _10108_/B _09987_/X vssd1 vssd1 vccd1 vccd1 _12453_/D sky130_fd_sc_hd__nor3b_1
XANTENNA_output59_A _13760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11088_ _13843_/A _12698_/Q _11101_/S vssd1 vssd1 vccd1 vccd1 _11089_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10039_ _09982_/A _10097_/C _10053_/B _10097_/B vssd1 vssd1 vccd1 vccd1 _10040_/B
+ sky130_fd_sc_hd__a31o_1
X_13340__496 vssd1 vssd1 vccd1 vccd1 _13340__496/HI _14093_/A sky130_fd_sc_hd__conb_1
XFILLER_36_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13729_ _13729_/A _07018_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[18] sky130_fd_sc_hd__ebufn_8
XFILLER_31_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07250_ _07253_/A _07250_/B _07260_/C vssd1 vssd1 vccd1 vccd1 _07251_/A sky130_fd_sc_hd__or3_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07181_ _07181_/A vssd1 vssd1 vccd1 vccd1 _07181_/X sky130_fd_sc_hd__clkbuf_1
X_13234__390 vssd1 vssd1 vccd1 vccd1 _13234__390/HI _13889_/A sky130_fd_sc_hd__conb_1
XFILLER_145_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09096__B _09096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07328__C _07739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12181__A1 _11153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09822_ _09822_/A vssd1 vssd1 vccd1 vccd1 _12382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10731__A2 _10703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater81_A _14126_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ _10648_/A vssd1 vssd1 vccd1 vccd1 _09753_/X sky130_fd_sc_hd__buf_6
XFILLER_101_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06965_ _06972_/A _06965_/B vssd1 vssd1 vccd1 vccd1 _06966_/A sky130_fd_sc_hd__or2_1
XFILLER_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08704_ _08561_/X _08565_/X _08566_/X _08567_/X _08632_/X _08634_/X vssd1 vssd1 vccd1
+ vccd1 _08704_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09684_ _09684_/A vssd1 vssd1 vccd1 vccd1 _12348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06896_ _07328_/A _06898_/B _06898_/C vssd1 vssd1 vccd1 vccd1 _06897_/A sky130_fd_sc_hd__or3_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ _08624_/X _08626_/X _08628_/X _08631_/X _08632_/X _08634_/X vssd1 vssd1 vccd1
+ vccd1 _08635_/X sky130_fd_sc_hd__mux4_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13362__A _13362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08566_ _12441_/Q _12442_/Q _12443_/Q _12444_/Q _08559_/X _08560_/X vssd1 vssd1 vccd1
+ vccd1 _08566_/X sky130_fd_sc_hd__mux4_2
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07517_ _07517_/A _07517_/B _07524_/C vssd1 vssd1 vccd1 vccd1 _07518_/A sky130_fd_sc_hd__or3_1
X_08497_ _08389_/X _08390_/X _08469_/X _08496_/X _08492_/X _08424_/X vssd1 vssd1 vccd1
+ vccd1 _08497_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07448_ _07448_/A vssd1 vssd1 vccd1 vccd1 _07448_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07379_ _07393_/A vssd1 vssd1 vccd1 vccd1 _07391_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_108_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09118_ _09116_/X _09100_/X _09117_/X _09109_/X vssd1 vssd1 vccd1 vccd1 _12212_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10390_ _13650_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10390_/X sky130_fd_sc_hd__or2_1
XFILLER_129_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09049_ _11384_/B vssd1 vssd1 vccd1 vccd1 _13944_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_163_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13283__439 vssd1 vssd1 vccd1 vccd1 _13283__439/HI _13988_/A sky130_fd_sc_hd__conb_1
X_12060_ _12060_/A _12062_/B _12059_/Y vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__or3b_2
X_11011_ _11011_/A _11011_/B _11011_/C _11011_/D vssd1 vssd1 vccd1 vccd1 _11022_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_145_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09734__B _13555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12160__B _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12962_ _12962_/CLK _12962_/D vssd1 vssd1 vccd1 vccd1 _12962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input10_A peripheralBus_address[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09750__A _10645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _12894_/Q _13366_/A vssd1 vssd1 vccd1 vccd1 _11915_/C sky130_fd_sc_hd__xor2_1
XFILLER_73_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _12895_/CLK _12893_/D vssd1 vssd1 vccd1 vccd1 _12893_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13177__333 vssd1 vssd1 vccd1 vccd1 _13177__333/HI _13770_/A sky130_fd_sc_hd__conb_1
X_11844_ _11852_/A _11844_/B vssd1 vssd1 vccd1 vccd1 _11845_/A sky130_fd_sc_hd__and2_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08526__S1 _09146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11775_/A _11775_/B _11775_/C _11775_/D vssd1 vssd1 vccd1 vccd1 _11786_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _13514_/A _07584_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
X_10726_ _13785_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10726_/X sky130_fd_sc_hd__or2_1
XFILLER_159_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13218__374 vssd1 vssd1 vccd1 vccd1 _13218__374/HI _13857_/A sky130_fd_sc_hd__conb_1
XFILLER_158_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13445_ _13445_/A _07765_/X vssd1 vssd1 vccd1 vccd1 _13765_/Z sky130_fd_sc_hd__ebufn_8
X_10657_ _13716_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10657_/X sky130_fd_sc_hd__or2_1
XFILLER_70_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09197__A _09281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13376_ _13376_/A _08318_/X vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__ebufn_8
X_10588_ _10608_/S vssd1 vssd1 vccd1 vccd1 _10601_/S sky130_fd_sc_hd__clkbuf_2
X_12327_ _12331_/CLK _12327_/D vssd1 vssd1 vccd1 vccd1 _13457_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12258_ _12258_/CLK _12258_/D vssd1 vssd1 vccd1 vccd1 _12258_/Q sky130_fd_sc_hd__dfxtp_1
X_11209_ _11209_/A vssd1 vssd1 vccd1 vccd1 _12728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189_ _14098_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12189_/X sky130_fd_sc_hd__or2_1
XFILLER_110_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06750_ _06750_/A vssd1 vssd1 vccd1 vccd1 _06750_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06681_ _06722_/A vssd1 vssd1 vccd1 vccd1 _06692_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_52_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ _12234_/Q _12235_/Q _12236_/Q _12237_/Q _08373_/X _08374_/X vssd1 vssd1 vccd1
+ vccd1 _08420_/X sky130_fd_sc_hd__mux4_2
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08351_ _08351_/A vssd1 vssd1 vccd1 vccd1 _08360_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07302_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07314_/C sky130_fd_sc_hd__clkbuf_1
X_08282_ _08282_/A vssd1 vssd1 vccd1 vccd1 _08282_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07233_ _08177_/A vssd1 vssd1 vccd1 vccd1 _07739_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07164_ _07164_/A vssd1 vssd1 vccd1 vccd1 _07164_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10401__A1 _09763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07095_ _07095_/A vssd1 vssd1 vccd1 vccd1 _07095_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13011__167 vssd1 vssd1 vccd1 vccd1 _13011__167/HI _13422_/A sky130_fd_sc_hd__conb_1
XFILLER_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10480__S _10480_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09805_ _09805_/A vssd1 vssd1 vccd1 vccd1 _12377_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input2_A peripheralBus_address[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07997_ _07997_/A _08005_/B _08002_/C vssd1 vssd1 vccd1 vccd1 _07998_/A sky130_fd_sc_hd__or3_1
XFILLER_86_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09736_ _09736_/A _09736_/B _09736_/C vssd1 vssd1 vccd1 vccd1 _09736_/Y sky130_fd_sc_hd__nor3_1
X_06948_ _06948_/A _06953_/B vssd1 vssd1 vccd1 vccd1 _06949_/A sky130_fd_sc_hd__or2_1
XFILLER_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09667_ _09667_/A vssd1 vssd1 vccd1 vccd1 _12343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06879_ _06879_/A vssd1 vssd1 vccd1 vccd1 _06890_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08618_ _12453_/Q vssd1 vssd1 vccd1 vccd1 _10111_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09598_ _12310_/Q _13553_/A vssd1 vssd1 vccd1 vccd1 _09602_/A sky130_fd_sc_hd__xor2_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08186__A _08186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07090__A _07090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08549_ _08708_/A vssd1 vssd1 vccd1 vccd1 _08549_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ _11565_/C _11604_/B _11560_/C vssd1 vssd1 vccd1 vccd1 _11561_/A sky130_fd_sc_hd__and3b_1
XFILLER_23_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ _10538_/A vssd1 vssd1 vccd1 vccd1 _10511_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09729__B _13558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ _11491_/A vssd1 vssd1 vccd1 vccd1 _12802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10442_ _10480_/S vssd1 vssd1 vccd1 vccd1 _10456_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_156_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08352__C _08360_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10373_ _10373_/A _10373_/B _10373_/C vssd1 vssd1 vccd1 vccd1 _10373_/Y sky130_fd_sc_hd__nor3_1
XFILLER_151_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12112_ _12115_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12113_/A sky130_fd_sc_hd__and2_1
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09745__A _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12043_ _12930_/Q _13369_/A vssd1 vssd1 vccd1 vccd1 _12045_/C sky130_fd_sc_hd__xor2_1
XFILLER_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09464__B _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07265__A _07291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13994_ _13994_/A _06300_/X vssd1 vssd1 vccd1 vccd1 _13994_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11656__B1 _11569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12945_ _12952_/CLK _12945_/D vssd1 vssd1 vccd1 vccd1 _14071_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12876_ _12904_/CLK _12876_/D vssd1 vssd1 vccd1 vccd1 _14004_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _14009_/Z _14009_/A _11840_/S vssd1 vssd1 vccd1 vccd1 _11828_/B sky130_fd_sc_hd__mux2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11758_ _11758_/A vssd1 vssd1 vccd1 vccd1 _12867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10709_ _10709_/A vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__clkbuf_1
X_11689_ _11689_/A _11695_/C vssd1 vssd1 vccd1 vccd1 _11690_/C sky130_fd_sc_hd__nand2_1
XFILLER_146_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13428_ _13428_/A _07810_/X vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_139_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13359_ _13359_/A _08169_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[0] sky130_fd_sc_hd__ebufn_8
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09126__A_N input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09655__A _14110_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07920_ _07920_/A vssd1 vssd1 vccd1 vccd1 _07931_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_130_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07175__A _07248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ _07851_/A vssd1 vssd1 vccd1 vccd1 _07851_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10698__A1 _10385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06802_ _06802_/A vssd1 vssd1 vccd1 vccd1 _06802_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__12917__CLK _12917_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07782_ _07782_/A _07792_/B _07787_/C vssd1 vssd1 vccd1 vccd1 _07783_/A sky130_fd_sc_hd__or3_1
Xinput2 peripheralBus_address[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09521_ _11064_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09521_/X sky130_fd_sc_hd__or2_1
X_06733_ _06733_/A _06738_/B _06738_/C vssd1 vssd1 vccd1 vccd1 _06734_/A sky130_fd_sc_hd__or3_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09452_ _09455_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09453_/A sky130_fd_sc_hd__and2_1
XFILLER_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06664_ _06673_/A _06664_/B _06664_/C vssd1 vssd1 vccd1 vccd1 _06665_/A sky130_fd_sc_hd__or3_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _12246_/Q vssd1 vssd1 vccd1 vccd1 _09321_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__11144__B _13940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09383_ _09382_/A _09379_/B _09236_/X vssd1 vssd1 vccd1 vccd1 _09384_/B sky130_fd_sc_hd__o21ai_1
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06595_ _06597_/A _06602_/B _06602_/C vssd1 vssd1 vccd1 vccd1 _06596_/A sky130_fd_sc_hd__or3_1
XFILLER_52_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08334_ _08334_/A vssd1 vssd1 vccd1 vccd1 _08334_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08734__A _13777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08265_ _08265_/A vssd1 vssd1 vccd1 vccd1 _08265_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11160__A _11160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07216_ _07220_/A _07216_/B _07228_/C vssd1 vssd1 vccd1 vccd1 _07217_/A sky130_fd_sc_hd__or3_1
X_08196_ _08196_/A vssd1 vssd1 vccd1 vccd1 _08196_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07147_ _08364_/B _07863_/B _07969_/B vssd1 vssd1 vccd1 vccd1 _07148_/A sky130_fd_sc_hd__or3_1
XFILLER_133_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08674__S0 _08602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07078_ _07120_/A vssd1 vssd1 vccd1 vccd1 _07091_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_126_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10223__B _13756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07813__A _07868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09719_ _12354_/Q _13564_/A vssd1 vssd1 vccd1 vccd1 _09719_/Y sky130_fd_sc_hd__xnor2_1
X_10991_ _11078_/A _10991_/B vssd1 vssd1 vccd1 vccd1 _10992_/A sky130_fd_sc_hd__and2_1
X_12730_ _12743_/CLK _12730_/D vssd1 vssd1 vccd1 vccd1 _12730_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12661_ _12687_/CLK _12661_/D vssd1 vssd1 vccd1 vccd1 _12661_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11616_/C _11612_/B vssd1 vssd1 vccd1 vccd1 _12832_/D sky130_fd_sc_hd__nor2_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12592_ _12598_/CLK _12592_/D vssd1 vssd1 vccd1 vccd1 _13719_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11543_ _12816_/Q vssd1 vssd1 vccd1 vccd1 _11627_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09459__B _13555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13289__445 vssd1 vssd1 vccd1 vccd1 _13289__445/HI _13994_/A sky130_fd_sc_hd__conb_1
X_11474_ _11474_/A vssd1 vssd1 vccd1 vccd1 _11489_/S sky130_fd_sc_hd__buf_2
XFILLER_109_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10425_ _10650_/A vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__clkbuf_2
X_10356_ _12514_/Q _13756_/A vssd1 vssd1 vccd1 vccd1 _10356_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_151_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10287_ _10285_/X _10278_/X _10286_/X _10283_/X vssd1 vssd1 vccd1 vccd1 _12497_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_repeater112_A peripheralBus_data[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10414__A _11189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11326__C1 _11319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ _12933_/Q _14076_/A _12029_/S vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output41_A _13596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13977_ _13977_/A _06347_/X vssd1 vssd1 vccd1 vccd1 _14009_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_74_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _12929_/CLK _12928_/D vssd1 vssd1 vccd1 vccd1 _12928_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06339__A _07045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _12904_/CLK _12859_/D vssd1 vssd1 vccd1 vccd1 _12859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06380_ _08338_/A vssd1 vssd1 vccd1 vccd1 _08349_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08050_ _08052_/A _08110_/B _08057_/C vssd1 vssd1 vccd1 vccd1 _08051_/A sky130_fd_sc_hd__or3_1
X_07001_ _07007_/A _07007_/B vssd1 vssd1 vccd1 vccd1 _07002_/A sky130_fd_sc_hd__or2_1
XFILLER_134_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08952_ _13970_/A vssd1 vssd1 vccd1 vccd1 _08952_/X sky130_fd_sc_hd__buf_2
X_07903_ _07908_/A _07903_/B _07903_/C vssd1 vssd1 vccd1 vccd1 _07904_/A sky130_fd_sc_hd__or3_1
XANTENNA__11139__B _13942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13082__238 vssd1 vssd1 vccd1 vccd1 _13082__238/HI _13577_/A sky130_fd_sc_hd__conb_1
X_08883_ _10613_/B vssd1 vssd1 vccd1 vccd1 _13754_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07834_ _07834_/A vssd1 vssd1 vccd1 vccd1 _07834_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07765_ _07765_/A vssd1 vssd1 vccd1 vccd1 _07765_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13123__279 vssd1 vssd1 vccd1 vccd1 _13123__279/HI _13664_/A sky130_fd_sc_hd__conb_1
XANTENNA__11155__A _11185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ _09631_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__or2_1
X_06716_ _06748_/A vssd1 vssd1 vccd1 vccd1 _06733_/A sky130_fd_sc_hd__clkbuf_1
X_07696_ _07699_/A _07696_/B _07704_/C vssd1 vssd1 vccd1 vccd1 _07697_/A sky130_fd_sc_hd__or3_1
XFILLER_64_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09435_ _13432_/A _12284_/Q _09448_/S vssd1 vssd1 vccd1 vccd1 _09436_/B sky130_fd_sc_hd__mux2_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06647_ _06647_/A vssd1 vssd1 vccd1 vccd1 _06647_/X sky130_fd_sc_hd__clkbuf_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13370__A _13370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _09366_/A vssd1 vssd1 vccd1 vccd1 _12266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06578_ _08035_/A vssd1 vssd1 vccd1 vccd1 _06633_/A sky130_fd_sc_hd__clkbuf_2
X_08317_ _08324_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__or2_1
XFILLER_165_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09297_ _09329_/C _09300_/C vssd1 vssd1 vccd1 vccd1 _09299_/A sky130_fd_sc_hd__and2_1
X_08248_ _08251_/A _08248_/B _08251_/C vssd1 vssd1 vccd1 vccd1 _08249_/A sky130_fd_sc_hd__or3_1
X_13017__173 vssd1 vssd1 vccd1 vccd1 _13017__173/HI _13444_/A sky130_fd_sc_hd__conb_1
XFILLER_165_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08179_ _08179_/A vssd1 vssd1 vccd1 vccd1 _08179_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10210_ _10317_/A vssd1 vssd1 vccd1 vccd1 _10298_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07808__A _08064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ _13850_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11190_/X sky130_fd_sc_hd__or2_1
XFILLER_106_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10141_ _10148_/B _10142_/B _09978_/X vssd1 vssd1 vccd1 vccd1 _10143_/A sky130_fd_sc_hd__o21ai_1
XFILLER_106_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10072_ _12447_/Q vssd1 vssd1 vccd1 vccd1 _10099_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13900_ _13900_/A _06557_/X vssd1 vssd1 vccd1 vccd1 _14028_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13831_ _13831_/A _06747_/X vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08358__B _08358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10974_ _10974_/A vssd1 vssd1 vccd1 vccd1 _12669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13762_ _13762_/A _06937_/X vssd1 vssd1 vccd1 vccd1 _14082_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ _12726_/CLK _12713_/D vssd1 vssd1 vccd1 vccd1 _13841_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ _13693_/A _07112_/X vssd1 vssd1 vccd1 vccd1 _14077_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12644_ _12647_/CLK _12644_/D vssd1 vssd1 vccd1 vccd1 _12644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _12589_/CLK _12575_/D vssd1 vssd1 vccd1 vccd1 _12575_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10409__A _10409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11526_ _11531_/C _11526_/B vssd1 vssd1 vccd1 vccd1 _12811_/D sky130_fd_sc_hd__nor2_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11457_ _11457_/A _11457_/B vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__nor2_2
X_10408_ _11184_/A vssd1 vssd1 vccd1 vccd1 _10408_/X sky130_fd_sc_hd__buf_4
X_11388_ _12761_/Q _11388_/B vssd1 vssd1 vccd1 vccd1 _11388_/X sky130_fd_sc_hd__and2_1
XFILLER_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10339_ _13659_/A _12513_/Q _10342_/S vssd1 vssd1 vccd1 vccd1 _10340_/B sky130_fd_sc_hd__mux2_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater105 peripheralBus_data[21] vssd1 vssd1 vccd1 vccd1 _13988_/Z sky130_fd_sc_hd__buf_12
XANTENNA__13455__A _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ _12928_/Q _14071_/A _12012_/S vssd1 vssd1 vccd1 vccd1 _12010_/B sky130_fd_sc_hd__mux2_1
Xrepeater116 peripheralBus_data[17] vssd1 vssd1 vccd1 vccd1 _14112_/Z sky130_fd_sc_hd__buf_12
XFILLER_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater127 _13979_/Z vssd1 vssd1 vccd1 vccd1 _14075_/Z sky130_fd_sc_hd__buf_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07550_ _07550_/A vssd1 vssd1 vccd1 vccd1 _07550_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06501_ _06528_/A vssd1 vssd1 vccd1 vccd1 _06512_/B sky130_fd_sc_hd__clkbuf_1
X_07481_ _08314_/A vssd1 vssd1 vccd1 vccd1 _08089_/A sky130_fd_sc_hd__buf_4
XFILLER_62_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09220_ _12233_/Q vssd1 vssd1 vccd1 vccd1 _09315_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__11703__A _11703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06432_ _06432_/A vssd1 vssd1 vccd1 vccd1 _06432_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09151_ _09623_/A vssd1 vssd1 vccd1 vccd1 _10648_/A sky130_fd_sc_hd__buf_4
XFILLER_147_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06363_ _06363_/A vssd1 vssd1 vccd1 vccd1 _06363_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08102_ _08102_/A vssd1 vssd1 vccd1 vccd1 _08102_/X sky130_fd_sc_hd__clkbuf_1
X_09082_ _11687_/A _12850_/Q _12851_/Q _12852_/Q _09067_/X _09068_/X vssd1 vssd1 vccd1
+ vccd1 _09082_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06294_ _08186_/A vssd1 vssd1 vccd1 vccd1 _08266_/A sky130_fd_sc_hd__clkbuf_4
X_08033_ _08039_/A _08033_/B _08044_/C vssd1 vssd1 vccd1 vccd1 _08034_/A sky130_fd_sc_hd__or3_1
XFILLER_116_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07628__A _08035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09984_ _09982_/X _09984_/B _10157_/B vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__and3b_1
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08935_ _08930_/X _08931_/X _08932_/X _08933_/X _08924_/X _08934_/X vssd1 vssd1 vccd1
+ vccd1 _08935_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10989__A _11206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13365__A _13365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08866_ _10907_/B _12652_/Q _12653_/Q _12654_/Q _08733_/X _08735_/X vssd1 vssd1 vccd1
+ vccd1 _08866_/X sky130_fd_sc_hd__mux4_2
XFILLER_84_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07363__A _07403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07817_ _07817_/A vssd1 vssd1 vccd1 vccd1 _08110_/C sky130_fd_sc_hd__clkbuf_4
X_08797_ _08788_/X _08796_/X _08863_/S vssd1 vssd1 vccd1 vccd1 _10163_/C sky130_fd_sc_hd__mux2_1
XFILLER_72_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10501__B _13747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08178__B _08358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11069__A1 _10548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ _07756_/A _07753_/B _07748_/C vssd1 vssd1 vccd1 vccd1 _07749_/A sky130_fd_sc_hd__or3_1
XFILLER_53_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07679_ _07679_/A vssd1 vssd1 vccd1 vccd1 _07679_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09418_ _13427_/A _12279_/Q _09431_/S vssd1 vssd1 vccd1 vccd1 _09419_/B sky130_fd_sc_hd__mux2_1
X_10690_ _10703_/S vssd1 vssd1 vccd1 vccd1 _10690_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09349_ _09347_/X _09372_/B _09349_/C vssd1 vssd1 vccd1 vccd1 _09350_/A sky130_fd_sc_hd__and3b_1
XFILLER_32_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12360_ _12367_/CLK _12360_/D vssd1 vssd1 vccd1 vccd1 _13489_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11311_ _10670_/X _11299_/X _11310_/X _11306_/X vssd1 vssd1 vccd1 vccd1 _12753_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12291_ _12301_/CLK _12291_/D vssd1 vssd1 vccd1 vccd1 _13570_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_4_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14030_ _14030_/A _08194_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
X_11242_ _13882_/A _12738_/Q _11248_/S vssd1 vssd1 vccd1 vccd1 _11243_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06442__A _06442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12163__B _13365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08360__C _08360_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11173_ _13844_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11173_/X sky130_fd_sc_hd__or2_1
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10124_ _10130_/C _10126_/C _10114_/X _10123_/Y vssd1 vssd1 vccd1 vccd1 _12457_/D
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__09753__A _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10055_ _10060_/C _10062_/B _10055_/C vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__and3b_1
XANTENNA__09472__B _13559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08369__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13814_ _13814_/A _06794_/X vssd1 vssd1 vccd1 vccd1 _13974_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13745_ _13745_/A _06978_/X vssd1 vssd1 vccd1 vccd1 _14097_/Z sky130_fd_sc_hd__ebufn_8
X_10957_ _10957_/A vssd1 vssd1 vccd1 vccd1 _12664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13676_ _13676_/A _07157_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
X_10888_ _10891_/B _10888_/B vssd1 vssd1 vccd1 vccd1 _12646_/D sky130_fd_sc_hd__nor2_1
X_12627_ _12647_/CLK _12627_/D vssd1 vssd1 vccd1 vccd1 _12627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12558_ _12974_/CLK _12558_/D vssd1 vssd1 vccd1 vccd1 _13686_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11509_ _11658_/A _12807_/Q _12808_/Q vssd1 vssd1 vccd1 vccd1 _11512_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12489_ _12492_/CLK _12489_/D vssd1 vssd1 vccd1 vccd1 _13619_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13345__501 vssd1 vssd1 vccd1 vccd1 _13345__501/HI _14114_/A sky130_fd_sc_hd__conb_1
XANTENNA__06352__A _06547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06981_ _08266_/A vssd1 vssd1 vccd1 vccd1 _07033_/A sky130_fd_sc_hd__buf_4
XANTENNA__09036__S0 _08941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08720_ _10148_/A _10149_/A _12465_/Q _12466_/Q _09929_/A _08709_/X vssd1 vssd1 vccd1
+ vccd1 _08720_/X sky130_fd_sc_hd__mux4_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _09397_/D vssd1 vssd1 vccd1 vccd1 _13554_/A sky130_fd_sc_hd__buf_4
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07602_ _07602_/A vssd1 vssd1 vccd1 vccd1 _07602_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08582_ _12434_/Q _12435_/Q _10029_/A _12437_/Q _08556_/X _08557_/X vssd1 vssd1 vccd1
+ vccd1 _08582_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07533_ _07533_/A vssd1 vssd1 vccd1 vccd1 _07590_/A sky130_fd_sc_hd__buf_2
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07464_ _07466_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07465_/A sky130_fd_sc_hd__or2_1
XFILLER_50_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09372_/B sky130_fd_sc_hd__buf_2
X_06415_ _06913_/A vssd1 vssd1 vccd1 vccd1 _06425_/B sky130_fd_sc_hd__clkbuf_1
X_07395_ _07395_/A vssd1 vssd1 vccd1 vccd1 _07395_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09134_ _09134_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _09161_/A sky130_fd_sc_hd__and2_1
XANTENNA__09838__A _10173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06346_ _06346_/A _06349_/B _06349_/C vssd1 vssd1 vccd1 vccd1 _06347_/A sky130_fd_sc_hd__or3_1
XANTENNA__08742__A _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09065_ _10940_/D vssd1 vssd1 vccd1 vccd1 _13946_/A sky130_fd_sc_hd__buf_4
XFILLER_147_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06277_ _11789_/A _07319_/C _11789_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11457_/B
+ sky130_fd_sc_hd__or4b_4
X_08016_ _08025_/A _08020_/B _08016_/C vssd1 vssd1 vccd1 vccd1 _08017_/A sky130_fd_sc_hd__or3_1
XFILLER_151_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07358__A _07371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13088__244 vssd1 vssd1 vccd1 vccd1 _13088__244/HI _13597_/A sky130_fd_sc_hd__conb_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08180__C _08180_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09967_ _10107_/A _09967_/B _09967_/C vssd1 vssd1 vccd1 vccd1 _09977_/A sky130_fd_sc_hd__and3_1
X_13129__285 vssd1 vssd1 vccd1 vccd1 _13129__285/HI _13670_/A sky130_fd_sc_hd__conb_1
X_08918_ _13968_/A vssd1 vssd1 vccd1 vccd1 _08918_/X sky130_fd_sc_hd__buf_4
XANTENNA__10512__A _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ _13527_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09898_/X sky130_fd_sc_hd__or2_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08849_ _10162_/C vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__buf_4
XANTENNA__10231__B _13757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _11860_/A vssd1 vssd1 vccd1 vccd1 _12890_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _10864_/B _10790_/C _10809_/C _10864_/A vssd1 vssd1 vccd1 vccd1 _10812_/C
+ sky130_fd_sc_hd__a31o_1
X_11791_ _11843_/S vssd1 vssd1 vccd1 vccd1 _11805_/S sky130_fd_sc_hd__buf_2
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ _13530_/A _07544_/X vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_8
X_10742_ _10885_/A _10806_/C _10806_/D vssd1 vssd1 vccd1 vccd1 _10742_/X sky130_fd_sc_hd__and3_1
XANTENNA__12158__B _13370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13461_ _13461_/A _07725_/X vssd1 vssd1 vccd1 vccd1 _14037_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_41_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10673_ _10673_/A vssd1 vssd1 vccd1 vccd1 _10673_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12412_ _12414_/CLK _12412_/D vssd1 vssd1 vccd1 vccd1 _13588_/A sky130_fd_sc_hd__dfxtp_2
X_13392_ _13392_/A _08365_/X vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_127_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12343_ _12367_/CLK _12343_/D vssd1 vssd1 vccd1 vccd1 _12343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12274_ _12274_/CLK _12274_/D vssd1 vssd1 vccd1 vccd1 _12274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11225_ _13877_/A _12733_/Q _11231_/S vssd1 vssd1 vccd1 vccd1 _11226_/B sky130_fd_sc_hd__mux2_1
X_14013_ _14013_/A _08123_/X vssd1 vssd1 vccd1 vccd1 _14077_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09483__A _09513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11156_ _11412_/A _11156_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _11199_/B sky130_fd_sc_hd__nor3_4
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06900__A _06900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10107_ _10107_/A _10111_/C _10133_/B vssd1 vssd1 vccd1 vccd1 _10108_/B sky130_fd_sc_hd__and3_1
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11087_ _11124_/S vssd1 vssd1 vccd1 vccd1 _11101_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10038_ _10112_/A _10053_/B _10086_/C vssd1 vssd1 vccd1 vccd1 _10045_/C sky130_fd_sc_hd__and3_1
XFILLER_64_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11150__B1 _13953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11989_ _12922_/Q _14065_/A _11995_/S vssd1 vssd1 vccd1 vccd1 _11990_/B sky130_fd_sc_hd__mux2_1
XFILLER_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11453__A1 _10552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13728_ _13728_/A _07020_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[17] sky130_fd_sc_hd__ebufn_8
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_50_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13659_ _13659_/A _07201_/X vssd1 vssd1 vccd1 vccd1 _14075_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09658__A _09711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ _07180_/A _07190_/B _07187_/C vssd1 vssd1 vccd1 vccd1 _07181_/A sky130_fd_sc_hd__or3_1
XFILLER_118_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12084__A _12084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10716__A0 _13974_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09582__A0 _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ _09834_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__and2_1
XFILLER_59_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07906__A _11154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06810__A _07857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09752_ _09750_/X _09741_/X _09751_/X _09748_/X vssd1 vssd1 vccd1 vccd1 _12360_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06964_ _06964_/A vssd1 vssd1 vccd1 vccd1 _06964_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_repeater74_A peripheralBus_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ _09848_/B vssd1 vssd1 vccd1 vccd1 _13562_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11147__B _13939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09683_ _09686_/A _09683_/B vssd1 vssd1 vccd1 vccd1 _09684_/A sky130_fd_sc_hd__and2_1
X_06895_ _06895_/A vssd1 vssd1 vccd1 vccd1 _06895_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09885__A1 _09753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _08695_/A vssd1 vssd1 vccd1 vccd1 _08634_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08565_ _12437_/Q _12438_/Q _12439_/Q _12440_/Q _08559_/X _08560_/X vssd1 vssd1 vccd1
+ vccd1 _08565_/X sky130_fd_sc_hd__mux4_2
XFILLER_70_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07516_ _07516_/A vssd1 vssd1 vccd1 vccd1 _07516_/X sky130_fd_sc_hd__clkbuf_1
X_08496_ _09362_/C _12265_/Q _09362_/A _09368_/A _08445_/X _08446_/X vssd1 vssd1 vccd1
+ vccd1 _08496_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_18_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07447_ _07454_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07448_/A sky130_fd_sc_hd__or2_1
XFILLER_13_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07378_ _07378_/A vssd1 vssd1 vccd1 vccd1 _07378_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_3_5_0_clk_A clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ _14109_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _09117_/X sky130_fd_sc_hd__or2_1
XFILLER_108_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06329_ _06333_/A _06336_/B _06336_/C vssd1 vssd1 vccd1 vccd1 _06330_/A sky130_fd_sc_hd__or3_1
XANTENNA__09287__B _09389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10507__A _11151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09048_ _09045_/X _09047_/X _13972_/A vssd1 vssd1 vccd1 vccd1 _11384_/B sky130_fd_sc_hd__mux2_4
XANTENNA__10226__B _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10707__A0 _14099_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _12664_/Q _13938_/A vssd1 vssd1 vccd1 vccd1 _11011_/D sky130_fd_sc_hd__xor2_1
XFILLER_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12961_ _12961_/CLK _12961_/D vssd1 vssd1 vccd1 vccd1 _12961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13553__A _13553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11912_ _12902_/Q _13374_/A vssd1 vssd1 vccd1 vccd1 _11915_/B sky130_fd_sc_hd__xor2_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12892_ _12895_/CLK _12892_/D vssd1 vssd1 vccd1 vccd1 _12892_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11843_ peripheralBus_data[15] _14014_/A _11843_/S vssd1 vssd1 vccd1 vccd1 _11844_/B
+ sky130_fd_sc_hd__mux2_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11073__A _11124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11435__A1 _10665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _12868_/Q _13373_/A vssd1 vssd1 vccd1 vccd1 _11775_/D sky130_fd_sc_hd__xor2_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13513_/A _07586_/X vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_14_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _10725_/A vssd1 vssd1 vccd1 vccd1 _12609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13444_ _13444_/A _07767_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
X_10656_ _10686_/B vssd1 vssd1 vccd1 vccd1 _10671_/B sky130_fd_sc_hd__clkbuf_1
X_13375_ _13375_/A _08316_/X vssd1 vssd1 vccd1 vccd1 _14111_/Z sky130_fd_sc_hd__ebufn_8
X_10587_ _10971_/A vssd1 vssd1 vccd1 vccd1 _10602_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12326_ _12331_/CLK _12326_/D vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12257_ _12264_/CLK _12257_/D vssd1 vssd1 vccd1 vccd1 _12257_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09925__B _11460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11208_ _11221_/A _11208_/B vssd1 vssd1 vccd1 vccd1 _11209_/A sky130_fd_sc_hd__and2_1
XANTENNA__07726__A _07892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12188_ _10645_/A _12182_/X _12186_/X _12187_/X vssd1 vssd1 vccd1 vccd1 _12972_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11139_ _12701_/Q _13942_/A vssd1 vssd1 vccd1 vccd1 _11143_/A sky130_fd_sc_hd__xor2_1
XFILLER_95_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06680_ _06680_/A vssd1 vssd1 vccd1 vccd1 _06692_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07461__A _07473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08276__B _08276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08350_ _08350_/A vssd1 vssd1 vccd1 vccd1 _08350_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07301_ _07301_/A vssd1 vssd1 vccd1 vccd1 _07301_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08281_ _08288_/A _08285_/B vssd1 vssd1 vccd1 vccd1 _08282_/A sky130_fd_sc_hd__or2_1
XFILLER_32_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11711__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07232_ _07232_/A vssd1 vssd1 vccd1 vccd1 _07232_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07163_ _07166_/A _07163_/B _07173_/C vssd1 vssd1 vccd1 vccd1 _07164_/A sky130_fd_sc_hd__or3_1
XFILLER_118_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07094_ _07094_/A _07105_/B _07101_/C vssd1 vssd1 vccd1 vccd1 _07095_/A sky130_fd_sc_hd__or3_1
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11158__A _13839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09804_ _09817_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__and2_1
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07996_ _07996_/A vssd1 vssd1 vccd1 vccd1 _07996_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09735_ _09735_/A _09735_/B _09735_/C _09735_/D vssd1 vssd1 vccd1 vccd1 _09736_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06947_ _06947_/A vssd1 vssd1 vccd1 vccd1 _06947_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13373__A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _09669_/A _09666_/B vssd1 vssd1 vccd1 vccd1 _09667_/A sky130_fd_sc_hd__and2_1
X_06878_ _06878_/A vssd1 vssd1 vccd1 vccd1 _06878_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07371__A _07371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08617_ _12447_/Q _12448_/Q _12449_/Q _10097_/A _08578_/X _08579_/X vssd1 vssd1 vccd1
+ vccd1 _08617_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10873__C1 _10895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09597_/A _09597_/B _09597_/C _09597_/D vssd1 vssd1 vccd1 vccd1 _09608_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _13584_/A vssd1 vssd1 vccd1 vccd1 _08708_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08479_ _08479_/A vssd1 vssd1 vccd1 vccd1 _09152_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09491__C1 _09192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13250__406 vssd1 vssd1 vccd1 vccd1 _13250__406/HI _13921_/A sky130_fd_sc_hd__conb_1
XFILLER_24_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10510_ _11285_/B _10512_/B _11410_/C vssd1 vssd1 vccd1 vccd1 _10538_/A sky130_fd_sc_hd__or3_2
X_11490_ _11490_/A _11490_/B vssd1 vssd1 vccd1 vccd1 _11491_/A sky130_fd_sc_hd__or2_1
X_10441_ _10441_/A vssd1 vssd1 vccd1 vccd1 _12537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10372_ _10372_/A _10372_/B _10372_/C _10372_/D vssd1 vssd1 vccd1 vccd1 _10373_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_156_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12111_ _12955_/Q _14097_/A _12118_/S vssd1 vssd1 vccd1 vccd1 _12112_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12042_ _12926_/Q _13365_/A vssd1 vssd1 vccd1 vccd1 _12045_/B sky130_fd_sc_hd__xor2_1
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13144__300 vssd1 vssd1 vccd1 vccd1 _13144__300/HI _13701_/A sky130_fd_sc_hd__conb_1
XANTENNA__11068__A _11195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09761__A _13492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13993_ _13993_/A _06302_/X vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_105_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ _12952_/CLK _12944_/D vssd1 vssd1 vccd1 vccd1 _14070_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08377__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__A _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _12961_/CLK _12875_/D vssd1 vssd1 vccd1 vccd1 _14003_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11826_ _11843_/S vssd1 vssd1 vccd1 vccd1 _11840_/S sky130_fd_sc_hd__buf_2
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11757_ _11757_/A _11757_/B vssd1 vssd1 vccd1 vccd1 _11758_/A sky130_fd_sc_hd__and2_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10708_ _10720_/A _10708_/B vssd1 vssd1 vccd1 vccd1 _10709_/A sky130_fd_sc_hd__or2_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11688_ _11688_/A _11688_/B _11688_/C _11688_/D vssd1 vssd1 vccd1 vccd1 _11695_/C
+ sky130_fd_sc_hd__and4_1
X_13427_ _13427_/A _07814_/X vssd1 vssd1 vccd1 vccd1 _14035_/Z sky130_fd_sc_hd__ebufn_8
X_10639_ _10639_/A _12060_/A vssd1 vssd1 vccd1 vccd1 _10686_/B sky130_fd_sc_hd__nor2_4
XANTENNA__10919__B1 _10936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11592__B1 _11505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ _12334_/CLK _12309_/D vssd1 vssd1 vccd1 vccd1 _12309_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09655__B _09655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07456__A _07468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07850_ _07962_/A _07854_/B _07852_/C vssd1 vssd1 vccd1 vccd1 _07851_/A sky130_fd_sc_hd__or3_1
XFILLER_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06801_ _06801_/A _06806_/B _06806_/C vssd1 vssd1 vccd1 vccd1 _06802_/A sky130_fd_sc_hd__or3_1
X_07781_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07792_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput3 peripheralBus_address[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
X_09520_ _13435_/A _09513_/X _09519_/X _09509_/X vssd1 vssd1 vccd1 vccd1 _12304_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06732_ _06732_/A vssd1 vssd1 vccd1 vccd1 _06732_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09451_ _13437_/A _12289_/Q _09454_/S vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__mux2_1
X_06663_ _06663_/A vssd1 vssd1 vccd1 vccd1 _06663_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08402_ _08395_/X _08398_/X _08400_/X _08401_/X _08382_/X _08383_/X vssd1 vssd1 vccd1
+ vccd1 _08402_/X sky130_fd_sc_hd__mux4_1
X_09382_ _09382_/A _09382_/B _09382_/C vssd1 vssd1 vccd1 vccd1 _09388_/C sky130_fd_sc_hd__and3_1
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06594_ _06594_/A vssd1 vssd1 vccd1 vccd1 _06594_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__12072__A1 _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08333_ _08336_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08334_/A sky130_fd_sc_hd__or2_1
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08371__S0 _08368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ _08264_/A _08274_/B _08264_/C vssd1 vssd1 vccd1 vccd1 _08265_/A sky130_fd_sc_hd__or3_1
X_07215_ _07230_/A vssd1 vssd1 vccd1 vccd1 _07228_/C sky130_fd_sc_hd__clkbuf_1
X_08195_ _08198_/A _08195_/B _08198_/C vssd1 vssd1 vccd1 vccd1 _08196_/A sky130_fd_sc_hd__or3_1
XFILLER_146_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09846__A _09846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _07146_/A vssd1 vssd1 vccd1 vccd1 _07146_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08674__S1 _08603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13368__A _13368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ _07077_/A vssd1 vssd1 vccd1 vccd1 _07077_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07366__A _07393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06270__A _08364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ _07979_/A _07979_/B vssd1 vssd1 vccd1 vccd1 _07980_/A sky130_fd_sc_hd__or2_1
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09718_ _12342_/Q _09851_/B vssd1 vssd1 vccd1 vccd1 _09718_/X sky130_fd_sc_hd__and2_1
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10990_ _13820_/A _12674_/Q _10990_/S vssd1 vssd1 vccd1 vccd1 _10991_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08197__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09649_ _09878_/A vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12660_/CLK _12660_/D vssd1 vssd1 vccd1 vccd1 _12660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11640_/B _11609_/A _11569_/X vssd1 vssd1 vccd1 vccd1 _11612_/B sky130_fd_sc_hd__o21ai_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_116_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _12251_/CLK sky130_fd_sc_hd__clkbuf_16
X_12591_ _12593_/CLK _12591_/D vssd1 vssd1 vccd1 vccd1 _13718_/A sky130_fd_sc_hd__dfxtp_1
X_11542_ _11542_/A _11542_/B vssd1 vssd1 vccd1 vccd1 _12815_/D sky130_fd_sc_hd__nor2_1
XANTENNA__11070__B _11070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11473_ _11473_/A vssd1 vssd1 vccd1 vccd1 _12796_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_2_2_0_clk_A clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09756__A _10652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ _10667_/A vssd1 vssd1 vccd1 vccd1 _10650_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09475__B _13553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10355_ _12502_/Q _13744_/A vssd1 vssd1 vccd1 vccd1 _10355_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _13627_/A _10291_/B vssd1 vssd1 vccd1 vccd1 _10286_/X sky130_fd_sc_hd__or2_1
XFILLER_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12025_ _12025_/A vssd1 vssd1 vccd1 vccd1 _12932_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_repeater105_A peripheralBus_data[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13976_ _13976_/A _06350_/X vssd1 vssd1 vccd1 vccd1 _13976_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA_output34_A _13980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12927_ _12929_/CLK _12927_/D vssd1 vssd1 vccd1 vccd1 _12927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12858_ _12961_/CLK _12858_/D vssd1 vssd1 vccd1 vccd1 _12858_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _14068_/Z _14004_/A _11823_/S vssd1 vssd1 vccd1 vccd1 _11810_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_107_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _12340_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12923_/CLK _12789_/D vssd1 vssd1 vccd1 vccd1 _13915_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10065__B1 _09994_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07000_ _07000_/A vssd1 vssd1 vccd1 vccd1 _07000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08951_ _12820_/Q _12821_/Q _12822_/Q _12823_/Q _08921_/X _08922_/X vssd1 vssd1 vccd1
+ vccd1 _08951_/X sky130_fd_sc_hd__mux4_2
XFILLER_69_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07902_ _07902_/A vssd1 vssd1 vccd1 vccd1 _07902_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08882_ _08877_/X _08880_/X _10710_/A vssd1 vssd1 vccd1 vccd1 _10613_/B sky130_fd_sc_hd__mux2_4
XFILLER_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07833_ _07843_/A _07840_/B _08180_/C vssd1 vssd1 vccd1 vccd1 _07834_/A sky130_fd_sc_hd__or3_1
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07764_ _07769_/A _07766_/B _07774_/C vssd1 vssd1 vccd1 vccd1 _07765_/A sky130_fd_sc_hd__or3_1
X_09503_ _13428_/A _09500_/X _09502_/X _09496_/X vssd1 vssd1 vccd1 vccd1 _12297_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06715_ _06715_/A vssd1 vssd1 vccd1 vccd1 _06715_/X sky130_fd_sc_hd__clkbuf_1
X_07695_ _07695_/A vssd1 vssd1 vccd1 vccd1 _07695_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09434_ _09454_/S vssd1 vssd1 vccd1 vccd1 _09448_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06646_ _06646_/A _06651_/B _06651_/C vssd1 vssd1 vccd1 vccd1 _06647_/A sky130_fd_sc_hd__or3_1
XANTENNA__08745__A _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09365_ _09380_/A _09365_/B _09365_/C vssd1 vssd1 vccd1 vccd1 _09366_/A sky130_fd_sc_hd__and3_1
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06577_ _06577_/A vssd1 vssd1 vccd1 vccd1 _08035_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__11171__A _11185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08316_ _08316_/A vssd1 vssd1 vccd1 vccd1 _08316_/X sky130_fd_sc_hd__clkbuf_1
X_09296_ _12252_/Q vssd1 vssd1 vccd1 vccd1 _09329_/C sky130_fd_sc_hd__clkbuf_1
X_08247_ _08247_/A vssd1 vssd1 vccd1 vccd1 _08247_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08178_ _08358_/A _08358_/B _08184_/C vssd1 vssd1 vccd1 vccd1 _08179_/A sky130_fd_sc_hd__or3_1
XFILLER_118_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07129_ _07129_/A vssd1 vssd1 vccd1 vccd1 _07129_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10140_ _10140_/A vssd1 vssd1 vccd1 vccd1 _12461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10234__B _13755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10071_ _10071_/A vssd1 vssd1 vccd1 vccd1 _12446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11346__A _11363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ _13830_/A _06750_/X vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_63_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08358__C _08360_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13761_ _13761_/A _06940_/X vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__ebufn_8
X_10973_ _10986_/A _10973_/B vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__and2_1
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13256__412 vssd1 vssd1 vccd1 vccd1 _13256__412/HI _13927_/A sky130_fd_sc_hd__conb_1
XANTENNA__13561__A _13561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ _12726_/CLK _12712_/D vssd1 vssd1 vccd1 vccd1 _13840_/A sky130_fd_sc_hd__dfxtp_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _13692_/A _07114_/X vssd1 vssd1 vccd1 vccd1 _14108_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12643_ _12647_/CLK _12643_/D vssd1 vssd1 vccd1 vccd1 _12643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09988__B1 _09987_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12574_ _12598_/CLK _12574_/D vssd1 vssd1 vccd1 vccd1 _12574_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11512__C _11682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11795__A0 _14064_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11525_ _11625_/D _11523_/A _11521_/X vssd1 vssd1 vccd1 vccd1 _11526_/B sky130_fd_sc_hd__o21ai_1
XFILLER_156_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09486__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11456_ _11634_/A vssd1 vssd1 vccd1 vccd1 _11689_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10407_ _09773_/X _10395_/X _10406_/X _10398_/X vssd1 vssd1 vccd1 vccd1 _12527_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11387_ _12761_/Q _11388_/B vssd1 vssd1 vccd1 vccd1 _11387_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10425__A _10650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10338_ _10338_/A vssd1 vssd1 vccd1 vccd1 _12512_/D sky130_fd_sc_hd__clkbuf_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _10667_/A vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater106 _13987_/Z vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__buf_12
X_12008_ _12008_/A vssd1 vssd1 vccd1 vccd1 _12927_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater117 _14079_/Z vssd1 vssd1 vccd1 vccd1 _13983_/Z sky130_fd_sc_hd__buf_12
Xrepeater128 peripheralBus_data[12] vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__buf_12
XFILLER_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10160__A _10160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13959_ _13959_/A _06399_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[24] sky130_fd_sc_hd__ebufn_8
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06500_ _06500_/A vssd1 vssd1 vccd1 vccd1 _06500_/X sky130_fd_sc_hd__clkbuf_1
X_07480_ _07480_/A vssd1 vssd1 vccd1 vccd1 _08314_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06431_ _06440_/A _06437_/B vssd1 vssd1 vccd1 vccd1 _06432_/A sky130_fd_sc_hd__or2_1
XFILLER_62_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09979__B1 _09978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09150_ _14066_/Z vssd1 vssd1 vccd1 vccd1 _09623_/A sky130_fd_sc_hd__buf_4
X_06362_ _06822_/A _06362_/B _06362_/C vssd1 vssd1 vccd1 vccd1 _06363_/A sky130_fd_sc_hd__or3_1
XFILLER_147_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08101_ _08101_/A _08101_/B _08105_/C vssd1 vssd1 vccd1 vccd1 _08102_/A sky130_fd_sc_hd__or3_1
X_09081_ _08972_/X _08976_/X _08975_/X _08978_/X _09024_/X _09030_/X vssd1 vssd1 vccd1
+ vccd1 _09081_/X sky130_fd_sc_hd__mux4_1
X_06293_ _06442_/A vssd1 vssd1 vccd1 vccd1 _06308_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_163_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09396__A _09867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ _08072_/A vssd1 vssd1 vccd1 vccd1 _08044_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_163_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10335__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ _09981_/B _09972_/X _09981_/A vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__a21o_1
XFILLER_115_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08934_ _13971_/A vssd1 vssd1 vccd1 vccd1 _08934_/X sky130_fd_sc_hd__buf_2
XFILLER_69_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08865_ _08765_/X _08768_/X _08771_/X _08772_/X _08826_/X _08859_/X vssd1 vssd1 vccd1
+ vccd1 _08865_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11166__A _11195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07816_ _07816_/A vssd1 vssd1 vccd1 vccd1 _07816_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10070__A _10160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08796_ _08790_/X _08791_/X _08793_/X _08795_/X _08748_/X _08749_/X vssd1 vssd1 vccd1
+ vccd1 _08796_/X sky130_fd_sc_hd__mux4_1
X_07747_ _07747_/A vssd1 vssd1 vccd1 vccd1 _07747_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08565__S0 _08559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07678_ _07686_/A _07683_/B _07678_/C vssd1 vssd1 vccd1 vccd1 _07679_/A sky130_fd_sc_hd__or3_1
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09417_ _09454_/S vssd1 vssd1 vccd1 vccd1 _09431_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06629_ _06629_/A vssd1 vssd1 vccd1 vccd1 _06629_/X sky130_fd_sc_hd__clkbuf_1
X_09348_ _09352_/C _09344_/B _09352_/B vssd1 vssd1 vccd1 vccd1 _09349_/C sky130_fd_sc_hd__a21o_1
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10229__B _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09279_ _09279_/A vssd1 vssd1 vccd1 vccd1 _12247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _13880_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11310_/X sky130_fd_sc_hd__or2_1
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12290_ _12290_/CLK _12290_/D vssd1 vssd1 vccd1 vccd1 _12290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11241_ _11363_/A vssd1 vssd1 vccd1 vccd1 _11255_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11172_ _11199_/B vssd1 vssd1 vccd1 vccd1 _11182_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_107_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13556__A _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ _10123_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _10123_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10054_ _10052_/B _10045_/X _10052_/A vssd1 vssd1 vccd1 vccd1 _10055_/C sky130_fd_sc_hd__a21o_1
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13813_ _13813_/A _06798_/X vssd1 vssd1 vccd1 vccd1 _13973_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09122__A1 _09120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13744_ _13744_/A _06980_/X vssd1 vssd1 vccd1 vccd1 _14096_/Z sky130_fd_sc_hd__ebufn_8
X_10956_ _10969_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10957_/A sky130_fd_sc_hd__and2_1
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13675_ _13675_/A _07159_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10887_ _10908_/C _10894_/D _10798_/X vssd1 vssd1 vccd1 vccd1 _10888_/B sky130_fd_sc_hd__o21ai_1
X_12626_ _12634_/CLK _12626_/D vssd1 vssd1 vccd1 vccd1 _12626_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10139__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12557_ _12974_/CLK _12557_/D vssd1 vssd1 vccd1 vccd1 _13685_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11508_ _11634_/A vssd1 vssd1 vccd1 vccd1 _11658_/A sky130_fd_sc_hd__buf_2
X_12488_ _12492_/CLK _12488_/D vssd1 vssd1 vccd1 vccd1 _13618_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_144_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11439_ _11452_/B vssd1 vssd1 vccd1 vccd1 _11450_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_125_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10743__A1 _10885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11940__A0 _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _06980_/A vssd1 vssd1 vccd1 vccd1 _06980_/X sky130_fd_sc_hd__clkbuf_1
X_14089_ _14089_/A _08145_/X vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_140_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09036__S1 _08942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08650_ _08635_/X _08648_/X _08712_/S vssd1 vssd1 vccd1 vccd1 _09397_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07601_ _07601_/A _07613_/B _07608_/C vssd1 vssd1 vccd1 vccd1 _07602_/A sky130_fd_sc_hd__or3_1
X_08581_ _12436_/Q vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11714__A _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07532_ _07532_/A vssd1 vssd1 vccd1 vccd1 _07532_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07463_ _07463_/A vssd1 vssd1 vccd1 vccd1 _07463_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _09379_/A _12228_/Q _12229_/Q vssd1 vssd1 vccd1 vccd1 _09204_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06414_ _08338_/A vssd1 vssd1 vccd1 vccd1 _06913_/A sky130_fd_sc_hd__buf_2
X_07394_ _07396_/A _07404_/B _07401_/C vssd1 vssd1 vccd1 vccd1 _07395_/A sky130_fd_sc_hd__or3_1
X_09133_ _09370_/A vssd1 vssd1 vccd1 vccd1 _09379_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06345_ _06345_/A vssd1 vssd1 vccd1 vccd1 _06345_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09064_ _09058_/X _09062_/X _09089_/S vssd1 vssd1 vccd1 vccd1 _10940_/D sky130_fd_sc_hd__mux2_1
X_06276_ input6/X vssd1 vssd1 vccd1 vccd1 _11789_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_08015_ _08015_/A vssd1 vssd1 vccd1 vccd1 _08015_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11931__A0 _14096_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13376__A _13376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _13592_/A _13591_/A _09965_/X vssd1 vssd1 vccd1 vccd1 _09967_/C sky130_fd_sc_hd__or3b_1
XFILLER_89_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08917_ _12811_/Q _12812_/Q _12813_/Q _12814_/Q _08915_/X _08916_/X vssd1 vssd1 vccd1
+ vccd1 _08917_/X sky130_fd_sc_hd__mux4_1
X_09897_ _09767_/X _09888_/X _09896_/X _09892_/X vssd1 vssd1 vccd1 vccd1 _12398_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _12356_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08189__B _08189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_clk_A clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ _08844_/X _08847_/X _08863_/S vssd1 vssd1 vccd1 vccd1 _10162_/C sky130_fd_sc_hd__mux2_1
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08779_ _08886_/A vssd1 vssd1 vccd1 vccd1 _08779_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _10872_/A _10880_/C vssd1 vssd1 vccd1 vccd1 _10878_/B sky130_fd_sc_hd__and2_1
X_11790_ _11790_/A _11924_/B _11924_/C vssd1 vssd1 vccd1 vccd1 _11843_/S sky130_fd_sc_hd__or3_2
XFILLER_150_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ _10915_/A vssd1 vssd1 vccd1 vccd1 _10885_/A sky130_fd_sc_hd__buf_2
XFILLER_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13460_ _13460_/A _07728_/X vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_8
X_10672_ _10670_/X _10655_/X _10671_/X _10668_/X vssd1 vssd1 vccd1 vccd1 _12593_/D
+ sky130_fd_sc_hd__o211a_1
X_12411_ _12418_/CLK _12411_/D vssd1 vssd1 vccd1 vccd1 _13587_/A sky130_fd_sc_hd__dfxtp_1
X_13391_ _13391_/A _08161_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[0] sky130_fd_sc_hd__ebufn_8
XFILLER_154_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk _12881_/CLK vssd1 vssd1 vccd1 vccd1 _12929_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08710__S0 _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12342_ _12367_/CLK _12342_/D vssd1 vssd1 vccd1 vccd1 _12342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12174__B _13363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12273_ _12274_/CLK _12273_/D vssd1 vssd1 vccd1 vccd1 _12273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14012_ _14012_/A _08129_/X vssd1 vssd1 vccd1 vccd1 _14012_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA_clkbuf_4_12_0_clk_A clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ _11363_/A vssd1 vssd1 vccd1 vccd1 _11239_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09764__A _13493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11155_ _11185_/A vssd1 vssd1 vccd1 vccd1 _11155_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10106_ _09982_/A _10133_/B _10111_/C vssd1 vssd1 vccd1 vccd1 _10108_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11086_ _11086_/A vssd1 vssd1 vccd1 vccd1 _12697_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_87_clk _12438_/CLK vssd1 vssd1 vccd1 vccd1 _12451_/CLK sky130_fd_sc_hd__clkbuf_16
X_10037_ _10097_/B _10097_/C vssd1 vssd1 vccd1 vccd1 _10086_/C sky130_fd_sc_hd__and2_1
XFILLER_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11988_ _11988_/A vssd1 vssd1 vccd1 vccd1 _12921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13727_ _13727_/A _07024_/X vssd1 vssd1 vccd1 vccd1 _13983_/Z sky130_fd_sc_hd__ebufn_8
X_10939_ _10939_/A _10939_/B _10939_/C _10939_/D vssd1 vssd1 vccd1 vccd1 _10942_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__09939__A _09939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13658_ _13658_/A _07204_/X vssd1 vssd1 vccd1 vccd1 _14106_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _12811_/CLK _12609_/D vssd1 vssd1 vccd1 vccd1 _13784_/A sky130_fd_sc_hd__dfxtp_1
X_13589_ _13589_/A _07395_/X vssd1 vssd1 vccd1 vccd1 _14037_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_129_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_clk _12917_/CLK vssd1 vssd1 vccd1 vccd1 _12908_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ _13527_/A _12382_/Q _09820_/S vssd1 vssd1 vccd1 vccd1 _09821_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13161__317 vssd1 vssd1 vccd1 vccd1 _13161__317/HI _13734_/A sky130_fd_sc_hd__conb_1
X_09751_ _13489_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09751_/X sky130_fd_sc_hd__or2_1
XFILLER_113_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06963_ _06972_/A _06965_/B vssd1 vssd1 vccd1 vccd1 _06964_/A sky130_fd_sc_hd__or2_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_78_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _12652_/CLK sky130_fd_sc_hd__clkbuf_16
X_08702_ _08696_/X _08700_/X _09941_/A vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__mux2_2
XANTENNA__13924__A _13924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ _13494_/A _12348_/Q _09685_/S vssd1 vssd1 vccd1 vccd1 _09683_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06894_ _07328_/A _06898_/B _06898_/C vssd1 vssd1 vccd1 vccd1 _06895_/A sky130_fd_sc_hd__or3_1
XFILLER_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08633_ _13587_/A vssd1 vssd1 vccd1 vccd1 _08695_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater67_A _14070_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202__358 vssd1 vssd1 vccd1 vccd1 _13202__358/HI _13825_/A sky130_fd_sc_hd__conb_1
XFILLER_82_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11444__A _12084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _08552_/X _08555_/X _08558_/X _08561_/X _08670_/A _08563_/X vssd1 vssd1 vccd1
+ vccd1 _08564_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07515_ _07517_/A _07517_/B _07524_/C vssd1 vssd1 vccd1 vccd1 _07516_/A sky130_fd_sc_hd__or3_1
X_08495_ _12267_/Q vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13055__211 vssd1 vssd1 vccd1 vccd1 _13055__211/HI _13514_/A sky130_fd_sc_hd__conb_1
X_07446_ _07446_/A vssd1 vssd1 vccd1 vccd1 _07446_/X sky130_fd_sc_hd__clkbuf_1
X_07377_ _07382_/A _07377_/B _07388_/C vssd1 vssd1 vccd1 vccd1 _07378_/A sky130_fd_sc_hd__or3_1
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09116_ _10548_/A vssd1 vssd1 vccd1 vccd1 _09116_/X sky130_fd_sc_hd__clkbuf_8
X_06328_ _06328_/A vssd1 vssd1 vccd1 vccd1 _06328_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09047_ _08959_/X _08960_/X _09020_/X _09046_/X _09030_/A _08934_/X vssd1 vssd1 vccd1
+ vccd1 _09047_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10523__A _10650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09949_ _09949_/A vssd1 vssd1 vccd1 vccd1 _12414_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_69_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _12802_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_161_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12960_ _12962_/CLK _12960_/D vssd1 vssd1 vccd1 vccd1 _12960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11911_ _12889_/Q _13361_/A vssd1 vssd1 vccd1 vccd1 _11915_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07832__A _08335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12895_/CLK _12891_/D vssd1 vssd1 vccd1 vccd1 _12891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11842_/A vssd1 vssd1 vccd1 vccd1 _12885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12169__B _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _12864_/Q _13369_/A vssd1 vssd1 vccd1 vccd1 _11775_/C sky130_fd_sc_hd__xor2_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _13512_/A _07589_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09759__A _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _11481_/A _10724_/B vssd1 vssd1 vccd1 vccd1 _10725_/A sky130_fd_sc_hd__or2_1
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13443_ _13443_/A _07770_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
X_10655_ _10673_/A vssd1 vssd1 vccd1 vccd1 _10655_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_127_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13374_ _13374_/A _08313_/X vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_70_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10586_ _10586_/A vssd1 vssd1 vccd1 vccd1 _12575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12325_ _12325_/CLK _12325_/D vssd1 vssd1 vccd1 vccd1 _13455_/A sky130_fd_sc_hd__dfxtp_2
XANTENNA_repeater135_A peripheralBus_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09494__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12256_ _12258_/CLK _12256_/D vssd1 vssd1 vccd1 vccd1 _12256_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06911__A _08168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ _13872_/A _12728_/Q _11281_/B vssd1 vssd1 vccd1 vccd1 _11208_/B sky130_fd_sc_hd__mux2_1
XFILLER_122_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12187_ _12200_/A vssd1 vssd1 vccd1 vccd1 _12187_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11138_ _11138_/A _11138_/B _11138_/C _11138_/D vssd1 vssd1 vccd1 vccd1 _11149_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13744__A _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11069_ _10548_/X _11055_/X _11067_/X _11068_/X vssd1 vssd1 vccd1 vccd1 _12692_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_0_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _12274_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10882__B1 _10798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07300_ _07307_/A _07303_/B _07300_/C vssd1 vssd1 vccd1 vccd1 _07301_/A sky130_fd_sc_hd__or3_1
XANTENNA__10634__B1 _13759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08280_ _08280_/A vssd1 vssd1 vccd1 vccd1 _08280_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07231_ _07239_/A _07231_/B _07246_/C vssd1 vssd1 vccd1 vccd1 _07232_/A sky130_fd_sc_hd__or3_1
X_07162_ _07162_/A vssd1 vssd1 vccd1 vccd1 _07173_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__09252__B1 _09248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07093_ _07120_/A vssd1 vssd1 vccd1 vccd1 _07105_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_117_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06821__A _06967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09803_ _13522_/A _12377_/Q _09871_/B vssd1 vssd1 vccd1 vccd1 _09804_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07995_ _08180_/A _07995_/B _08180_/C vssd1 vssd1 vccd1 vccd1 _07996_/A sky130_fd_sc_hd__or3_1
XFILLER_75_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ _12345_/Q _13555_/A vssd1 vssd1 vccd1 vccd1 _09735_/D sky130_fd_sc_hd__xor2_1
XFILLER_28_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09851__B _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06946_ _06948_/A _06953_/B vssd1 vssd1 vccd1 vccd1 _06947_/A sky130_fd_sc_hd__or2_1
XFILLER_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ _13489_/A _12343_/Q _09738_/B vssd1 vssd1 vccd1 vccd1 _09666_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06877_ _06877_/A _06884_/B _06884_/C vssd1 vssd1 vccd1 vccd1 _06878_/A sky130_fd_sc_hd__or3_1
X_08616_ _12450_/Q vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09596_ _12322_/Q _13565_/A vssd1 vssd1 vccd1 vccd1 _09597_/D sky130_fd_sc_hd__xor2_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06268__A _11457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _12424_/Q vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08478_ _11705_/B vssd1 vssd1 vccd1 vccd1 _13364_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07429_ _07429_/A vssd1 vssd1 vccd1 vccd1 _07429_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10440_ _10444_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__and2_1
XFILLER_6_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13330__486 vssd1 vssd1 vccd1 vccd1 _13330__486/HI _14083_/A sky130_fd_sc_hd__conb_1
XFILLER_164_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _12501_/Q _13743_/A vssd1 vssd1 vccd1 vccd1 _10372_/D sky130_fd_sc_hd__xor2_1
XFILLER_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ _12110_/A vssd1 vssd1 vccd1 vccd1 _12954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12041_ _12923_/Q _13362_/A vssd1 vssd1 vccd1 vccd1 _12045_/A sky130_fd_sc_hd__xor2_1
XFILLER_78_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13564__A _13564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13992_ _13992_/A _06304_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_19_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224__380 vssd1 vssd1 vccd1 vccd1 _13224__380/HI _13863_/A sky130_fd_sc_hd__conb_1
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12943_ _12946_/CLK _12943_/D vssd1 vssd1 vccd1 vccd1 _14069_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_64_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ _12904_/CLK _12874_/D vssd1 vssd1 vccd1 vccd1 _14002_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _11825_/A vssd1 vssd1 vccd1 vccd1 _12880_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11756_ _12867_/Q _14012_/A _11760_/S vssd1 vssd1 vccd1 vccd1 _11757_/B sky130_fd_sc_hd__mux2_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06906__A _06955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_79_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _14099_/Z _08876_/X _10723_/S vssd1 vssd1 vccd1 vccd1 _10708_/B sky130_fd_sc_hd__mux2_1
X_11687_ _11687_/A _11687_/B _11687_/C vssd1 vssd1 vccd1 vccd1 _11688_/D sky130_fd_sc_hd__and3_1
XANTENNA__10428__A _13786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13426_ _13426_/A _07816_/X vssd1 vssd1 vccd1 vccd1 _14034_/Z sky130_fd_sc_hd__ebufn_8
X_10638_ _10673_/A vssd1 vssd1 vccd1 vccd1 _10638_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10569_ _10988_/A vssd1 vssd1 vccd1 vccd1 _10971_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12308_ _12313_/CLK _12308_/D vssd1 vssd1 vccd1 vccd1 _12308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06641__A _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11259__A _12740_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12239_ _12242_/CLK _12239_/D vssd1 vssd1 vccd1 vccd1 _12239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06800_ _06800_/A vssd1 vssd1 vccd1 vccd1 _06800_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07780_ _07780_/A vssd1 vssd1 vccd1 vccd1 _07780_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput4 peripheralBus_address[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10910__B1_N _10820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06731_ _06733_/A _06738_/B _06738_/C vssd1 vssd1 vccd1 vccd1 _06732_/A sky130_fd_sc_hd__or3_1
XANTENNA__11706__B _11706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09450_ _09450_/A vssd1 vssd1 vccd1 vccd1 _12288_/D sky130_fd_sc_hd__clkbuf_1
X_06662_ _06673_/A _06664_/B _06664_/C vssd1 vssd1 vccd1 vccd1 _06663_/A sky130_fd_sc_hd__or3_1
XFILLER_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08401_ _12241_/Q _12242_/Q _12243_/Q _12244_/Q _08376_/X _08377_/X vssd1 vssd1 vccd1
+ vccd1 _08401_/X sky130_fd_sc_hd__mux4_2
X_09381_ _09381_/A vssd1 vssd1 vccd1 vccd1 _12270_/D sky130_fd_sc_hd__clkbuf_1
X_13273__429 vssd1 vssd1 vccd1 vccd1 _13273__429/HI _13964_/A sky130_fd_sc_hd__conb_1
X_06593_ _06597_/A _06602_/B _06602_/C vssd1 vssd1 vccd1 vccd1 _06594_/A sky130_fd_sc_hd__or3_1
X_08332_ _08332_/A vssd1 vssd1 vccd1 vccd1 _08332_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11280__B1 _13952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08371__S1 _08370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08263_ _08263_/A vssd1 vssd1 vccd1 vccd1 _08274_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_4_0_0_clk_A clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07214_ _07214_/A vssd1 vssd1 vccd1 vccd1 _07214_/X sky130_fd_sc_hd__clkbuf_1
X_08194_ _08194_/A vssd1 vssd1 vccd1 vccd1 _08194_/X sky130_fd_sc_hd__clkbuf_1
X_07145_ _07152_/A _07145_/B _07160_/C vssd1 vssd1 vccd1 vccd1 _07146_/A sky130_fd_sc_hd__or3_1
XFILLER_105_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07076_ _07079_/A _07076_/B _07088_/C vssd1 vssd1 vccd1 vccd1 _07077_/A sky130_fd_sc_hd__or3_1
X_13167__323 vssd1 vssd1 vccd1 vccd1 _13167__323/HI _13740_/A sky130_fd_sc_hd__conb_1
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13208__364 vssd1 vssd1 vccd1 vccd1 _13208__364/HI _13831_/A sky130_fd_sc_hd__conb_1
XFILLER_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07978_ _07978_/A vssd1 vssd1 vccd1 vccd1 _07978_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09717_ _12342_/Q _13552_/A vssd1 vssd1 vccd1 vccd1 _09717_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06929_ _06936_/A _06929_/B vssd1 vssd1 vccd1 vccd1 _06930_/A sky130_fd_sc_hd__or2_1
XFILLER_67_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ _10667_/A vssd1 vssd1 vccd1 vccd1 _09878_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10846__B1 _10781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09579_/A _09579_/B vssd1 vssd1 vccd1 vccd1 _09580_/A sky130_fd_sc_hd__and2_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11640_/B _11640_/C _11610_/C vssd1 vssd1 vccd1 vccd1 _11616_/C sky130_fd_sc_hd__and3_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12593_/CLK _12590_/D vssd1 vssd1 vccd1 vccd1 _13717_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06726__A _11790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ _11627_/D _11547_/D _11540_/X vssd1 vssd1 vccd1 vccd1 _11542_/B sky130_fd_sc_hd__o21ai_1
XFILLER_156_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10248__A _11028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11472_ _11481_/A _11472_/B vssd1 vssd1 vccd1 vccd1 _11473_/A sky130_fd_sc_hd__or2_1
XFILLER_149_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13559__A _13559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _13662_/A _10423_/B vssd1 vssd1 vccd1 vccd1 _10423_/X sky130_fd_sc_hd__or2_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10354_ _12502_/Q _10614_/B vssd1 vssd1 vccd1 vccd1 _10354_/X sky130_fd_sc_hd__and2_1
XFILLER_152_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10285_ _11061_/A vssd1 vssd1 vccd1 vccd1 _10285_/X sky130_fd_sc_hd__buf_4
XANTENNA__11326__A1 _10552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12024_ _12030_/A _12024_/B vssd1 vssd1 vccd1 vccd1 _12025_/A sky130_fd_sc_hd__and2_1
XFILLER_104_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10711__A _11039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13975_ _13975_/A _06354_/X vssd1 vssd1 vccd1 vccd1 _14103_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_34_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12926_ _12929_/CLK _12926_/D vssd1 vssd1 vccd1 vccd1 _12926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09711__S _09711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12857_ _12873_/CLK _12857_/D vssd1 vssd1 vccd1 vccd1 _12857_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13001__157 vssd1 vssd1 vccd1 vccd1 _13001__157/HI _13412_/A sky130_fd_sc_hd__conb_1
XFILLER_21_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11808_ _11843_/S vssd1 vssd1 vccd1 vccd1 _11823_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__06636__A input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _12938_/CLK _12788_/D vssd1 vssd1 vccd1 vccd1 _13914_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11261__B _11388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11739_ _12862_/Q _14007_/A _11743_/S vssd1 vssd1 vccd1 vccd1 _11740_/B sky130_fd_sc_hd__mux2_1
XFILLER_159_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09207__B1 _09206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09758__A1 _09756_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13469__A _13469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ _13409_/A _08100_/X vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_128_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08950_ _12816_/Q _12817_/Q _11562_/C _12819_/Q _08915_/X _08916_/X vssd1 vssd1 vccd1
+ vccd1 _08950_/X sky130_fd_sc_hd__mux4_2
XANTENNA__11317__A1 _11189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07901_ _07908_/A _07903_/B _07903_/C vssd1 vssd1 vccd1 vccd1 _07902_/A sky130_fd_sc_hd__or3_1
XFILLER_102_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08881_ _13780_/A vssd1 vssd1 vccd1 vccd1 _10710_/A sky130_fd_sc_hd__buf_2
XFILLER_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09930__A1 _09139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__A _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07832_ _08335_/A vssd1 vssd1 vccd1 vccd1 _08180_/C sky130_fd_sc_hd__buf_2
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07763_ _07763_/A vssd1 vssd1 vccd1 vccd1 _07774_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09502_ _11170_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09502_/X sky130_fd_sc_hd__or2_1
X_06714_ _06714_/A _06719_/B _06719_/C vssd1 vssd1 vccd1 vccd1 _06715_/A sky130_fd_sc_hd__or3_1
XFILLER_37_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07694_ _07699_/A _07696_/B _07704_/C vssd1 vssd1 vccd1 vccd1 _07695_/A sky130_fd_sc_hd__or3_1
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09433_ _09433_/A vssd1 vssd1 vccd1 vccd1 _12283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06645_ _06645_/A vssd1 vssd1 vccd1 vccd1 _06645_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _09379_/A _09364_/B vssd1 vssd1 vccd1 vccd1 _09365_/C sky130_fd_sc_hd__nand2_1
X_06576_ _06604_/A vssd1 vssd1 vccd1 vccd1 _06589_/B sky130_fd_sc_hd__clkbuf_1
X_08315_ _08324_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08316_/A sky130_fd_sc_hd__or2_1
X_09295_ _09295_/A vssd1 vssd1 vccd1 vccd1 _12251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08246_ _08251_/A _08248_/B _08251_/C vssd1 vssd1 vccd1 vccd1 _08247_/A sky130_fd_sc_hd__or3_1
XFILLER_21_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09749__A1 _09139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ _08177_/A vssd1 vssd1 vccd1 vccd1 _08358_/B sky130_fd_sc_hd__buf_2
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07128_ _07135_/A _07131_/B _07128_/C vssd1 vssd1 vccd1 vccd1 _07129_/A sky130_fd_sc_hd__or3_1
XFILLER_118_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06281__A input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07059_ _08266_/A vssd1 vssd1 vccd1 vccd1 _08364_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10070_ _10160_/A _10070_/B _10070_/C vssd1 vssd1 vccd1 vccd1 _10071_/A sky130_fd_sc_hd__and3_1
XFILLER_0_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13760_ _13760_/A _06942_/X vssd1 vssd1 vccd1 vccd1 _14112_/Z sky130_fd_sc_hd__ebufn_8
X_10972_ _13815_/A _12669_/Q _10972_/S vssd1 vssd1 vccd1 vccd1 _10973_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09685__A0 _13495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13295__451 vssd1 vssd1 vccd1 vccd1 _13295__451/HI _14016_/A sky130_fd_sc_hd__conb_1
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ _12726_/CLK _12711_/D vssd1 vssd1 vccd1 vccd1 _13839_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13691_ _13691_/A _07116_/X vssd1 vssd1 vccd1 vccd1 _14075_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_70_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12642_ _12813_/CLK _12642_/D vssd1 vssd1 vccd1 vccd1 _12642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13336__492 vssd1 vssd1 vccd1 vccd1 _13336__492/HI _14089_/A sky130_fd_sc_hd__conb_1
XFILLER_157_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12573_ _12598_/CLK _12573_/D vssd1 vssd1 vccd1 vccd1 _12573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09767__A _10662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ _11680_/A _11625_/D _11628_/A vssd1 vssd1 vccd1 vccd1 _11531_/C sky130_fd_sc_hd__and3_1
X_11455_ _11680_/A vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__buf_2
XANTENNA__10706__A _10706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _13656_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10406_/X sky130_fd_sc_hd__or2_1
XFILLER_137_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11386_ _12773_/Q _11386_/B vssd1 vssd1 vccd1 vccd1 _11386_/X sky130_fd_sc_hd__and2_1
XFILLER_140_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10337_ _10349_/A _10337_/B vssd1 vssd1 vccd1 vccd1 _10338_/A sky130_fd_sc_hd__and2_1
XFILLER_98_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _13621_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10268_/X sky130_fd_sc_hd__or2_1
XFILLER_105_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09912__A1 _09112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ _12013_/A _12007_/B vssd1 vssd1 vccd1 vccd1 _12008_/A sky130_fd_sc_hd__and2_1
Xrepeater107 peripheralBus_data[20] vssd1 vssd1 vccd1 vccd1 _13987_/Z sky130_fd_sc_hd__buf_12
Xrepeater118 peripheralBus_data[16] vssd1 vssd1 vccd1 vccd1 _14079_/Z sky130_fd_sc_hd__buf_12
X_10199_ _10199_/A vssd1 vssd1 vccd1 vccd1 _12476_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater129 peripheralBus_data[12] vssd1 vssd1 vccd1 vccd1 _13979_/Z sky130_fd_sc_hd__buf_12
XFILLER_66_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13752__A _13752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__A0 _13492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13958_ _13958_/A _06401_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[23] sky130_fd_sc_hd__ebufn_8
XANTENNA__11483__A0 _13974_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ _12919_/CLK _12909_/D vssd1 vssd1 vccd1 vccd1 _14036_/A sky130_fd_sc_hd__dfxtp_1
X_13889_ _13889_/A _06588_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[18] sky130_fd_sc_hd__ebufn_8
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06430_ _06442_/A vssd1 vssd1 vccd1 vccd1 _06440_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06366__A _06547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06361_ _06361_/A vssd1 vssd1 vccd1 vccd1 _06822_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09099__D _12062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ _08100_/A vssd1 vssd1 vccd1 vccd1 _08100_/X sky130_fd_sc_hd__clkbuf_1
X_09080_ _11386_/B vssd1 vssd1 vccd1 vccd1 _13948_/A sky130_fd_sc_hd__buf_2
X_06292_ _06292_/A vssd1 vssd1 vccd1 vccd1 _06292_/X sky130_fd_sc_hd__clkbuf_1
X_08031_ _08031_/A vssd1 vssd1 vccd1 vccd1 _08031_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09982_ _09982_/A _10030_/A vssd1 vssd1 vccd1 vccd1 _09982_/X sky130_fd_sc_hd__and2_1
XFILLER_115_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08933_ _12835_/Q _12836_/Q _12837_/Q _12838_/Q _08921_/X _08922_/X vssd1 vssd1 vccd1
+ vccd1 _08933_/X sky130_fd_sc_hd__mux4_2
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08864_ _10164_/A vssd1 vssd1 vccd1 vccd1 _13751_/A sky130_fd_sc_hd__buf_6
X_07815_ _07868_/A _07820_/B _07815_/C vssd1 vssd1 vccd1 vccd1 _07816_/A sky130_fd_sc_hd__or3_1
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08795_ _12644_/Q _12645_/Q _12646_/Q _10908_/B _08785_/X _08786_/X vssd1 vssd1 vccd1
+ vccd1 _08795_/X sky130_fd_sc_hd__mux4_2
XFILLER_123_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13279__435 vssd1 vssd1 vccd1 vccd1 _13279__435/HI _13984_/A sky130_fd_sc_hd__conb_1
X_07746_ _07756_/A _07753_/B _07748_/C vssd1 vssd1 vccd1 vccd1 _07747_/A sky130_fd_sc_hd__or3_1
XFILLER_53_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10277__A1 _09773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__S1 _08560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ _07677_/A vssd1 vssd1 vccd1 vccd1 _07677_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09416_ _09416_/A vssd1 vssd1 vccd1 vccd1 _12278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06628_ _06646_/A _06630_/B _06630_/C vssd1 vssd1 vccd1 vccd1 _06629_/A sky130_fd_sc_hd__or3_1
X_09347_ _09347_/A _09363_/A _09368_/C vssd1 vssd1 vccd1 vccd1 _09347_/X sky130_fd_sc_hd__and3_1
X_06559_ _06569_/A _06561_/B _06561_/C vssd1 vssd1 vccd1 vccd1 _06560_/A sky130_fd_sc_hd__or3_1
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12993__149 vssd1 vssd1 vccd1 vccd1 _12993__149/HI _13390_/A sky130_fd_sc_hd__conb_1
XFILLER_21_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ _09276_/X _09389_/A _09278_/C vssd1 vssd1 vccd1 vccd1 _09279_/A sky130_fd_sc_hd__and3b_1
XFILLER_148_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08229_ _08238_/A _08235_/B _08238_/C vssd1 vssd1 vccd1 vccd1 _08230_/A sky130_fd_sc_hd__or3_1
XANTENNA__11121__S _11124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ _11240_/A vssd1 vssd1 vccd1 vccd1 _12737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11171_ _11185_/A vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10122_ _10126_/C _10126_/D _10130_/C vssd1 vssd1 vccd1 vccd1 _10123_/B sky130_fd_sc_hd__a21o_1
XFILLER_106_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10053_ _13583_/A _10053_/B _10086_/C _10100_/A vssd1 vssd1 vccd1 vccd1 _10060_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input26_A peripheralBus_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13812_ _13812_/A _06800_/X vssd1 vssd1 vccd1 vccd1 _14068_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_29_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10955_ _13810_/A _12664_/Q _10955_/S vssd1 vssd1 vccd1 vccd1 _10956_/B sky130_fd_sc_hd__mux2_1
X_13743_ _13743_/A _07970_/X vssd1 vssd1 vccd1 vccd1 _13775_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13674_ _13674_/A _07161_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
X_10886_ _10915_/A _10922_/B vssd1 vssd1 vccd1 vccd1 _10894_/D sky130_fd_sc_hd__and2_1
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ _12625_/CLK _12625_/D vssd1 vssd1 vccd1 vccd1 _12625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13072__228 vssd1 vssd1 vccd1 vccd1 _13072__228/HI _13547_/A sky130_fd_sc_hd__conb_1
XFILLER_8_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ _12565_/CLK _12556_/D vssd1 vssd1 vccd1 vccd1 _13684_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11507_ _11634_/A _12808_/Q _12807_/Q vssd1 vssd1 vccd1 vccd1 _11514_/B sky130_fd_sc_hd__and3_1
XFILLER_157_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12487_ _12492_/CLK _12487_/D vssd1 vssd1 vccd1 vccd1 _13617_/A sky130_fd_sc_hd__dfxtp_1
X_13113__269 vssd1 vssd1 vccd1 vccd1 _13113__269/HI _13638_/A sky130_fd_sc_hd__conb_1
X_11438_ _11438_/A vssd1 vssd1 vccd1 vccd1 _11438_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13747__A _13747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11369_ _11369_/A vssd1 vssd1 vccd1 vccd1 _12771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _14088_/A _08143_/X vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__ebufn_8
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07600_ _07615_/A vssd1 vssd1 vccd1 vccd1 _07613_/B sky130_fd_sc_hd__clkbuf_1
X_08580_ _12430_/Q _12431_/Q _12432_/Q _12433_/Q _08578_/X _08579_/X vssd1 vssd1 vccd1
+ vccd1 _08580_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13007__163 vssd1 vssd1 vccd1 vccd1 _13007__163/HI _13418_/A sky130_fd_sc_hd__conb_1
XANTENNA__10259__A1 _09750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07480__A _07480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07531_ _07531_/A _07531_/B _07538_/C vssd1 vssd1 vccd1 vccd1 _07532_/A sky130_fd_sc_hd__or3_1
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07462_ _07466_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07463_/A sky130_fd_sc_hd__or2_1
XFILLER_62_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09201_ _09269_/A _12229_/Q _12228_/Q vssd1 vssd1 vccd1 vccd1 _09201_/X sky130_fd_sc_hd__and3_1
X_06413_ _06413_/A vssd1 vssd1 vccd1 vccd1 _06413_/X sky130_fd_sc_hd__clkbuf_1
X_07393_ _07393_/A vssd1 vssd1 vccd1 vccd1 _07404_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09132_ _09269_/A vssd1 vssd1 vccd1 vccd1 _09370_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06344_ _06346_/A _06349_/B _06349_/C vssd1 vssd1 vccd1 vccd1 _06345_/A sky130_fd_sc_hd__or3_1
XANTENNA__06824__A _09125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ _13972_/A vssd1 vssd1 vccd1 vccd1 _09089_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06275_ input7/X vssd1 vssd1 vccd1 vccd1 _11789_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08014_ _08025_/A _08020_/B _08016_/C vssd1 vssd1 vccd1 vccd1 _08015_/A sky130_fd_sc_hd__or3_1
XFILLER_118_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09854__B _13561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11931__A1 _14032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09965_ _09851_/B _09397_/C _09397_/D _09867_/B _13589_/A _13590_/A vssd1 vssd1 vccd1
+ vccd1 _09965_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08916_ _13969_/A vssd1 vssd1 vccd1 vccd1 _08916_/X sky130_fd_sc_hd__buf_2
XFILLER_134_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09896_ _13526_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09896_/X sky130_fd_sc_hd__or2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10512__C _11156_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08847_ _08791_/X _08795_/X _08793_/X _08846_/X _08837_/X _08838_/X vssd1 vssd1 vccd1
+ vccd1 _08847_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08778_ _10614_/B vssd1 vssd1 vccd1 vccd1 _13744_/A sky130_fd_sc_hd__buf_4
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07390__A _07403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _07729_/A vssd1 vssd1 vccd1 vccd1 _07742_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10740_ _10806_/D _10895_/A vssd1 vssd1 vccd1 vccd1 _12614_/D sky130_fd_sc_hd__nor2_1
XFILLER_41_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _13720_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10671_/X sky130_fd_sc_hd__or2_1
XFILLER_41_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12410_ _12470_/CLK _12410_/D vssd1 vssd1 vccd1 vccd1 _13586_/A sky130_fd_sc_hd__dfxtp_2
X_13390_ _13390_/A _08350_/X vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__ebufn_8
X_12341_ _12349_/CLK _12341_/D vssd1 vssd1 vccd1 vccd1 _12341_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10422__A1 _09116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06453__B _07845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12272_ _12274_/CLK _12272_/D vssd1 vssd1 vccd1 vccd1 _12272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14011_ _14011_/A _08074_/X vssd1 vssd1 vccd1 vccd1 _14075_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__13567__A _13567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _11929_/A vssd1 vssd1 vccd1 vccd1 _11363_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_153_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11154_ _11410_/A _11154_/B _11410_/C vssd1 vssd1 vccd1 vccd1 _11185_/A sky130_fd_sc_hd__or3_4
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11087__A _11124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10105_ _10105_/A vssd1 vssd1 vccd1 vccd1 _12452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11085_ _11095_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11086_/A sky130_fd_sc_hd__and2_1
XFILLER_88_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10036_ _10097_/C _10089_/A _10035_/Y vssd1 vssd1 vccd1 vccd1 _12437_/D sky130_fd_sc_hd__a21oi_1
XFILLER_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06909__A _08168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ _11996_/A _11987_/B vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__and2_1
XFILLER_16_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ _13726_/A _07026_/X vssd1 vssd1 vccd1 vccd1 _14078_/Z sky130_fd_sc_hd__ebufn_8
X_10938_ _10938_/A _10938_/B _10938_/C _10938_/D vssd1 vssd1 vccd1 vccd1 _10942_/A
+ sky130_fd_sc_hd__or4_1
XANTENNA__10661__A1 _10659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13657_ _13657_/A _07207_/X vssd1 vssd1 vccd1 vccd1 _14105_/Z sky130_fd_sc_hd__ebufn_8
X_10869_ _10876_/C _10869_/B _10869_/C _10869_/D vssd1 vssd1 vccd1 vccd1 _10871_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_83_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12608_ _12811_/CLK _12608_/D vssd1 vssd1 vccd1 vccd1 _13783_/A sky130_fd_sc_hd__dfxtp_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13588_ _13588_/A _07397_/X vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10413__A1 _10408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12539_ _12554_/CLK _12539_/D vssd1 vssd1 vccd1 vccd1 _12539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10613__B _10613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06810__C _07947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _10645_/A vssd1 vssd1 vccd1 vccd1 _09750_/X sky130_fd_sc_hd__buf_6
X_06962_ _06974_/A vssd1 vssd1 vccd1 vccd1 _06972_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_140_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08701_ _13588_/A vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09690__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09681_ _09681_/A vssd1 vssd1 vccd1 vccd1 _12347_/D sky130_fd_sc_hd__clkbuf_1
X_06893_ _07371_/A vssd1 vssd1 vccd1 vccd1 _07328_/A sky130_fd_sc_hd__buf_2
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08632_ _13586_/A vssd1 vssd1 vccd1 vccd1 _08632_/X sky130_fd_sc_hd__buf_2
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06819__A _06983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13241__397 vssd1 vssd1 vccd1 vccd1 _13241__397/HI _13896_/A sky130_fd_sc_hd__conb_1
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08563_ _13587_/A vssd1 vssd1 vccd1 vccd1 _08563_/X sky130_fd_sc_hd__buf_2
XFILLER_120_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13940__A _13940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07514_ _07514_/A vssd1 vssd1 vccd1 vccd1 _07514_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _12264_/Q vssd1 vssd1 vccd1 vccd1 _09362_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07445_ _07454_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07446_/A sky130_fd_sc_hd__or2_1
X_13094__250 vssd1 vssd1 vccd1 vccd1 _13094__250/HI _13603_/A sky130_fd_sc_hd__conb_1
XANTENNA__09849__B _13562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07376_ _07403_/A vssd1 vssd1 vccd1 vccd1 _07388_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_148_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09115_ peripheralBus_data[14] vssd1 vssd1 vccd1 vccd1 _10548_/A sky130_fd_sc_hd__buf_4
X_06327_ _06333_/A _06336_/B _06336_/C vssd1 vssd1 vccd1 vccd1 _06328_/A sky130_fd_sc_hd__or3_1
XANTENNA__09270__A1 _09347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135__291 vssd1 vssd1 vccd1 vccd1 _13135__291/HI _13676_/A sky130_fd_sc_hd__conb_1
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09046_ _12844_/Q _12845_/Q _12846_/Q _12847_/Q _08967_/X _08968_/X vssd1 vssd1 vccd1
+ vccd1 _09046_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07385__A _07964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09948_ _10700_/A _09948_/B vssd1 vssd1 vccd1 vccd1 _09949_/A sky130_fd_sc_hd__or2_1
X_09879_ _09124_/X _09874_/X _09877_/X _09878_/X vssd1 vssd1 vccd1 vccd1 _12391_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11910_ _11910_/A _11910_/B _11910_/C _11910_/D vssd1 vssd1 vccd1 vccd1 _11921_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _12895_/CLK _12890_/D vssd1 vssd1 vccd1 vccd1 _12890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06729__A _06729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__A input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11841_ _11852_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _11842_/A sky130_fd_sc_hd__and2_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999__155 vssd1 vssd1 vccd1 vccd1 _12999__155/HI _13410_/A sky130_fd_sc_hd__conb_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11772_ _12860_/Q _13365_/A vssd1 vssd1 vccd1 vccd1 _11775_/B sky130_fd_sc_hd__xor2_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13511_/A _07592_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11840__A0 peripheralBus_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _13976_/Z _13784_/A _10723_/S vssd1 vssd1 vccd1 vccd1 _10724_/B sky130_fd_sc_hd__mux2_1
XFILLER_158_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13442_ _13442_/A _07773_/X vssd1 vssd1 vccd1 vccd1 _13666_/Z sky130_fd_sc_hd__ebufn_8
X_10654_ _10652_/X _10638_/X _10653_/X _10650_/X vssd1 vssd1 vccd1 vccd1 _12588_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06464__A _06729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13373_ _13373_/A _08310_/X vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__ebufn_8
X_10585_ _10585_/A _10585_/B vssd1 vssd1 vccd1 vccd1 _10586_/A sky130_fd_sc_hd__and2_1
XFILLER_126_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12324_ _12367_/CLK _12324_/D vssd1 vssd1 vccd1 vccd1 _13569_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_127_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12255_ _12258_/CLK _12255_/D vssd1 vssd1 vccd1 vccd1 _12255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11206_ _11206_/A vssd1 vssd1 vccd1 vccd1 _11221_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12186_ _14097_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12186_/X sky130_fd_sc_hd__or2_1
X_11137_ _12697_/Q _13938_/A vssd1 vssd1 vccd1 vccd1 _11138_/D sky130_fd_sc_hd__xor2_1
XFILLER_95_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output57_A _13570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ _11195_/A vssd1 vssd1 vccd1 vccd1 _11068_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10019_ _10024_/C _10062_/B _10019_/C vssd1 vssd1 vccd1 vccd1 _10020_/A sky130_fd_sc_hd__and3b_1
XFILLER_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06639__A _11924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11264__B _13945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13078__234 vssd1 vssd1 vccd1 vccd1 _13078__234/HI _13573_/A sky130_fd_sc_hd__conb_1
XANTENNA__13760__A _13760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13709_ _13709_/A _07067_/X vssd1 vssd1 vccd1 vccd1 _14125_/Z sky130_fd_sc_hd__ebufn_8
X_07230_ _07230_/A vssd1 vssd1 vccd1 vccd1 _07246_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13119__275 vssd1 vssd1 vccd1 vccd1 _13119__275/HI _13644_/A sky130_fd_sc_hd__conb_1
X_07161_ _07161_/A vssd1 vssd1 vccd1 vccd1 _07161_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07092_ _07092_/A vssd1 vssd1 vccd1 vccd1 _07092_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13935__A _13935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ _09836_/A vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09960__C1 _09959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07994_ _07994_/A vssd1 vssd1 vccd1 vccd1 _07994_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_141_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07933__A _11154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ _12349_/Q _13559_/A vssd1 vssd1 vccd1 vccd1 _09735_/C sky130_fd_sc_hd__xor2_1
X_06945_ _06945_/A vssd1 vssd1 vccd1 vccd1 _06945_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11455__A _11680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09664_ _09664_/A vssd1 vssd1 vccd1 vccd1 _12342_/D sky130_fd_sc_hd__clkbuf_1
X_06876_ _06876_/A vssd1 vssd1 vccd1 vccd1 _06876_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08610__S0 _08575_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08615_ _10099_/D _12444_/Q _12445_/Q _10098_/B _08553_/X _08554_/X vssd1 vssd1 vccd1
+ vccd1 _08615_/X sky130_fd_sc_hd__mux4_1
X_09595_ _12311_/Q _13554_/A vssd1 vssd1 vccd1 vccd1 _09597_/C sky130_fd_sc_hd__xor2_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _11708_/D vssd1 vssd1 vccd1 vccd1 _13374_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_24_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08477_ _08474_/X _08476_/X _13396_/A vssd1 vssd1 vccd1 vccd1 _11705_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11902__B _13370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07428_ _07430_/A _07435_/B vssd1 vssd1 vccd1 vccd1 _07429_/A sky130_fd_sc_hd__or2_1
XANTENNA__06284__A _06694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07359_ _07369_/A _07364_/B _07361_/C vssd1 vssd1 vccd1 vccd1 _07360_/A sky130_fd_sc_hd__or3_1
XFILLER_136_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11050__A1 _10665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10370_ _12506_/Q _13748_/A vssd1 vssd1 vccd1 vccd1 _10372_/C sky130_fd_sc_hd__xor2_1
XFILLER_156_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09029_ _10938_/C vssd1 vssd1 vccd1 vccd1 _13941_/A sky130_fd_sc_hd__buf_6
XFILLER_2_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12040_ _12040_/A _12040_/B _12040_/C _12040_/D vssd1 vssd1 vccd1 vccd1 _12057_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08004__A _08004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13991_ _13991_/A _06309_/X vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12942_ _12946_/CLK _12942_/D vssd1 vssd1 vccd1 vccd1 _14068_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06459__A _08276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _12873_/CLK _12873_/D vssd1 vssd1 vccd1 vccd1 _14001_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _11834_/A _11824_/B vssd1 vssd1 vccd1 vccd1 _11825_/A sky130_fd_sc_hd__and2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11755_/A vssd1 vssd1 vccd1 vccd1 _12866_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10706_ _10706_/A vssd1 vssd1 vccd1 vccd1 _10723_/S sky130_fd_sc_hd__clkbuf_2
X_11686_ _11687_/B _11680_/X _11687_/A vssd1 vssd1 vccd1 vccd1 _11690_/B sky130_fd_sc_hd__a21o_1
X_13425_ _13425_/A _07819_/X vssd1 vssd1 vccd1 vccd1 _14033_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_127_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10637_ _10637_/A _10637_/B vssd1 vssd1 vccd1 vccd1 _10673_/A sky130_fd_sc_hd__or2_2
XFILLER_155_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10568_ _10568_/A vssd1 vssd1 vccd1 vccd1 _12570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ _12325_/CLK _12307_/D vssd1 vssd1 vccd1 vccd1 _13438_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10499_ _10499_/A _10499_/B _10499_/C _10499_/D vssd1 vssd1 vccd1 vccd1 _10505_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_46_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12238_ _12242_/CLK _12238_/D vssd1 vssd1 vccd1 vccd1 _12238_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13755__A _13755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ _12960_/Q _13366_/A vssd1 vssd1 vccd1 vccd1 _12171_/C sky130_fd_sc_hd__xor2_1
XFILLER_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 peripheralBus_address[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_06730_ _06730_/A vssd1 vssd1 vccd1 vccd1 _06730_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06661_ _06675_/A vssd1 vssd1 vccd1 vccd1 _06673_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08400_ _12237_/Q _09258_/D _12239_/Q _12240_/Q _08396_/X _08397_/X vssd1 vssd1 vccd1
+ vccd1 _08400_/X sky130_fd_sc_hd__mux4_2
X_09380_ _09380_/A _09380_/B _09380_/C vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__and3_1
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06592_ _06633_/A vssd1 vssd1 vccd1 vccd1 _06602_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ _08336_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08332_/A sky130_fd_sc_hd__or2_1
X_08262_ _08262_/A vssd1 vssd1 vccd1 vccd1 _08262_/X sky130_fd_sc_hd__clkbuf_1
X_07213_ _07220_/A _07216_/B _07213_/C vssd1 vssd1 vccd1 vccd1 _07214_/A sky130_fd_sc_hd__or3_1
X_08193_ _08198_/A _08195_/B _08198_/C vssd1 vssd1 vccd1 vccd1 _08194_/A sky130_fd_sc_hd__or3_1
X_07144_ _07162_/A vssd1 vssd1 vccd1 vccd1 _07160_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07075_ _07090_/A vssd1 vssd1 vccd1 vccd1 _07088_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_145_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09862__B _13558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07977_ _08075_/A _08075_/B _07977_/C vssd1 vssd1 vccd1 vccd1 _07978_/A sky130_fd_sc_hd__or3_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11185__A _11185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ _12352_/Q _13562_/A vssd1 vssd1 vccd1 vccd1 _09716_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06928_ _06928_/A vssd1 vssd1 vccd1 vccd1 _06928_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09647_ _09846_/A vssd1 vssd1 vccd1 vccd1 _10667_/A sky130_fd_sc_hd__buf_4
XFILLER_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06859_ _06900_/A vssd1 vssd1 vccd1 vccd1 _06870_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _13469_/A _12322_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09579_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08529_ _11708_/A vssd1 vssd1 vccd1 vccd1 _13371_/A sky130_fd_sc_hd__buf_4
XANTENNA__11124__S _11124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09102__B _12062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ _11582_/C vssd1 vssd1 vccd1 vccd1 _11540_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11471_ _14066_/Z _09030_/X _11499_/B vssd1 vssd1 vccd1 vccd1 _11472_/B sky130_fd_sc_hd__mux2_1
XFILLER_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10422_ _09116_/X _10409_/X _10421_/X _10412_/X vssd1 vssd1 vccd1 vccd1 _12532_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10353_ _12512_/Q _10613_/B vssd1 vssd1 vccd1 vccd1 _10353_/X sky130_fd_sc_hd__and2_1
XANTENNA__10264__A _10278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10782__B1 _10781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ _09186_/X _10278_/X _10282_/X _10283_/X vssd1 vssd1 vccd1 vccd1 _12496_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11326__A2 _11312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12023_ _12932_/Q _14075_/A _12029_/S vssd1 vssd1 vccd1 vccd1 _12024_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08822__S0 _08807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13974_ _13974_/A _06356_/X vssd1 vssd1 vccd1 vccd1 _13974_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_46_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12925_ _12929_/CLK _12925_/D vssd1 vssd1 vccd1 vccd1 _12925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _12873_/CLK _12856_/D vssd1 vssd1 vccd1 vccd1 _12856_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13040__196 vssd1 vssd1 vccd1 vccd1 _13040__196/HI _13483_/A sky130_fd_sc_hd__conb_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11807_/A vssd1 vssd1 vccd1 vccd1 _12875_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _12923_/CLK _12787_/D vssd1 vssd1 vccd1 vccd1 _13913_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _11738_/A vssd1 vssd1 vccd1 vccd1 _12861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11669_ _11669_/A vssd1 vssd1 vccd1 vccd1 _12844_/D sky130_fd_sc_hd__clkbuf_1
X_13408_ _13408_/A _08098_/X vssd1 vssd1 vccd1 vccd1 _14112_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_127_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06371__B _07822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09963__A _13596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07900_ _07900_/A vssd1 vssd1 vccd1 vccd1 _07900_/X sky130_fd_sc_hd__clkbuf_1
X_08880_ _08822_/X _08825_/X _08855_/X _08879_/X _08810_/X _08876_/X vssd1 vssd1 vccd1
+ vccd1 _08880_/X sky130_fd_sc_hd__mux4_1
X_07831_ _08166_/A vssd1 vssd1 vccd1 vccd1 _08335_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_111_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10621__B _13757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07762_ _07762_/A vssd1 vssd1 vccd1 vccd1 _07762_/X sky130_fd_sc_hd__clkbuf_1
X_09501_ _09526_/B vssd1 vssd1 vccd1 vccd1 _09511_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06713_ _06713_/A vssd1 vssd1 vccd1 vccd1 _06713_/X sky130_fd_sc_hd__clkbuf_1
X_07693_ _07693_/A vssd1 vssd1 vccd1 vccd1 _07704_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09432_ _09439_/A _09432_/B vssd1 vssd1 vccd1 vccd1 _09433_/A sky130_fd_sc_hd__and2_1
X_06644_ _06646_/A _06651_/B _06651_/C vssd1 vssd1 vccd1 vccd1 _06645_/A sky130_fd_sc_hd__or3_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09363_ _09363_/A _09368_/C _09368_/D vssd1 vssd1 vccd1 vccd1 _09364_/B sky130_fd_sc_hd__and3_1
X_06575_ _06575_/A vssd1 vssd1 vccd1 vccd1 _06575_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08314_ _08314_/A vssd1 vssd1 vccd1 vccd1 _08324_/A sky130_fd_sc_hd__clkbuf_4
X_09294_ _09300_/C _09389_/A _09294_/C vssd1 vssd1 vccd1 vccd1 _09295_/A sky130_fd_sc_hd__and3b_1
XFILLER_20_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08245_ _08245_/A vssd1 vssd1 vccd1 vccd1 _08245_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09857__B _13565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08176_ _10693_/A vssd1 vssd1 vccd1 vccd1 _08358_/A sky130_fd_sc_hd__buf_2
XFILLER_146_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07127_ _07127_/A vssd1 vssd1 vccd1 vccd1 _07127_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10084__A _10146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09873__A _11412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ _07058_/A vssd1 vssd1 vccd1 vccd1 _07058_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07393__A _07393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10819__A1 _10885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _10971_/A vssd1 vssd1 vccd1 vccd1 _10986_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12710_ _12710_/CLK _12710_/D vssd1 vssd1 vccd1 vccd1 _13953_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__07840__B _07840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13690_ _13690_/A _07119_/X vssd1 vssd1 vccd1 vccd1 _14106_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_71_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12641_ _12813_/CLK _12641_/D vssd1 vssd1 vccd1 vccd1 _12641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_16_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ _12598_/CLK _12572_/D vssd1 vssd1 vccd1 vccd1 _12572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11523_ _11523_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _12810_/D sky130_fd_sc_hd__nor2_1
XFILLER_156_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06472__A _06481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11454_ _13967_/A vssd1 vssd1 vccd1 vccd1 _11680_/A sky130_fd_sc_hd__buf_2
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10405_ _09770_/X _10395_/X _10404_/X _10398_/X vssd1 vssd1 vccd1 vccd1 _12526_/D
+ sky130_fd_sc_hd__o211a_1
X_11385_ _12773_/Q _11386_/B vssd1 vssd1 vccd1 vccd1 _11385_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10336_ _13658_/A _12512_/Q _10342_/S vssd1 vssd1 vccd1 vccd1 _10337_/B sky130_fd_sc_hd__mux2_1
XFILLER_152_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11818__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_clk clkbuf_4_9_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clk/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater110_A peripheralBus_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _09160_/X _10264_/X _10266_/X _10256_/X vssd1 vssd1 vccd1 vccd1 _12490_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10722__A input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12006_ _12927_/Q _14070_/A _12012_/S vssd1 vssd1 vccd1 vccd1 _12007_/B sky130_fd_sc_hd__mux2_1
Xrepeater108 _14096_/Z vssd1 vssd1 vccd1 vccd1 _14064_/Z sky130_fd_sc_hd__buf_12
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10198_ _10208_/A _10198_/B vssd1 vssd1 vccd1 vccd1 _10199_/A sky130_fd_sc_hd__and2_1
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater119 peripheralBus_data[16] vssd1 vssd1 vccd1 vccd1 _14111_/Z sky130_fd_sc_hd__buf_12
XFILLER_120_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13957_ _13957_/A _06404_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12908_ _12908_/CLK _12908_/D vssd1 vssd1 vccd1 vccd1 _14035_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13888_ _13888_/A _06590_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[17] sky130_fd_sc_hd__ebufn_8
XANTENNA__11272__B _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12839_ _12842_/CLK _12839_/D vssd1 vssd1 vccd1 vccd1 _12839_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09958__A _13594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06360_ _06360_/A vssd1 vssd1 vccd1 vccd1 _06360_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06291_ _06303_/A _07845_/A _07979_/A vssd1 vssd1 vccd1 vccd1 _06292_/A sky130_fd_sc_hd__or3_1
X_08030_ _08039_/A _08033_/B _08030_/C vssd1 vssd1 vccd1 vccd1 _08031_/A sky130_fd_sc_hd__or3_1
XFILLER_163_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10616__B _13756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06813__C _09097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09981_ _09981_/A _09981_/B _12422_/Q _12421_/Q vssd1 vssd1 vccd1 vccd1 _10030_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_103_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08932_ _12831_/Q _12832_/Q _12833_/Q _12834_/Q _08921_/X _08922_/X vssd1 vssd1 vccd1
+ vccd1 _08932_/X sky130_fd_sc_hd__mux4_2
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08863_ _08860_/X _08862_/X _08863_/S vssd1 vssd1 vccd1 vccd1 _10164_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10351__B _13752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13943__A _13943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07814_ _07814_/A vssd1 vssd1 vccd1 vccd1 _07814_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08794_ _12647_/Q vssd1 vssd1 vccd1 vccd1 _10908_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07745_ _07798_/A vssd1 vssd1 vccd1 vccd1 _07756_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11463__A _14063_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07676_ _07686_/A _07683_/B _07678_/C vssd1 vssd1 vccd1 vccd1 _07677_/A sky130_fd_sc_hd__or3_1
X_09415_ _09422_/A _09415_/B vssd1 vssd1 vccd1 vccd1 _09416_/A sky130_fd_sc_hd__and2_1
XFILLER_53_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06627_ _06675_/A vssd1 vssd1 vccd1 vccd1 _06646_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09346_ _09352_/B _09352_/C _09346_/C vssd1 vssd1 vccd1 vccd1 _09368_/C sky130_fd_sc_hd__and3_1
X_06558_ _06599_/A vssd1 vssd1 vccd1 vccd1 _06569_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09587__B _09848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09277_ _09284_/D _09276_/C _09321_/C vssd1 vssd1 vccd1 vccd1 _09278_/C sky130_fd_sc_hd__a21o_1
X_06489_ _08276_/B vssd1 vssd1 vccd1 vccd1 _06499_/C sky130_fd_sc_hd__clkbuf_1
X_08228_ _08228_/A vssd1 vssd1 vccd1 vccd1 _08238_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_165_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08159_ _08177_/A vssd1 vssd1 vccd1 vccd1 _08174_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_106_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11170_ _11170_/A vssd1 vssd1 vccd1 vccd1 _11170_/X sky130_fd_sc_hd__buf_6
X_10121_ _12457_/Q vssd1 vssd1 vccd1 vccd1 _10130_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07835__B _07840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10052_ _10052_/A _10052_/B _10052_/C _10052_/D vssd1 vssd1 vccd1 vccd1 _10100_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__09108__A _11443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08012__A _08186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13811_ _13811_/A _06802_/X vssd1 vssd1 vccd1 vccd1 _14067_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA_input19_A peripheralBus_address[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13742_ _13742_/A _06988_/X vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11465__A1 _11689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ _10971_/A vssd1 vssd1 vccd1 vccd1 _10969_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13673_ _13673_/A _07164_/X vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_44_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10885_ _10885_/A _10908_/C _10922_/B vssd1 vssd1 vccd1 vccd1 _10891_/B sky130_fd_sc_hd__and3_1
X_12624_ _12625_/CLK _12624_/D vssd1 vssd1 vccd1 vccd1 _12624_/Q sky130_fd_sc_hd__dfxtp_1
X_12555_ _12555_/CLK _12555_/D vssd1 vssd1 vccd1 vccd1 _13683_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ _11506_/A vssd1 vssd1 vccd1 vccd1 _12807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12486_ _12492_/CLK _12486_/D vssd1 vssd1 vccd1 vccd1 _13616_/A sky130_fd_sc_hd__dfxtp_1
X_11437_ _10670_/X _11425_/X _11436_/X _11430_/X vssd1 vssd1 vccd1 vccd1 _12786_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ _11377_/A _11368_/B vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__and2_1
XFILLER_140_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _10332_/A _10319_/B vssd1 vssd1 vccd1 vccd1 _10320_/A sky130_fd_sc_hd__and2_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14087_/A _08058_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_113_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11299_ _11312_/A vssd1 vssd1 vccd1 vccd1 _11299_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11267__B _13938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09897__A1 _09767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07530_ _07530_/A vssd1 vssd1 vccd1 vccd1 _07530_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06377__A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07461_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07471_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_62_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352__508 vssd1 vssd1 vccd1 vccd1 _13352__508/HI _14121_/A sky130_fd_sc_hd__conb_1
X_09200_ _09200_/A vssd1 vssd1 vccd1 vccd1 _12228_/D sky130_fd_sc_hd__clkbuf_1
X_06412_ _06416_/A _06412_/B vssd1 vssd1 vccd1 vccd1 _06413_/A sky130_fd_sc_hd__or2_1
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09688__A _09967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07392_ _07392_/A vssd1 vssd1 vccd1 vccd1 _07392_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09131_ _13391_/A vssd1 vssd1 vccd1 vccd1 _09269_/A sky130_fd_sc_hd__buf_2
X_06343_ _06343_/A vssd1 vssd1 vccd1 vccd1 _06343_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09062_ _09004_/X _09008_/X _09036_/X _09061_/X _09056_/X _08996_/X vssd1 vssd1 vccd1
+ vccd1 _09062_/X sky130_fd_sc_hd__mux4_1
X_06274_ input4/X _09097_/B _09097_/C vssd1 vssd1 vccd1 vccd1 _07319_/C sky130_fd_sc_hd__or3_1
XFILLER_135_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08013_ _08067_/A vssd1 vssd1 vccd1 vccd1 _08025_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__13938__A _13938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10719__A0 _14103_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13246__402 vssd1 vssd1 vccd1 vccd1 _13246__402/HI _13901_/A sky130_fd_sc_hd__conb_1
XFILLER_143_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09964_ _09112_/X _09934_/S _09963_/X _09959_/X vssd1 vssd1 vccd1 vccd1 _12420_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09337__B1 _09236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08915_ _13968_/A vssd1 vssd1 vccd1 vccd1 _08915_/X sky130_fd_sc_hd__clkbuf_4
X_09895_ _09763_/X _09888_/X _09894_/X _09892_/X vssd1 vssd1 vccd1 vccd1 _12397_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _12648_/Q _10907_/D _12650_/Q _12651_/Q _08739_/X _08740_/X vssd1 vssd1 vccd1
+ vccd1 _08846_/X sky130_fd_sc_hd__mux4_2
XANTENNA__08767__A _13777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _10163_/B vssd1 vssd1 vccd1 vccd1 _10614_/B sky130_fd_sc_hd__buf_2
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11447__A1 _11061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _07728_/A vssd1 vssd1 vccd1 vccd1 _07728_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07659_ _07659_/A _07669_/B _07664_/C vssd1 vssd1 vccd1 vccd1 _07660_/A sky130_fd_sc_hd__or3_1
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10670_ _10670_/A vssd1 vssd1 vccd1 vccd1 _10670_/X sky130_fd_sc_hd__buf_6
XFILLER_159_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ _09329_/A _09329_/B _09329_/C vssd1 vssd1 vccd1 vccd1 _09331_/C sky130_fd_sc_hd__and3_1
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ _12340_/CLK _12340_/D vssd1 vssd1 vccd1 vccd1 _13470_/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__08007__A _08022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12271_ _12274_/CLK _12271_/D vssd1 vssd1 vccd1 vccd1 _12271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _14010_/A _08136_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[11] sky130_fd_sc_hd__ebufn_8
X_11222_ _11222_/A vssd1 vssd1 vccd1 vccd1 _12732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11153_ _11153_/A vssd1 vssd1 vccd1 vccd1 _11153_/X sky130_fd_sc_hd__buf_4
X_10104_ _10133_/B _10135_/B _10104_/C vssd1 vssd1 vccd1 vccd1 _10105_/A sky130_fd_sc_hd__and3b_1
XFILLER_49_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11084_ _13842_/A _12697_/Q _11151_/B vssd1 vssd1 vccd1 vccd1 _11085_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09879__A1 _09124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ _10097_/C _10089_/A _09978_/X vssd1 vssd1 vccd1 vccd1 _10035_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13583__A _13583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ _12921_/Q _14064_/A _11995_/S vssd1 vssd1 vccd1 vccd1 _11987_/B sky130_fd_sc_hd__mux2_1
X_13725_ _13725_/A _07028_/X vssd1 vssd1 vccd1 vccd1 _14077_/Z sky130_fd_sc_hd__ebufn_8
X_10937_ _10937_/A vssd1 vssd1 vccd1 vccd1 _12660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11831__A _11834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13656_ _13656_/A _07210_/X vssd1 vssd1 vccd1 vccd1 _14072_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06925__A _07480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10868_ _10874_/A _10875_/A _10876_/A _10868_/D vssd1 vssd1 vccd1 vccd1 _10871_/B
+ sky130_fd_sc_hd__and4_1
X_12607_ _12811_/CLK _12607_/D vssd1 vssd1 vccd1 vccd1 _13782_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11550__B _11604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09264__C1 _09263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ _13587_/A _07400_/X vssd1 vssd1 vccd1 vccd1 _14035_/Z sky130_fd_sc_hd__ebufn_8
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _10863_/A _10800_/B _10798_/X vssd1 vssd1 vccd1 vccd1 _10801_/A sky130_fd_sc_hd__o21ai_1
X_12538_ _12554_/CLK _12538_/D vssd1 vssd1 vccd1 vccd1 _12538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13758__A _13758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12469_ _12492_/CLK _12469_/D vssd1 vssd1 vccd1 vccd1 _12469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06961_ _06961_/A vssd1 vssd1 vccd1 vccd1 _06961_/X sky130_fd_sc_hd__clkbuf_1
X_08700_ _08643_/X _08646_/X _08674_/X _08699_/X _08694_/X _08695_/X vssd1 vssd1 vccd1
+ vccd1 _08700_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13493__A _13493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09680_ _09686_/A _09680_/B vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__and2_1
X_06892_ _09125_/A vssd1 vssd1 vccd1 vccd1 _07371_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08631_ _10029_/A _12437_/Q _10097_/B _12439_/Q _08629_/X _08630_/X vssd1 vssd1 vccd1
+ vccd1 _08631_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08562_ _13586_/A vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__clkbuf_2
X_07513_ _07517_/A _07517_/B _07524_/C vssd1 vssd1 vccd1 vccd1 _07514_/A sky130_fd_sc_hd__or3_1
X_08493_ _08378_/X _08381_/X _08386_/X _08388_/X _08492_/X _08424_/X vssd1 vssd1 vccd1
+ vccd1 _08493_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07444_ _07468_/A vssd1 vssd1 vccd1 vccd1 _07454_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09211__A _09347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__B _11460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07375_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07375_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09114_ _09112_/X _09100_/X _09113_/X _09109_/X vssd1 vssd1 vccd1 vccd1 _12211_/D
+ sky130_fd_sc_hd__o211a_1
X_06326_ _07045_/A vssd1 vssd1 vccd1 vccd1 _06336_/C sky130_fd_sc_hd__clkbuf_1
X_09045_ _08950_/X _08951_/X _08955_/X _08957_/X _09030_/A _08934_/X vssd1 vssd1 vccd1
+ vccd1 _09045_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09865__B _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09947_ _14102_/Z _13590_/A _09953_/S vssd1 vssd1 vccd1 vccd1 _09948_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09878_ _09878_/A vssd1 vssd1 vccd1 vccd1 _09878_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08829_ _08813_/X _08827_/X _08890_/S vssd1 vssd1 vccd1 vccd1 _10163_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06729__B _07323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ peripheralBus_data[14] _14013_/A _11840_/S vssd1 vssd1 vccd1 vccd1 _11841_/B
+ sky130_fd_sc_hd__mux2_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12093__A1 _11189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11771_ _12857_/Q _13362_/A vssd1 vssd1 vccd1 vccd1 _11775_/A sky130_fd_sc_hd__xor2_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11651__A _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ _13510_/A _07594_/X vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_8
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ input27/X vssd1 vssd1 vccd1 vccd1 _11481_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13441_ _13441_/A _07775_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_70_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10653_ _13715_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10653_/X sky130_fd_sc_hd__or2_1
X_13372_ _13372_/A _08308_/X vssd1 vssd1 vccd1 vccd1 _14108_/Z sky130_fd_sc_hd__ebufn_8
X_10584_ _13719_/A _12575_/Q _10584_/S vssd1 vssd1 vccd1 vccd1 _10585_/B sky130_fd_sc_hd__mux2_1
X_12323_ _12349_/CLK _12323_/D vssd1 vssd1 vccd1 vccd1 _12323_/Q sky130_fd_sc_hd__dfxtp_1
X_12254_ _12258_/CLK _12254_/D vssd1 vssd1 vccd1 vccd1 _12254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11205_ _11205_/A vssd1 vssd1 vccd1 vccd1 _12727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12185_ _11160_/X _12182_/X _12184_/X _12097_/X vssd1 vssd1 vccd1 vccd1 _12971_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09791__A _13593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11136_ _12700_/Q _13941_/A vssd1 vssd1 vccd1 vccd1 _11138_/C sky130_fd_sc_hd__xor2_1
XFILLER_150_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11067_ _13821_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11067_/X sky130_fd_sc_hd__or2_1
XANTENNA__10730__A _13787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10018_ _10021_/C _10016_/C _10021_/B vssd1 vssd1 vccd1 vccd1 _10019_/C sky130_fd_sc_hd__a21o_1
XFILLER_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08200__A _08240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11969_ _11978_/A _11969_/B vssd1 vssd1 vccd1 vccd1 _11970_/A sky130_fd_sc_hd__and2_1
XFILLER_60_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13708_ _13708_/A _07070_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_32_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13639_ _13639_/A _07257_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07160_ _07166_/A _07163_/B _07160_/C vssd1 vssd1 vccd1 vccd1 _07161_/A sky130_fd_sc_hd__or3_1
XFILLER_9_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07091_ _07094_/A _07091_/B _07101_/C vssd1 vssd1 vccd1 vccd1 _07092_/A sky130_fd_sc_hd__or3_1
XFILLER_118_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07486__A _08089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06390__A _07845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10624__B _13755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09801_ _09801_/A vssd1 vssd1 vccd1 vccd1 _12376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07993_ _07997_/A _08062_/B _07993_/C vssd1 vssd1 vccd1 vccd1 _07994_/A sky130_fd_sc_hd__or3_1
X_09732_ _12346_/Q _13556_/A vssd1 vssd1 vccd1 vccd1 _09735_/B sky130_fd_sc_hd__xor2_1
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06944_ _06948_/A _06953_/B vssd1 vssd1 vccd1 vccd1 _06945_/A sky130_fd_sc_hd__or2_1
XANTENNA__10640__A _10686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater72_A _14100_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _09669_/A _09663_/B vssd1 vssd1 vccd1 vccd1 _09664_/A sky130_fd_sc_hd__and2_1
XFILLER_28_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13358__514 vssd1 vssd1 vccd1 vccd1 _13358__514/HI peripheralBus_busy sky130_fd_sc_hd__conb_1
XANTENNA__08110__A _08110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ _06877_/A _06884_/B _06884_/C vssd1 vssd1 vccd1 vccd1 _06876_/A sky130_fd_sc_hd__or3_1
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08610__S1 _08576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13951__A _13951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ _12439_/Q _12440_/Q _12441_/Q _10052_/A _08578_/X _08579_/X vssd1 vssd1 vccd1
+ vccd1 _08614_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09594_ _12314_/Q _13557_/A vssd1 vssd1 vccd1 vccd1 _09597_/B sky130_fd_sc_hd__xor2_1
XFILLER_43_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _08541_/X _08544_/X _09162_/A vssd1 vssd1 vccd1 vccd1 _11708_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _08407_/X _08409_/X _08411_/X _08475_/X _08479_/A _08383_/X vssd1 vssd1 vccd1
+ vccd1 _08476_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ _07427_/A vssd1 vssd1 vccd1 vccd1 _07427_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09876__A _09915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07358_ _07371_/A vssd1 vssd1 vccd1 vccd1 _07369_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__10389__A1 _09750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11586__B1 _11540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06309_ _06309_/A vssd1 vssd1 vccd1 vccd1 _06309_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09595__B _13554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07289_ _07292_/A _07289_/B _07300_/C vssd1 vssd1 vccd1 vccd1 _07290_/A sky130_fd_sc_hd__or3_1
XFILLER_163_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09028_ _09025_/X _09027_/X _09043_/S vssd1 vssd1 vccd1 vccd1 _10938_/C sky130_fd_sc_hd__mux2_2
XFILLER_124_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07827__C _08349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07843__B _07854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10550__A _10650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ _13990_/A _06315_/X vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_93_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08506__A1 _08423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09116__A _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ _12946_/CLK _12941_/D vssd1 vssd1 vccd1 vccd1 _14067_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12872_ _12873_/CLK _12872_/D vssd1 vssd1 vccd1 vccd1 _14000_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11823_ _09638_/A _14008_/A _11823_/S vssd1 vssd1 vccd1 vccd1 _11824_/B sky130_fd_sc_hd__mux2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11757_/A _11754_/B vssd1 vssd1 vccd1 vccd1 _11755_/A sky130_fd_sc_hd__and2_1
XFILLER_14_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10705_/A vssd1 vssd1 vccd1 vccd1 _12603_/D sky130_fd_sc_hd__clkbuf_1
X_11685_ _11687_/B _11680_/X _11684_/Y vssd1 vssd1 vccd1 vccd1 _12848_/D sky130_fd_sc_hd__a21oi_1
XFILLER_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13151__307 vssd1 vssd1 vccd1 vccd1 _13151__307/HI _13708_/A sky130_fd_sc_hd__conb_1
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13424_ _13424_/A _07821_/X vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_8
X_10636_ _10636_/A vssd1 vssd1 vccd1 vccd1 _12583_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11577__B1 _11576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10567_ _10567_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _10568_/A sky130_fd_sc_hd__and2_1
XFILLER_154_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12306_ _12969_/CLK _12306_/D vssd1 vssd1 vccd1 vccd1 _13437_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_155_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10498_ _12541_/Q _13750_/A vssd1 vssd1 vccd1 vccd1 _10499_/D sky130_fd_sc_hd__xor2_1
X_12237_ _12242_/CLK _12237_/D vssd1 vssd1 vccd1 vccd1 _12237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12168_ _12968_/Q _13374_/A vssd1 vssd1 vccd1 vccd1 _12171_/B sky130_fd_sc_hd__xor2_1
XFILLER_69_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13045__201 vssd1 vssd1 vccd1 vccd1 _13045__201/HI _13504_/A sky130_fd_sc_hd__conb_1
XFILLER_122_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11556__A _11703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ _11204_/A _11119_/B vssd1 vssd1 vccd1 vccd1 _11120_/A sky130_fd_sc_hd__and2_1
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12099_ _14077_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__or2_1
XANTENNA__11275__B _13935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 peripheralBus_address[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11501__A0 _10939_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06369__B _07822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06660_ _06660_/A vssd1 vssd1 vccd1 vccd1 _06660_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06591_ _06604_/A vssd1 vssd1 vccd1 vccd1 _06602_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ _08330_/A vssd1 vssd1 vccd1 vccd1 _08330_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10619__B _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ _08264_/A _08261_/B _08264_/C vssd1 vssd1 vccd1 vccd1 _08262_/A sky130_fd_sc_hd__or3_1
XFILLER_165_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07212_ _07212_/A vssd1 vssd1 vccd1 vccd1 _07212_/X sky130_fd_sc_hd__clkbuf_1
X_08192_ _08192_/A vssd1 vssd1 vccd1 vccd1 _08192_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07143_ _07143_/A vssd1 vssd1 vccd1 vccd1 _07143_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10635__A _11151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07074_ _07074_/A vssd1 vssd1 vccd1 vccd1 _07074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08105__A _08110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__B _10614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13946__A _13946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10543__A1 _10414_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11466__A _14064_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _07976_/A vssd1 vssd1 vccd1 vccd1 _07976_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09715_ _12352_/Q _09848_/B vssd1 vssd1 vccd1 vccd1 _09715_/X sky130_fd_sc_hd__and2_1
XFILLER_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06927_ _06936_/A _06929_/B vssd1 vssd1 vccd1 vccd1 _06928_/A sky130_fd_sc_hd__or2_1
XFILLER_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08595__S0 _08556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ _11061_/A _09653_/B vssd1 vssd1 vccd1 vccd1 _09646_/X sky130_fd_sc_hd__or2_1
XFILLER_28_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06858_ _06858_/A vssd1 vssd1 vccd1 vccd1 _06858_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11913__B _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _09577_/A vssd1 vssd1 vccd1 vccd1 _12321_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ _06789_/A vssd1 vssd1 vccd1 vccd1 _06789_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08528_ _08522_/X _08527_/X _08528_/S vssd1 vssd1 vccd1 vccd1 _11708_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06295__A _08266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ _12260_/Q vssd1 vssd1 vccd1 vccd1 _09346_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10248__C _10693_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11470_ _11470_/A vssd1 vssd1 vccd1 vccd1 _12795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10421_ _13661_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10421_/X sky130_fd_sc_hd__or2_1
XFILLER_109_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ _12512_/Q _13754_/A vssd1 vssd1 vccd1 vccd1 _10352_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10283_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10283_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07854__A _07857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ _12022_/A vssd1 vssd1 vccd1 vccd1 _12931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10534__A1 _09770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08822__S1 _08808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13973_ _13973_/A _06358_/X vssd1 vssd1 vccd1 vccd1 _13973_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12924_ _12929_/CLK _12924_/D vssd1 vssd1 vccd1 vccd1 _12924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12855_ _12873_/CLK _12855_/D vssd1 vssd1 vccd1 vccd1 _12855_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _11816_/A _11806_/B vssd1 vssd1 vccd1 vccd1 _11807_/A sky130_fd_sc_hd__and2_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11798__A0 _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12786_/CLK _12786_/D vssd1 vssd1 vccd1 vccd1 _13912_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11740_/A _11737_/B vssd1 vssd1 vccd1 vccd1 _11738_/A sky130_fd_sc_hd__and2_1
X_11668_ _11703_/A _11668_/B _11668_/C vssd1 vssd1 vccd1 vccd1 _11669_/A sky130_fd_sc_hd__and3_1
X_13407_ _13407_/A _08086_/X vssd1 vssd1 vccd1 vccd1 _14079_/Z sky130_fd_sc_hd__ebufn_8
X_10619_ _12573_/Q _13749_/A vssd1 vssd1 vccd1 vccd1 _10622_/B sky130_fd_sc_hd__xor2_1
XFILLER_127_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11599_ _11641_/D vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06371__C _07822_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09963__B _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11286__A _11325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ _09125_/B vssd1 vssd1 vccd1 vccd1 _08166_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07761_ _07769_/A _07766_/B _07761_/C vssd1 vssd1 vccd1 vccd1 _07762_/A sky130_fd_sc_hd__or3_1
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09500_ _09513_/A vssd1 vssd1 vccd1 vccd1 _09500_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08577__S0 _08575_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06712_ _06714_/A _06719_/B _06719_/C vssd1 vssd1 vccd1 vccd1 _06713_/A sky130_fd_sc_hd__or3_1
XFILLER_37_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07692_ _07692_/A vssd1 vssd1 vccd1 vccd1 _07692_/X sky130_fd_sc_hd__clkbuf_1
X_13320__476 vssd1 vssd1 vccd1 vccd1 _13320__476/HI _14057_/A sky130_fd_sc_hd__conb_1
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09431_ _13431_/A _12283_/Q _09431_/S vssd1 vssd1 vccd1 vccd1 _09432_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06643_ _06643_/A vssd1 vssd1 vccd1 vccd1 _06643_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09362_ _09362_/A _09362_/B _09362_/C _09362_/D vssd1 vssd1 vccd1 vccd1 _09368_/D
+ sky130_fd_sc_hd__and4_1
X_06574_ _06584_/A _06574_/B _06574_/C vssd1 vssd1 vccd1 vccd1 _06575_/A sky130_fd_sc_hd__or3_1
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08313_ _08313_/A vssd1 vssd1 vccd1 vccd1 _08313_/X sky130_fd_sc_hd__clkbuf_1
X_09293_ _09330_/D _09292_/C _09330_/C vssd1 vssd1 vccd1 vccd1 _09294_/C sky130_fd_sc_hd__a21o_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08244_ _08251_/A _08248_/B _08251_/C vssd1 vssd1 vccd1 vccd1 _08245_/A sky130_fd_sc_hd__or3_1
XFILLER_165_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08175_ _08175_/A vssd1 vssd1 vccd1 vccd1 _08175_/X sky130_fd_sc_hd__clkbuf_1
X_13214__370 vssd1 vssd1 vccd1 vccd1 _13214__370/HI _13837_/A sky130_fd_sc_hd__conb_1
XFILLER_21_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07126_ _07135_/A _07131_/B _07128_/C vssd1 vssd1 vccd1 vccd1 _07127_/A sky130_fd_sc_hd__or3_1
XFILLER_119_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11961__A0 peripheralBus_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07057_ _07979_/A _07979_/B vssd1 vssd1 vccd1 vccd1 _07058_/A sky130_fd_sc_hd__or2_1
XFILLER_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07674__A _07923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11908__B _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07959_ _07959_/A vssd1 vssd1 vccd1 vccd1 _07959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08568__S0 _08559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__A _11924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10970_ _10970_/A vssd1 vssd1 vccd1 vccd1 _12668_/D sky130_fd_sc_hd__clkbuf_1
X_09629_ _11170_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09629_/X sky130_fd_sc_hd__or2_1
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12640_ _12820_/CLK _12640_/D vssd1 vssd1 vccd1 vccd1 _12640_/Q sky130_fd_sc_hd__dfxtp_1
X_12571_ _12589_/CLK _12571_/D vssd1 vssd1 vccd1 vccd1 _12571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _12710_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _11518_/A _11517_/A _11521_/X vssd1 vssd1 vccd1 vccd1 _11523_/B sky130_fd_sc_hd__o21ai_1
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11453_ _10552_/A _11438_/A _11452_/X _11444_/X vssd1 vssd1 vccd1 vccd1 _12792_/D
+ sky130_fd_sc_hd__o211a_1
X_10404_ _13655_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10404_/X sky130_fd_sc_hd__or2_1
XFILLER_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11384_ _12769_/Q _11384_/B vssd1 vssd1 vccd1 vccd1 _11384_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_164_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10335_ _10479_/A vssd1 vssd1 vccd1 vccd1 _10349_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13263__419 vssd1 vssd1 vccd1 vccd1 _13263__419/HI _13934_/A sky130_fd_sc_hd__conb_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10266_ _13620_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10266_/X sky130_fd_sc_hd__or2_1
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12005_ _12005_/A vssd1 vssd1 vccd1 vccd1 _12926_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_repeater103_A peripheralBus_data[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater109 _13616_/Z vssd1 vssd1 vccd1 vccd1 _14096_/Z sky130_fd_sc_hd__buf_12
X_10197_ _13623_/A _12476_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _10198_/B sky130_fd_sc_hd__mux2_1
XFILLER_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11834__A _11834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13956_ _13956_/A _06407_/X vssd1 vssd1 vccd1 vccd1 _13988_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output32_A _13978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12907_ _12919_/CLK _12907_/D vssd1 vssd1 vccd1 vccd1 _14034_/A sky130_fd_sc_hd__dfxtp_1
X_13887_ _13887_/A _06594_/X vssd1 vssd1 vccd1 vccd1 _14079_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13157__313 vssd1 vssd1 vccd1 vccd1 _13157__313/HI _13730_/A sky130_fd_sc_hd__conb_1
X_12838_ _12842_/CLK _12838_/D vssd1 vssd1 vccd1 vccd1 _12838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _12786_/CLK _12769_/D vssd1 vssd1 vccd1 vccd1 _12769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _12586_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06290_ _08364_/A vssd1 vssd1 vccd1 vccd1 _06303_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 peripheralBus_address[5] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09974__A _09977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09980_ _09981_/B _09972_/X _09979_/Y vssd1 vssd1 vccd1 vccd1 _12423_/D sky130_fd_sc_hd__a21oi_1
XFILLER_89_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08931_ _12827_/Q _12828_/Q _12829_/Q _12830_/Q _08928_/X _08929_/X vssd1 vssd1 vccd1
+ vccd1 _08931_/X sky130_fd_sc_hd__mux4_2
XFILLER_130_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08862_ _08756_/X _08757_/X _08833_/X _08861_/X _08748_/X _08749_/X vssd1 vssd1 vccd1
+ vccd1 _08862_/X sky130_fd_sc_hd__mux4_1
X_07813_ _07868_/A _07820_/B _07815_/C vssd1 vssd1 vccd1 vccd1 _07814_/A sky130_fd_sc_hd__or3_1
XFILLER_85_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08793_ _10876_/B _12641_/Q _12642_/Q _10874_/A _08785_/X _08786_/X vssd1 vssd1 vccd1
+ vccd1 _08793_/X sky130_fd_sc_hd__mux4_2
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07744_ _07923_/A vssd1 vssd1 vccd1 vccd1 _07798_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07675_ _07729_/A vssd1 vssd1 vccd1 vccd1 _07686_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09414_ _13426_/A _12278_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _09415_/B sky130_fd_sc_hd__mux2_1
XFILLER_13_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08970__S0 _08967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06626_ _06626_/A vssd1 vssd1 vccd1 vccd1 _06626_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09345_ _09352_/C _09352_/D _09344_/Y _09263_/X vssd1 vssd1 vccd1 vccd1 _12261_/D
+ sky130_fd_sc_hd__o211a_1
X_06557_ _06557_/A vssd1 vssd1 vccd1 vccd1 _06557_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_32_clk _12759_/CLK vssd1 vssd1 vccd1 vccd1 _12782_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09276_ _09321_/C _09284_/D _09276_/C vssd1 vssd1 vccd1 vccd1 _09276_/X sky130_fd_sc_hd__and3_1
X_06488_ _06528_/A vssd1 vssd1 vccd1 vccd1 _06499_/B sky130_fd_sc_hd__clkbuf_1
X_08227_ _08240_/A vssd1 vssd1 vccd1 vccd1 _08238_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__10095__A _10146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08158_ _10693_/A vssd1 vssd1 vccd1 vccd1 _08174_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11934__A0 _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ _07109_/A vssd1 vssd1 vccd1 vccd1 _07109_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08089_ _08089_/A _08089_/B vssd1 vssd1 vccd1 vccd1 _08090_/A sky130_fd_sc_hd__or2_1
XFILLER_161_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10120_ _10126_/C _10114_/X _10119_/Y vssd1 vssd1 vccd1 vccd1 _12456_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__07835__C _08180_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _12369_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10051_ _10052_/B _10045_/X _10050_/Y vssd1 vssd1 vccd1 vccd1 _12441_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__11162__A1 _11160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11654__A _11680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ _13810_/A _06805_/X vssd1 vssd1 vccd1 vccd1 _14066_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13741_ _13741_/A _06990_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[30] sky130_fd_sc_hd__ebufn_8
XANTENNA__09124__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ _10953_/A vssd1 vssd1 vccd1 vccd1 _12663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13672_ _13672_/A _07167_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
X_10884_ _12646_/Q vssd1 vssd1 vccd1 vccd1 _10908_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12623_ _12625_/CLK _12623_/D vssd1 vssd1 vccd1 vccd1 _12623_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_23_clk _12881_/CLK vssd1 vssd1 vccd1 vccd1 _12867_/CLK sky130_fd_sc_hd__clkbuf_16
X_12554_ _12554_/CLK _12554_/D vssd1 vssd1 vccd1 vccd1 _13682_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11505_ _12807_/Q _11505_/B vssd1 vssd1 vccd1 vccd1 _11506_/A sky130_fd_sc_hd__and2b_1
XFILLER_129_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ _12492_/CLK _12485_/D vssd1 vssd1 vccd1 vccd1 _13615_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11436_ _13912_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11436_/X sky130_fd_sc_hd__or2_1
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11367_ _13914_/A _12771_/Q _11373_/S vssd1 vssd1 vccd1 vccd1 _11368_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _13653_/A _12507_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10319_/B sky130_fd_sc_hd__mux2_1
X_14086_ _14086_/A _08056_/X vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__ebufn_8
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _10652_/X _11284_/X _11297_/X _11293_/X vssd1 vssd1 vccd1 vccd1 _12748_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ _10278_/A vssd1 vssd1 vccd1 vccd1 _10249_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11283__B _11283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13939_ _13939_/A _06448_/X vssd1 vssd1 vccd1 vccd1 _14067_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA_clkbuf_leaf_62_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07460_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07460_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06411_ _06411_/A vssd1 vssd1 vccd1 vccd1 _06411_/X sky130_fd_sc_hd__clkbuf_1
X_07391_ _07396_/A _07391_/B _07401_/C vssd1 vssd1 vccd1 vccd1 _07392_/A sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_14_clk _12217_/CLK vssd1 vssd1 vccd1 vccd1 _12981_/CLK sky130_fd_sc_hd__clkbuf_16
X_09130_ _09152_/B vssd1 vssd1 vccd1 vccd1 _09130_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06342_ _06346_/A _06349_/B _06349_/C vssd1 vssd1 vccd1 vccd1 _06343_/A sky130_fd_sc_hd__or3_1
XANTENNA__06393__A _07861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__B1 _09392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ _11688_/A _11687_/C _12848_/Q _11687_/A _08941_/X _08942_/X vssd1 vssd1 vccd1
+ vccd1 _09061_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06273_ input8/X input11/X input10/X input9/X vssd1 vssd1 vccd1 vccd1 _09097_/C sky130_fd_sc_hd__or4b_2
X_08012_ _08186_/A vssd1 vssd1 vccd1 vccd1 _08067_/A sky130_fd_sc_hd__buf_2
XFILLER_144_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13285__441 vssd1 vssd1 vccd1 vccd1 _13285__441/HI _13990_/A sky130_fd_sc_hd__conb_1
XFILLER_143_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11458__B _11460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _13596_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09963_/X sky130_fd_sc_hd__or2_1
XANTENNA__08113__A _08122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08914_ _12807_/Q _12808_/Q _12809_/Q _11518_/A _08911_/X _08913_/X vssd1 vssd1 vccd1
+ vccd1 _08914_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13954__A _13954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09894_ _13525_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09894_/X sky130_fd_sc_hd__or2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13326__482 vssd1 vssd1 vccd1 vccd1 _13326__482/HI _14079_/A sky130_fd_sc_hd__conb_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_clk_A _12217_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _12649_/Q vssd1 vssd1 vccd1 vccd1 _10907_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08776_ _08770_/X _08775_/X _13780_/A vssd1 vssd1 vccd1 vccd1 _10163_/B sky130_fd_sc_hd__mux2_1
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ _07727_/A _07737_/B _07732_/C vssd1 vssd1 vccd1 vccd1 _07728_/A sky130_fd_sc_hd__or3_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08943__S0 _08941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ _07698_/A vssd1 vssd1 vccd1 vccd1 _07669_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06609_ _06609_/A vssd1 vssd1 vccd1 vccd1 _06609_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09598__B _13553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07589_ _07589_/A vssd1 vssd1 vccd1 vccd1 _07589_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_8_0_clk clkbuf_4_9_0_clk/A vssd1 vssd1 vccd1 vccd1 _12881_/CLK sky130_fd_sc_hd__clkbuf_2
X_09328_ _09328_/A _09328_/B _09328_/C vssd1 vssd1 vccd1 vccd1 _09331_/B sky130_fd_sc_hd__and3_1
XANTENNA__07399__A _07822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09259_ _09316_/A _09316_/B _09317_/C _09317_/D vssd1 vssd1 vccd1 vccd1 _09260_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_127_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _12274_/CLK _12270_/D vssd1 vssd1 vccd1 vccd1 _12270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ _11221_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11222_/A sky130_fd_sc_hd__and2_1
XFILLER_153_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11152_ _11152_/A vssd1 vssd1 vccd1 vccd1 _12710_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09119__A peripheralBus_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10103_ _10101_/B _10053_/B _10101_/D _10101_/A vssd1 vssd1 vccd1 vccd1 _10104_/C
+ sky130_fd_sc_hd__a31o_1
X_11083_ _11083_/A vssd1 vssd1 vccd1 vccd1 _12696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10034_ _12437_/Q vssd1 vssd1 vccd1 vccd1 _10097_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10699__S _10703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08839__A0 _08764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11985_ _11985_/A vssd1 vssd1 vccd1 vccd1 _12920_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09789__A hold2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10936_ _10936_/A _10936_/B _10936_/C vssd1 vssd1 vccd1 vccd1 _10937_/A sky130_fd_sc_hd__and3_1
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13724_ _13724_/A _07030_/X vssd1 vssd1 vccd1 vccd1 _14108_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_17_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13655_ _13655_/A _07212_/X vssd1 vssd1 vccd1 vccd1 _14103_/Z sky130_fd_sc_hd__ebufn_8
X_10867_ _10875_/B _10875_/C vssd1 vssd1 vccd1 vccd1 _10871_/A sky130_fd_sc_hd__and2_1
XANTENNA__10728__A _13786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _12802_/CLK _12606_/D vssd1 vssd1 vccd1 vccd1 _13781_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13586_ _13586_/A _07402_/X vssd1 vssd1 vccd1 vccd1 _14034_/Z sky130_fd_sc_hd__ebufn_8
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _10803_/A vssd1 vssd1 vccd1 vccd1 _10798_/X sky130_fd_sc_hd__buf_2
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12537_ _12554_/CLK _12537_/D vssd1 vssd1 vccd1 vccd1 _12537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13269__425 vssd1 vssd1 vccd1 vccd1 _13269__425/HI _13960_/A sky130_fd_sc_hd__conb_1
XFILLER_145_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ _12492_/CLK _12468_/D vssd1 vssd1 vccd1 vccd1 _12468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11419_ _13905_/A _11423_/B vssd1 vssd1 vccd1 vccd1 _11419_/X sky130_fd_sc_hd__or2_1
X_12399_ _12400_/CLK _12399_/D vssd1 vssd1 vccd1 vccd1 _13527_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10463__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06960_ _06960_/A _06965_/B vssd1 vssd1 vccd1 vccd1 _06961_/A sky130_fd_sc_hd__or2_1
X_14069_ _14069_/A _08009_/X vssd1 vssd1 vccd1 vccd1 _14069_/Z sky130_fd_sc_hd__ebufn_8
Xclkbuf_leaf_3_clk _12917_/CLK vssd1 vssd1 vccd1 vccd1 _12895_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12983__139 vssd1 vssd1 vccd1 vccd1 _12983__139/HI _13380_/A sky130_fd_sc_hd__conb_1
X_06891_ _06891_/A vssd1 vssd1 vccd1 vccd1 _06891_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08630_ _08709_/A vssd1 vssd1 vccd1 vccd1 _08630_/X sky130_fd_sc_hd__buf_2
XFILLER_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08561_ _12433_/Q _12434_/Q _12435_/Q _12436_/Q _08559_/X _08560_/X vssd1 vssd1 vccd1
+ vccd1 _08561_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07512_ _07553_/A vssd1 vssd1 vccd1 vccd1 _07524_/C sky130_fd_sc_hd__clkbuf_1
X_08492_ _13394_/A vssd1 vssd1 vccd1 vccd1 _08492_/X sky130_fd_sc_hd__buf_2
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07443_ _07443_/A vssd1 vssd1 vccd1 vccd1 _07443_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09255__B1 _09248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07374_ _07382_/A _07377_/B _07374_/C vssd1 vssd1 vccd1 vccd1 _07375_/A sky130_fd_sc_hd__or3_1
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08108__A _08110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09113_ _14108_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _09113_/X sky130_fd_sc_hd__or2_1
X_06325_ _06462_/A vssd1 vssd1 vccd1 vccd1 _06336_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__13949__A _13949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09044_ _10940_/A vssd1 vssd1 vccd1 vccd1 _13943_/A sky130_fd_sc_hd__buf_4
XFILLER_148_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09946_ _09946_/A vssd1 vssd1 vccd1 vccd1 _12413_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08778__A _10614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11916__B _13364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062__218 vssd1 vssd1 vccd1 vccd1 _13062__218/HI _13537_/A sky130_fd_sc_hd__conb_1
X_09877_ _13519_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09877_/X sky130_fd_sc_hd__or2_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08828_ _13780_/A vssd1 vssd1 vccd1 vccd1 _08890_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _08752_/X _08754_/X _08756_/X _08757_/X _08850_/A _08749_/X vssd1 vssd1 vccd1
+ vccd1 _08759_/X sky130_fd_sc_hd__mux4_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13103__259 vssd1 vssd1 vccd1 vccd1 _13103__259/HI _13612_/A sky130_fd_sc_hd__conb_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11770_ _11770_/A _11770_/B _11770_/C _11770_/D vssd1 vssd1 vccd1 vccd1 _11787_/A
+ sky130_fd_sc_hd__or4_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09402__A _09454_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10721_/A vssd1 vssd1 vccd1 vccd1 _12608_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10548__A _10548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13440_/A _07778_/X vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10652_ _10652_/A vssd1 vssd1 vccd1 vccd1 _10652_/X sky130_fd_sc_hd__buf_4
X_13371_ _13371_/A _08306_/X vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__ebufn_8
X_10583_ _10583_/A vssd1 vssd1 vccd1 vccd1 _12574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ _12349_/CLK _12322_/D vssd1 vssd1 vccd1 vccd1 _12322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07857__A _07857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11379__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ _12258_/CLK _12253_/D vssd1 vssd1 vccd1 vccd1 _12253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11204_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11205_/A sky130_fd_sc_hd__and2_1
XFILLER_107_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12184_ _14096_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12184_/X sky130_fd_sc_hd__or2_1
XFILLER_134_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11135_ _12708_/Q _13949_/A vssd1 vssd1 vccd1 vccd1 _11138_/B sky130_fd_sc_hd__xor2_1
XANTENNA__13594__A _13594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11066_ _11064_/X _11055_/X _11065_/X _11053_/X vssd1 vssd1 vccd1 vccd1 _12691_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10730__B _10732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ _10077_/A vssd1 vssd1 vccd1 vccd1 _10062_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_49_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12069__C1 _11497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11968_ _14107_/Z _14043_/A _11974_/S vssd1 vssd1 vccd1 vccd1 _11969_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13707_ _13707_/A _07072_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
X_10919_ _10921_/B _10915_/X _10936_/A vssd1 vssd1 vccd1 vccd1 _10919_/Y sky130_fd_sc_hd__o21ai_1
X_11899_ _11927_/A _11899_/B vssd1 vssd1 vccd1 vccd1 _11900_/A sky130_fd_sc_hd__and2_1
XFILLER_149_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09237__B1 _09236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13638_ _13638_/A _07259_/X vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__09788__A1 _09116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13569_ _13569_/A _07446_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_158_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07090_ _07090_/A vssd1 vssd1 vccd1 vccd1 _07101_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11289__A _13872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07486__B _08089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09982__A _09982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09800_ _09800_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__and2_1
XANTENNA__09960__A1 _09186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07992_ _07992_/A vssd1 vssd1 vccd1 vccd1 _07992_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09731_ _12341_/Q _13551_/A vssd1 vssd1 vccd1 vccd1 _09735_/A sky130_fd_sc_hd__xor2_1
X_06943_ _06955_/A vssd1 vssd1 vccd1 vccd1 _06953_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09662_ _13488_/A _12342_/Q _09738_/B vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__mux2_1
X_06874_ _07090_/A vssd1 vssd1 vccd1 vccd1 _06884_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__08110__B _08110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08613_ _08604_/X _08606_/X _08610_/X _08612_/X _08583_/X _08584_/X vssd1 vssd1 vccd1
+ vccd1 _08613_/X sky130_fd_sc_hd__mux4_1
XANTENNA_repeater65_A peripheralBus_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09593_ _12318_/Q _13561_/A vssd1 vssd1 vccd1 vccd1 _09597_/A sky130_fd_sc_hd__xor2_1
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08544_ _08461_/X _08488_/X _08516_/X _08543_/X _08467_/X _09157_/A vssd1 vssd1 vccd1
+ vccd1 _08544_/X sky130_fd_sc_hd__mux4_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06846__A _06900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08475_ _12261_/Q _12262_/Q _12263_/Q _12264_/Q _08396_/X _08397_/X vssd1 vssd1 vccd1
+ vccd1 _08475_/X sky130_fd_sc_hd__mux4_2
XFILLER_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07426_ _07430_/A _07435_/B vssd1 vssd1 vccd1 vccd1 _07427_/A sky130_fd_sc_hd__or2_1
XFILLER_50_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11898__S _11898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__A1 _09182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07357_ _07357_/A vssd1 vssd1 vccd1 vccd1 _07357_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06308_ _06320_/A _06308_/B _06308_/C vssd1 vssd1 vccd1 vccd1 _06309_/A sky130_fd_sc_hd__or3_1
XFILLER_136_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07288_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07300_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_108_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ _08976_/X _08980_/X _08978_/X _09026_/X _09024_/X _09013_/X vssd1 vssd1 vccd1
+ vccd1 _09027_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09929_ _09929_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _09929_/X sky130_fd_sc_hd__or2_1
XANTENNA__08506__A2 _08427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10849__B1 _10781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12940_ _12946_/CLK _12940_/D vssd1 vssd1 vccd1 vccd1 _14066_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _12873_/CLK _12871_/D vssd1 vssd1 vccd1 vccd1 _13999_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11822_/A vssd1 vssd1 vccd1 vccd1 _12879_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09132__A _09269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11753_ _12866_/Q _14011_/A _11760_/S vssd1 vssd1 vccd1 vccd1 _11754_/B sky130_fd_sc_hd__mux2_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10278__A _10278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10720_/A _10704_/B vssd1 vssd1 vccd1 vccd1 _10705_/A sky130_fd_sc_hd__or2_1
X_11684_ _11687_/B _11680_/X _11505_/B vssd1 vssd1 vccd1 vccd1 _11684_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_81_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13190__346 vssd1 vssd1 vccd1 vccd1 _13190__346/HI _13797_/A sky130_fd_sc_hd__conb_1
X_13423_ _13423_/A _08132_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[0] sky130_fd_sc_hd__ebufn_8
X_10635_ _11151_/A _10635_/B _10635_/C vssd1 vssd1 vccd1 vccd1 _10636_/A sky130_fd_sc_hd__and3_1
XFILLER_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07587__A _07615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10566_ _13714_/A _12570_/Q _10635_/B vssd1 vssd1 vccd1 vccd1 _10567_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12305_ _12331_/CLK _12305_/D vssd1 vssd1 vccd1 vccd1 _13436_/A sky130_fd_sc_hd__dfxtp_1
X_13231__387 vssd1 vssd1 vccd1 vccd1 _13231__387/HI _13870_/A sky130_fd_sc_hd__conb_1
XANTENNA__10217__S _10220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater133_A _13625_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10497_ _12536_/Q _13745_/A vssd1 vssd1 vccd1 vccd1 _10499_/C sky130_fd_sc_hd__xor2_1
XFILLER_142_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _12289_/CLK _12236_/D vssd1 vssd1 vccd1 vccd1 _12236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09942__A1 _09160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12167_ _12955_/Q _13361_/A vssd1 vssd1 vccd1 vccd1 _12171_/A sky130_fd_sc_hd__xor2_1
XFILLER_122_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13084__240 vssd1 vssd1 vccd1 vccd1 _13084__240/HI _13579_/A sky130_fd_sc_hd__conb_1
XFILLER_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11118_ _13852_/A _12707_/Q _11118_/S vssd1 vssd1 vccd1 vccd1 _11119_/B sky130_fd_sc_hd__mux2_1
XFILLER_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08211__A _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ _11064_/X _12088_/X _12096_/X _12097_/X vssd1 vssd1 vccd1 vccd1 _12950_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11049_ _13815_/A _11051_/B vssd1 vssd1 vccd1 vccd1 _11049_/X sky130_fd_sc_hd__or2_1
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 peripheralBus_address[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
X_13125__281 vssd1 vssd1 vccd1 vccd1 _13125__281/HI _13666_/A sky130_fd_sc_hd__conb_1
XANTENNA__06369__C _07822_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06590_ _06590_/A vssd1 vssd1 vccd1 vccd1 _06590_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06666__A _06680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09977__A _09977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ _08260_/A vssd1 vssd1 vccd1 vccd1 _08260_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08681__A1 _08568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07211_ _07220_/A _07216_/B _07213_/C vssd1 vssd1 vccd1 vccd1 _07212_/A sky130_fd_sc_hd__or3_1
XFILLER_165_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08191_ _08198_/A _08195_/B _08198_/C vssd1 vssd1 vccd1 vccd1 _08192_/A sky130_fd_sc_hd__or3_1
X_07142_ _07152_/A _07145_/B _07142_/C vssd1 vssd1 vccd1 vccd1 _07143_/A sky130_fd_sc_hd__or3_1
XFILLER_118_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07073_ _07079_/A _07076_/B _07073_/C vssd1 vssd1 vccd1 vccd1 _07074_/A sky130_fd_sc_hd__or3_1
XFILLER_160_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12989__145 vssd1 vssd1 vccd1 vccd1 _12989__145/HI _13386_/A sky130_fd_sc_hd__conb_1
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14123__A _14123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07975_ _08075_/A _08075_/B _07977_/C vssd1 vssd1 vccd1 vccd1 _07976_/A sky130_fd_sc_hd__or3_1
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08121__A _08121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10370__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09714_ _12350_/Q _13560_/A vssd1 vssd1 vccd1 vccd1 _09714_/Y sky130_fd_sc_hd__xnor2_1
X_06926_ _06974_/A vssd1 vssd1 vccd1 vccd1 _06936_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09645_ _13466_/A _09640_/X _09644_/X _09634_/X vssd1 vssd1 vccd1 vccd1 _12336_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08595__S1 _08557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06857_ _06863_/A _06857_/B _06857_/C vssd1 vssd1 vccd1 vccd1 _06858_/A sky130_fd_sc_hd__or3_1
XFILLER_55_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09576_ _09579_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__and2_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _06788_/A _06793_/B _06793_/C vssd1 vssd1 vccd1 vccd1 _06789_/A sky130_fd_sc_hd__or3_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08390_/X _08469_/X _08496_/X _08526_/X _08448_/X _08517_/X vssd1 vssd1 vccd1
+ vccd1 _08527_/X sky130_fd_sc_hd__mux4_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08458_ _09330_/A _12256_/Q _09328_/A _09336_/A _08445_/X _08446_/X vssd1 vssd1 vccd1
+ vccd1 _08458_/X sky130_fd_sc_hd__mux4_2
XFILLER_143_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09102__D _12062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07409_ _07409_/A vssd1 vssd1 vccd1 vccd1 _07409_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08389_ _12252_/Q _12253_/Q _12254_/Q _12255_/Q _08379_/X _08380_/X vssd1 vssd1 vccd1
+ vccd1 _08389_/X sky130_fd_sc_hd__mux4_2
X_10420_ _10288_/X _10409_/X _10419_/X _10412_/X vssd1 vssd1 vccd1 vccd1 _12531_/D
+ sky130_fd_sc_hd__o211a_1
X_10351_ _12510_/Q _13752_/A vssd1 vssd1 vccd1 vccd1 _10351_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_164_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10282_ _13626_/A _10291_/B vssd1 vssd1 vccd1 vccd1 _10282_/X sky130_fd_sc_hd__or2_1
X_13068__224 vssd1 vssd1 vccd1 vccd1 _13068__224/HI _13543_/A sky130_fd_sc_hd__conb_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12021_ _12030_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12022_/A sky130_fd_sc_hd__and2_1
XFILLER_105_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07854__B _07854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__A _09919_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13109__265 vssd1 vssd1 vccd1 vccd1 _13109__265/HI _13634_/A sky130_fd_sc_hd__conb_1
XANTENNA__13872__A _13872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13972_ _13972_/A _06360_/X vssd1 vssd1 vccd1 vccd1 _14068_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07870__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ _12923_/CLK _12923_/D vssd1 vssd1 vccd1 vccd1 _12923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _12935_/CLK _12854_/D vssd1 vssd1 vccd1 vccd1 _12854_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _09625_/A _14003_/A _11805_/S vssd1 vssd1 vccd1 vccd1 _11806_/B sky130_fd_sc_hd__mux2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _12786_/CLK _12785_/D vssd1 vssd1 vccd1 vccd1 _13911_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _12861_/Q _14006_/A _11743_/S vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__mux2_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11667_ _11676_/B _11667_/B vssd1 vssd1 vccd1 vccd1 _11668_/C sky130_fd_sc_hd__nand2_1
XFILLER_128_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13406_ _13406_/A _07978_/X vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_127_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10618_ _12577_/Q _13753_/A vssd1 vssd1 vccd1 vccd1 _10622_/A sky130_fd_sc_hd__xor2_1
XFILLER_128_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11598_ _11598_/A vssd1 vssd1 vccd1 vccd1 _12828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10549_ _13693_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10549_/X sky130_fd_sc_hd__or2_1
XFILLER_128_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12219_ _12295_/CLK _12219_/D vssd1 vssd1 vccd1 vccd1 _13396_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10930__C1 _10749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__A0 _13493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ _07760_/A vssd1 vssd1 vccd1 vccd1 _07760_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06711_ _06711_/A vssd1 vssd1 vccd1 vccd1 _06711_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11486__A0 _14103_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08577__S1 _08576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07691_ _07699_/A _07696_/B _07691_/C vssd1 vssd1 vccd1 vccd1 _07692_/A sky130_fd_sc_hd__or3_1
X_09430_ _09430_/A vssd1 vssd1 vccd1 vccd1 _12282_/D sky130_fd_sc_hd__clkbuf_1
X_06642_ _06729_/A _07323_/B _06651_/C vssd1 vssd1 vccd1 vccd1 _06643_/A sky130_fd_sc_hd__or3_1
XFILLER_25_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09361_ _09362_/B _09362_/C _09355_/B _09362_/A vssd1 vssd1 vccd1 vccd1 _09365_/B
+ sky130_fd_sc_hd__a31o_1
X_06573_ _06573_/A vssd1 vssd1 vccd1 vccd1 _06573_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08312_ _08312_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08313_/A sky130_fd_sc_hd__or2_1
X_09292_ _09330_/C _09330_/D _09292_/C vssd1 vssd1 vccd1 vccd1 _09300_/C sky130_fd_sc_hd__and3_1
XFILLER_60_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09500__A _09513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _08243_/A vssd1 vssd1 vccd1 vccd1 _08243_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08174_ _08174_/A _08174_/B _08184_/C vssd1 vssd1 vccd1 vccd1 _08175_/A sky130_fd_sc_hd__or3_1
XANTENNA__10365__B _13745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__A _08122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ _07125_/A vssd1 vssd1 vccd1 vccd1 _07125_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07056_ _07056_/A vssd1 vssd1 vccd1 vccd1 _07056_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09873__C _10637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09906__A1 _09182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10381__A _10423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07958_ _07983_/A _07971_/B _07962_/C vssd1 vssd1 vccd1 vccd1 _07959_/A sky130_fd_sc_hd__or3_1
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08786__A _13777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08568__S1 _08560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__B _11924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06909_ _08168_/A _06916_/B vssd1 vssd1 vccd1 vccd1 _06910_/A sky130_fd_sc_hd__or2_1
X_07889_ _07889_/A vssd1 vssd1 vccd1 vccd1 _07889_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09628_ _09655_/B vssd1 vssd1 vccd1 vccd1 _09638_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_28_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09559_ _09563_/A _09559_/B vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__and2_1
XFILLER_62_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12570_ _12599_/CLK _12570_/D vssd1 vssd1 vccd1 vccd1 _12570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11521_ _11582_/C vssd1 vssd1 vccd1 vccd1 _11521_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11452_ _13918_/A _11452_/B vssd1 vssd1 vccd1 vccd1 _11452_/X sky130_fd_sc_hd__or2_1
X_10403_ _09767_/X _10395_/X _10402_/X _10398_/X vssd1 vssd1 vccd1 vccd1 _12525_/D
+ sky130_fd_sc_hd__o211a_1
X_11383_ _11383_/A vssd1 vssd1 vccd1 vccd1 _12775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07865__A _07892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _10988_/A vssd1 vssd1 vccd1 vccd1 _10479_/A sky130_fd_sc_hd__buf_2
XFILLER_125_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _10293_/B vssd1 vssd1 vccd1 vccd1 _10276_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12004_ _12013_/A _12004_/B vssd1 vssd1 vccd1 vccd1 _12005_/A sky130_fd_sc_hd__and2_1
XFILLER_120_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10196_ _10196_/A vssd1 vssd1 vccd1 vccd1 _12475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13343__499 vssd1 vssd1 vccd1 vccd1 _13343__499/HI _14112_/A sky130_fd_sc_hd__conb_1
XFILLER_93_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11468__A0 _14097_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13955_ _13955_/A _06409_/X vssd1 vssd1 vccd1 vccd1 _13987_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12906_ _12908_/CLK _12906_/D vssd1 vssd1 vccd1 vccd1 _14033_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _13886_/A _06596_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
X_13196__352 vssd1 vssd1 vccd1 vccd1 _13196__352/HI _13803_/A sky130_fd_sc_hd__conb_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12842_/CLK _12837_/D vssd1 vssd1 vccd1 vccd1 _12837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12768_ _12768_/CLK _12768_/D vssd1 vssd1 vccd1 vccd1 _12768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13237__393 vssd1 vssd1 vccd1 vccd1 _13237__393/HI _13892_/A sky130_fd_sc_hd__conb_1
X_11719_ _12856_/Q _14001_/A _11726_/S vssd1 vssd1 vccd1 vccd1 _11720_/B sky130_fd_sc_hd__mux2_1
XFILLER_159_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12699_ _12699_/CLK _12699_/D vssd1 vssd1 vccd1 vccd1 _12699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput10 peripheralBus_address[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
Xinput21 peripheralBus_address[6] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__13777__A _13777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08930_ _11639_/C _12824_/Q _12825_/Q _12826_/Q _08928_/X _08929_/X vssd1 vssd1 vccd1
+ vccd1 _08930_/X sky130_fd_sc_hd__mux4_2
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08861_ _10907_/C _12651_/Q _10907_/A _12653_/Q _08807_/X _08808_/X vssd1 vssd1 vccd1
+ vccd1 _08861_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07812_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07868_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08792_ _12643_/Q vssd1 vssd1 vccd1 vccd1 _10874_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07743_ _07743_/A vssd1 vssd1 vccd1 vccd1 _07743_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07674_ _07923_/A vssd1 vssd1 vccd1 vccd1 _07729_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _09413_/A vssd1 vssd1 vccd1 vccd1 _12277_/D sky130_fd_sc_hd__clkbuf_1
X_06625_ _06625_/A _06630_/B _06630_/C vssd1 vssd1 vccd1 vccd1 _06626_/A sky130_fd_sc_hd__or3_1
XFILLER_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08970__S1 _08968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09344_ _09352_/C _09344_/B vssd1 vssd1 vccd1 vccd1 _09344_/Y sky130_fd_sc_hd__nand2_1
X_06556_ _06556_/A _06561_/B _06561_/C vssd1 vssd1 vccd1 vccd1 _06557_/A sky130_fd_sc_hd__or3_1
X_09275_ _09284_/D _09276_/C _09274_/Y vssd1 vssd1 vccd1 vccd1 _12246_/D sky130_fd_sc_hd__a21oi_1
X_06487_ _06487_/A vssd1 vssd1 vccd1 vccd1 _06487_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08226_ _08226_/A vssd1 vssd1 vccd1 vccd1 _08226_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _08157_/A vssd1 vssd1 vccd1 vccd1 _08157_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07108_ _07108_/A _07118_/B _07115_/C vssd1 vssd1 vccd1 vccd1 _07109_/A sky130_fd_sc_hd__or3_1
XFILLER_161_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11919__B _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ _08088_/A vssd1 vssd1 vccd1 vccd1 _08088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07039_ _07043_/A _07043_/B vssd1 vssd1 vccd1 vccd1 _07040_/A sky130_fd_sc_hd__or2_1
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13030__186 vssd1 vssd1 vccd1 vccd1 _13030__186/HI _13473_/A sky130_fd_sc_hd__conb_1
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10050_ _10052_/B _10045_/X _10123_/A vssd1 vssd1 vccd1 vccd1 _10050_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11698__B1 _11576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13740_ _13740_/A _06992_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[29] sky130_fd_sc_hd__ebufn_8
XFILLER_113_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10952_ _10952_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _10953_/A sky130_fd_sc_hd__and2_1
XFILLER_56_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13671_ _13671_/A _07170_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
X_10883_ _10922_/B _10883_/B vssd1 vssd1 vccd1 vccd1 _12645_/D sky130_fd_sc_hd__nor2_1
XFILLER_44_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12622_ _12625_/CLK _12622_/D vssd1 vssd1 vccd1 vccd1 _12622_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09140__A _09140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12553_ _12554_/CLK _12553_/D vssd1 vssd1 vccd1 vccd1 _13681_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11504_ _11520_/A vssd1 vssd1 vccd1 vccd1 _11505_/B sky130_fd_sc_hd__buf_4
X_12484_ _12656_/CLK _12484_/D vssd1 vssd1 vccd1 vccd1 _13762_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11435_ _10665_/X _11425_/X _11434_/X _11430_/X vssd1 vssd1 vccd1 vccd1 _12785_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11366_ _11366_/A vssd1 vssd1 vccd1 vccd1 _12770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10317_ _10317_/A vssd1 vssd1 vccd1 vccd1 _10332_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _14085_/A _08053_/X vssd1 vssd1 vccd1 vccd1 _14117_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_113_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11297_ _13875_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11297_/X sky130_fd_sc_hd__or2_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _11028_/B _12060_/A _10693_/C vssd1 vssd1 vccd1 vccd1 _10278_/A sky130_fd_sc_hd__or3_4
XFILLER_79_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10179_ _10179_/A vssd1 vssd1 vccd1 vccd1 _12470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12102__A1 _10552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11283__C _11410_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13938_ _13938_/A _06450_/X vssd1 vssd1 vccd1 vccd1 _14066_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_34_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06377__C _06377_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__A1 _10662_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ _13869_/A _06645_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[30] sky130_fd_sc_hd__ebufn_8
X_06410_ _06416_/A _06412_/B vssd1 vssd1 vccd1 vccd1 _06411_/A sky130_fd_sc_hd__or2_1
X_07390_ _07403_/A vssd1 vssd1 vccd1 vccd1 _07401_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10416__A1 _10414_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06341_ _06341_/A vssd1 vssd1 vccd1 vccd1 _06341_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ _12849_/Q vssd1 vssd1 vccd1 vccd1 _11687_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06272_ input14/X input13/X input16/X input15/X vssd1 vssd1 vccd1 vccd1 _09097_/B
+ sky130_fd_sc_hd__or4_4
X_08011_ _08011_/A vssd1 vssd1 vccd1 vccd1 _08011_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09962_ _09092_/X _09934_/S _09961_/X _09959_/X vssd1 vssd1 vccd1 vccd1 _12419_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_repeater95_A peripheralBus_data[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08913_ _09068_/A vssd1 vssd1 vccd1 vccd1 _08913_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_134_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09893_ _09160_/X _09888_/X _09890_/X _09892_/X vssd1 vssd1 vccd1 vccd1 _12396_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08844_ _08782_/X _08787_/X _08783_/X _08790_/X _08837_/X _08838_/X vssd1 vssd1 vccd1
+ vccd1 _08844_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08640__S0 _08575_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08775_ _08771_/X _08772_/X _08773_/X _08774_/X _08850_/A _08769_/X vssd1 vssd1 vccd1
+ vccd1 _08775_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07726_ _07892_/A vssd1 vssd1 vccd1 vccd1 _07737_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07657_ _07657_/A vssd1 vssd1 vccd1 vccd1 _07657_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08943__S1 _08942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__A _11490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06608_ _06610_/A _06616_/B _06616_/C vssd1 vssd1 vccd1 vccd1 _06609_/A sky130_fd_sc_hd__or3_1
X_07588_ _07588_/A _07598_/B _07593_/C vssd1 vssd1 vccd1 vccd1 _07589_/A sky130_fd_sc_hd__or3_1
XFILLER_159_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10407__A1 _09773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09327_ _09327_/A vssd1 vssd1 vccd1 vccd1 _12257_/D sky130_fd_sc_hd__clkbuf_1
X_06539_ _06539_/A vssd1 vssd1 vccd1 vccd1 _06539_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09258_ _09315_/A _09315_/B _09317_/A _09258_/D vssd1 vssd1 vccd1 vccd1 _09260_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_138_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08209_ _08209_/A vssd1 vssd1 vccd1 vccd1 _08209_/X sky130_fd_sc_hd__clkbuf_1
X_09189_ _13403_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _09189_/X sky130_fd_sc_hd__or2_1
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11220_ _13876_/A _12732_/Q _11231_/S vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__mux2_1
XFILLER_153_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11151_ _11151_/A _11151_/B _11151_/C vssd1 vssd1 vccd1 vccd1 _11152_/A sky130_fd_sc_hd__and3_1
XFILLER_150_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10102_ _10112_/B vssd1 vssd1 vccd1 vccd1 _10133_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11082_ _11095_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11083_/A sky130_fd_sc_hd__and2_1
XANTENNA__08536__A0 _08423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10033_ _10033_/A _10089_/A vssd1 vssd1 vccd1 vccd1 _12436_/D sky130_fd_sc_hd__nor2_1
XFILLER_76_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11384__B _11384_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A peripheralBus_address[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11984_ _11996_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _11985_/A sky130_fd_sc_hd__and2_1
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11843__A0 peripheralBus_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13723_ _13723_/A _07032_/X vssd1 vssd1 vccd1 vccd1 _14075_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__09789__B _09789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10935_ _12660_/Q _10935_/B vssd1 vssd1 vccd1 vccd1 _10936_/C sky130_fd_sc_hd__nand2_1
XFILLER_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13654_ _13654_/A _07214_/X vssd1 vssd1 vccd1 vccd1 _13974_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10866_ _10866_/A _10866_/B _10866_/C _10866_/D vssd1 vssd1 vccd1 vccd1 _10881_/B
+ sky130_fd_sc_hd__and4_1
X_12605_ _12802_/CLK _12605_/D vssd1 vssd1 vccd1 vccd1 _13780_/A sky130_fd_sc_hd__dfxtp_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13585_/A _07405_/X vssd1 vssd1 vccd1 vccd1 _14033_/Z sky130_fd_sc_hd__ebufn_8
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10797_ _10797_/A vssd1 vssd1 vccd1 vccd1 _12626_/D sky130_fd_sc_hd__clkbuf_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11071__A1 _10552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12536_ _12554_/CLK _12536_/D vssd1 vssd1 vccd1 vccd1 _12536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12467_ _12467_/CLK _12467_/D vssd1 vssd1 vccd1 vccd1 _12467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11418_ _11160_/X _11411_/X _11416_/X _11417_/X vssd1 vssd1 vccd1 vccd1 _12778_/D
+ sky130_fd_sc_hd__o211a_1
X_12398_ _12418_/CLK _12398_/D vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08214__A _08240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11349_ _11349_/A vssd1 vssd1 vccd1 vccd1 _12765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14068_ _14068_/A _08006_/X vssd1 vssd1 vccd1 vccd1 _14068_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06890_ _06890_/A _06898_/B _06898_/C vssd1 vssd1 vccd1 vccd1 _06891_/A sky130_fd_sc_hd__or3_1
XFILLER_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08560_ _13585_/A vssd1 vssd1 vccd1 vccd1 _08560_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07511_ _07511_/A vssd1 vssd1 vccd1 vccd1 _07511_/X sky130_fd_sc_hd__clkbuf_1
X_08491_ _11705_/D vssd1 vssd1 vccd1 vccd1 _13366_/A sky130_fd_sc_hd__buf_4
XFILLER_81_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07442_ _07442_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07443_/A sky130_fd_sc_hd__or2_1
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07373_ _07373_/A vssd1 vssd1 vccd1 vccd1 _07373_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09112_ _11064_/A vssd1 vssd1 vccd1 vccd1 _09112_/X sky130_fd_sc_hd__clkbuf_4
X_06324_ _06324_/A vssd1 vssd1 vccd1 vccd1 _06324_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09043_ _09040_/X _09042_/X _09043_/S vssd1 vssd1 vccd1 vccd1 _10940_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07947__B _07947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08861__S0 _08807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ _10700_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _09946_/A sky130_fd_sc_hd__or2_1
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09876_ _09915_/B vssd1 vssd1 vccd1 vccd1 _09886_/B sky130_fd_sc_hd__clkbuf_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10820__C _10820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08827_ _08815_/X _08818_/X _08822_/X _08825_/X _08826_/X _08812_/X vssd1 vssd1 vccd1
+ vccd1 _08827_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08758_ _13778_/A vssd1 vssd1 vccd1 vccd1 _08850_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13142__298 vssd1 vssd1 vccd1 vccd1 _13142__298/HI _13699_/A sky130_fd_sc_hd__conb_1
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _07709_/A vssd1 vssd1 vccd1 vccd1 _07709_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _08610_/X _08612_/X _08614_/X _08615_/X _08678_/X _08647_/X vssd1 vssd1 vccd1
+ vccd1 _08689_/X sky130_fd_sc_hd__mux4_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _10720_/A _10720_/B vssd1 vssd1 vccd1 vccd1 _10721_/A sky130_fd_sc_hd__or2_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10651_ _10648_/X _10638_/X _10649_/X _10650_/X vssd1 vssd1 vccd1 vccd1 _12587_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _13370_/A _08304_/X vssd1 vssd1 vccd1 vccd1 _14106_/Z sky130_fd_sc_hd__ebufn_8
X_10582_ _10585_/A _10582_/B vssd1 vssd1 vccd1 vccd1 _10583_/A sky130_fd_sc_hd__and2_1
XFILLER_70_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12321_ _12334_/CLK _12321_/D vssd1 vssd1 vccd1 vccd1 _12321_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07857__B _07962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13036__192 vssd1 vssd1 vccd1 vccd1 _13036__192/HI _13479_/A sky130_fd_sc_hd__conb_1
XFILLER_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12252_ _12258_/CLK _12252_/D vssd1 vssd1 vccd1 vccd1 _12252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11203_ _13871_/A _12727_/Q _11281_/B vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__mux2_1
X_12183_ _12208_/B vssd1 vssd1 vccd1 vccd1 _12193_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_150_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_61_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ _12704_/Q _13945_/A vssd1 vssd1 vccd1 vccd1 _11138_/A sky130_fd_sc_hd__xor2_1
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11065_ _13820_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11065_/X sky130_fd_sc_hd__or2_1
XFILLER_122_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08604__S0 _08602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06489__A _08276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10016_ _10021_/B _10021_/C _10016_/C vssd1 vssd1 vccd1 vccd1 _10024_/C sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_76_clk_A _12555_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11967_ _11967_/A vssd1 vssd1 vccd1 vccd1 _12915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10739__A _10820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13706_ _13706_/A _07074_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
X_10918_ _10918_/A vssd1 vssd1 vccd1 vccd1 _12654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11898_ _12902_/Q _14046_/A _11898_/S vssd1 vssd1 vccd1 vccd1 _11899_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13637_ _13637_/A _07261_/X vssd1 vssd1 vccd1 vccd1 _13765_/Z sky130_fd_sc_hd__ebufn_8
X_10849_ _10875_/B _10847_/A _10781_/X vssd1 vssd1 vccd1 vccd1 _10850_/B sky130_fd_sc_hd__o21ai_1
XFILLER_158_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11044__A1 _10394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A _12217_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13568_ _13568_/A _07448_/X vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_145_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12519_ _12522_/CLK _12519_/D vssd1 vssd1 vccd1 vccd1 _13648_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13499_ _13499_/A _07625_/X vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clk_A _12759_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13785__A _13785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07991_ _07997_/A _08184_/B _07993_/C vssd1 vssd1 vccd1 vccd1 _07992_/A sky130_fd_sc_hd__or3_1
XFILLER_141_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_clk clkbuf_4_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_09730_ _09730_/A _09730_/B _09730_/C _09730_/D vssd1 vssd1 vccd1 vccd1 _09736_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06942_ _06942_/A vssd1 vssd1 vccd1 vccd1 _06942_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09661_ _09661_/A vssd1 vssd1 vccd1 vccd1 _12341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06873_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07090_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__08110__C _08110_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ _10029_/B _10029_/A _12437_/Q _12438_/Q _08553_/X _08554_/X vssd1 vssd1 vccd1
+ vccd1 _08612_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09592_ _09587_/X _09588_/Y _09589_/Y _09590_/X _09591_/Y vssd1 vssd1 vccd1 vccd1
+ _09592_/X sky130_fd_sc_hd__o221a_1
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08543_ _09382_/A _09388_/B _12273_/Q _12274_/Q _09140_/A _09146_/A vssd1 vssd1 vccd1
+ vccd1 _08543_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08474_ _08398_/X _08401_/X _08400_/X _08406_/X _08517_/A _08467_/X vssd1 vssd1 vccd1
+ vccd1 _08474_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10368__B _13751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07425_ _08131_/C vssd1 vssd1 vccd1 vccd1 _07435_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11035__A1 _10645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07356_ _07356_/A _07364_/B _07361_/C vssd1 vssd1 vccd1 vccd1 _07357_/A sky130_fd_sc_hd__or3_1
XFILLER_164_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06307_ _06361_/A vssd1 vssd1 vccd1 vccd1 _06320_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07287_ _07287_/A vssd1 vssd1 vccd1 vccd1 _07287_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09026_ _11661_/B _12842_/Q _12843_/Q _12844_/Q _08967_/X _08968_/X vssd1 vssd1 vccd1
+ vccd1 _09026_/X sky130_fd_sc_hd__mux4_2
XFILLER_136_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11199__B _11199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09928_ _09124_/X _09921_/X _09927_/X _09916_/X vssd1 vssd1 vccd1 vccd1 _12407_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09859_ _12376_/Q _13553_/A vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__xor2_1
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12870_ _12903_/CLK _12870_/D vssd1 vssd1 vccd1 vccd1 _13378_/A sky130_fd_sc_hd__dfxtp_4
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11834_/A _11821_/B vssd1 vssd1 vccd1 vccd1 _11822_/A sky130_fd_sc_hd__and2_1
XFILLER_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11752_/A vssd1 vssd1 vccd1 vccd1 _12865_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _14098_/Z _08850_/X _10703_/S vssd1 vssd1 vccd1 vccd1 _10704_/B sky130_fd_sc_hd__mux2_1
XFILLER_81_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11683_/A vssd1 vssd1 vccd1 vccd1 _12847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07868__A _07868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13422_ _13422_/A _07838_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
X_10634_ _10611_/Y _10617_/X _10633_/Y _13759_/A vssd1 vssd1 vccd1 vccd1 _10635_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_139_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10565_ _10565_/A vssd1 vssd1 vccd1 vccd1 _12569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12304_ _12331_/CLK _12304_/D vssd1 vssd1 vccd1 vccd1 _13435_/A sky130_fd_sc_hd__dfxtp_1
X_10496_ _12546_/Q _13755_/A vssd1 vssd1 vccd1 vccd1 _10499_/B sky130_fd_sc_hd__xor2_1
XFILLER_6_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12235_ _12289_/CLK _12235_/D vssd1 vssd1 vccd1 vccd1 _12235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08825__S0 _08807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _12166_/A _12166_/B _12166_/C _12166_/D vssd1 vssd1 vccd1 vccd1 _12177_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold2_A hold2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ _11117_/A vssd1 vssd1 vccd1 vccd1 _12706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12097_ _12200_/A vssd1 vssd1 vccd1 vccd1 _12097_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output55_A _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11048_ _10662_/X _11041_/X _11047_/X _11039_/X vssd1 vssd1 vccd1 vccd1 _12685_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 peripheralBus_address[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09002__S0 _08967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07210_ _07210_/A vssd1 vssd1 vccd1 vccd1 _07210_/X sky130_fd_sc_hd__clkbuf_1
X_08190_ _08190_/A vssd1 vssd1 vccd1 vccd1 _08190_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06682__A _06686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07141_ _07141_/A vssd1 vssd1 vccd1 vccd1 _07141_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07072_ _07072_/A vssd1 vssd1 vccd1 vccd1 _07072_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07974_ _07974_/A vssd1 vssd1 vccd1 vccd1 _07974_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09713_ _09713_/A vssd1 vssd1 vccd1 vccd1 _12356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06925_ _07480_/A vssd1 vssd1 vccd1 vccd1 _06974_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09644_ _11189_/A _09653_/B vssd1 vssd1 vccd1 vccd1 _09644_/X sky130_fd_sc_hd__or2_1
X_06856_ _06856_/A vssd1 vssd1 vccd1 vccd1 _06856_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09575_ _13468_/A _12321_/Q _09575_/S vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__mux2_1
X_06787_ _06787_/A vssd1 vssd1 vccd1 vccd1 _06787_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10379__A _10409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _09377_/C _12269_/Q _09377_/A _09382_/A _09140_/A _09146_/A vssd1 vssd1 vccd1
+ vccd1 _08526_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08457_ _12258_/Q vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07408_ _07822_/A _07840_/B _07496_/C vssd1 vssd1 vccd1 vccd1 _07409_/A sky130_fd_sc_hd__or3_1
X_08388_ _12248_/Q _12249_/Q _09321_/B _12251_/Q _08376_/X _08377_/X vssd1 vssd1 vccd1
+ vccd1 _08388_/X sky130_fd_sc_hd__mux4_2
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07339_ _07393_/A vssd1 vssd1 vccd1 vccd1 _07351_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_164_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10350_ _10350_/A vssd1 vssd1 vccd1 vccd1 _12516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09009_ _08999_/X _09002_/X _09004_/X _09008_/X _08994_/X _08953_/X vssd1 vssd1 vccd1
+ vccd1 _09009_/X sky130_fd_sc_hd__mux4_1
X_10281_ _09182_/X _10278_/X _10280_/X _10270_/X vssd1 vssd1 vccd1 vccd1 _12495_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12020_ _12931_/Q _14074_/A _12029_/S vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07854__C _08180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13971_ _13971_/A _06363_/X vssd1 vssd1 vccd1 vccd1 _14099_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_19_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11495__A1 _13978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ _12923_/CLK _12922_/D vssd1 vssd1 vccd1 vccd1 _12922_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06767__A _07603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__B _13949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09143__A _14065_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ _12853_/CLK _12853_/D vssd1 vssd1 vccd1 vccd1 _12853_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11804_ _11804_/A vssd1 vssd1 vccd1 vccd1 _12874_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12786_/CLK _12784_/D vssd1 vssd1 vccd1 vccd1 _13910_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11735_/A vssd1 vssd1 vccd1 vccd1 _12860_/D sky130_fd_sc_hd__clkbuf_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _11676_/B _11667_/B vssd1 vssd1 vccd1 vccd1 _11668_/B sky130_fd_sc_hd__or2_1
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13405_ _13405_/A _07976_/X vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__ebufn_8
X_10617_ _10612_/Y _10613_/X _10614_/X _10615_/Y _10616_/Y vssd1 vssd1 vccd1 vccd1
+ _10617_/X sky130_fd_sc_hd__o221a_1
XFILLER_128_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11597_ _11595_/X _11604_/B _11597_/C vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__and3b_1
XANTENNA__10758__B1 _10757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08206__B _08208_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13348__504 vssd1 vssd1 vccd1 vccd1 _13348__504/HI _14117_/A sky130_fd_sc_hd__conb_1
XFILLER_128_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10548_ _10548_/A vssd1 vssd1 vccd1 vccd1 _10548_/X sky130_fd_sc_hd__buf_6
XFILLER_127_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10479_ _10479_/A vssd1 vssd1 vccd1 vccd1 _10567_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12218_ _12903_/CLK _12218_/D vssd1 vssd1 vccd1 vccd1 _13395_/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__11567__B _11604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12149_ _12149_/A _12149_/B vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__and2_1
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06710_ _06714_/A _06719_/B _06719_/C vssd1 vssd1 vccd1 vccd1 _06711_/A sky130_fd_sc_hd__or3_1
X_07690_ _07690_/A vssd1 vssd1 vccd1 vccd1 _07690_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06641_ _08184_/B vssd1 vssd1 vccd1 vccd1 _06651_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09360_ _09360_/A vssd1 vssd1 vccd1 vccd1 _12265_/D sky130_fd_sc_hd__clkbuf_1
X_06572_ _06584_/A _06574_/B _06574_/C vssd1 vssd1 vccd1 vccd1 _06573_/A sky130_fd_sc_hd__or3_1
X_08311_ _08335_/A vssd1 vssd1 vccd1 vccd1 _08321_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ _09330_/D _09292_/C _09290_/Y vssd1 vssd1 vccd1 vccd1 _12250_/D sky130_fd_sc_hd__a21oi_1
X_08242_ _08251_/A _08248_/B _08251_/C vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__or3_1
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08173_ _08173_/A vssd1 vssd1 vccd1 vccd1 _08173_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07124_ _07135_/A _07131_/B _07128_/C vssd1 vssd1 vccd1 vccd1 _07125_/A sky130_fd_sc_hd__or3_1
XFILLER_106_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07055_ _07055_/A _07055_/B vssd1 vssd1 vccd1 vccd1 _07056_/A sky130_fd_sc_hd__or2_1
XFILLER_106_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10662__A _10662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09367__B1 _09206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09228__A _13391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08132__A _08132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07957_ _07957_/A vssd1 vssd1 vccd1 vccd1 _07957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06908_ _06908_/A vssd1 vssd1 vccd1 vccd1 _06908_/X sky130_fd_sc_hd__clkbuf_1
X_07888_ _07894_/A _07890_/B _07890_/C vssd1 vssd1 vccd1 vccd1 _07889_/A sky130_fd_sc_hd__or3_1
XFILLER_56_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09627_ _09640_/A vssd1 vssd1 vccd1 vccd1 _09627_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06839_ _06850_/A _06843_/B _06843_/C vssd1 vssd1 vccd1 vccd1 _06840_/A sky130_fd_sc_hd__or3_1
XFILLER_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09558_ _13463_/A _12316_/Q _09558_/S vssd1 vssd1 vccd1 vccd1 _09559_/B sky130_fd_sc_hd__mux2_1
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08509_ _08506_/X _08508_/X _08528_/S vssd1 vssd1 vccd1 vccd1 _11707_/C sky130_fd_sc_hd__mux2_1
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09489_ _13424_/A _09483_/X _09488_/X _09192_/X vssd1 vssd1 vccd1 vccd1 _12293_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ _11520_/A vssd1 vssd1 vccd1 vccd1 _11582_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11451_ _10548_/A _11438_/X _11450_/X _11444_/X vssd1 vssd1 vccd1 vccd1 _12791_/D
+ sky130_fd_sc_hd__o211a_1
X_10402_ _13654_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10402_/X sky130_fd_sc_hd__or2_1
XFILLER_164_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11382_ _11723_/A _11382_/B vssd1 vssd1 vccd1 vccd1 _11383_/A sky130_fd_sc_hd__and2_1
XANTENNA__11668__A _11703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10333_ _10333_/A vssd1 vssd1 vccd1 vccd1 _12511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11387__B _11388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09138__A _14096_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ _10278_/A vssd1 vssd1 vccd1 vccd1 _10264_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12003_ _12926_/Q _14069_/A _12012_/S vssd1 vssd1 vccd1 vccd1 _12004_/B sky130_fd_sc_hd__mux2_1
X_10195_ _10208_/A _10195_/B vssd1 vssd1 vccd1 vccd1 _10196_/A sky130_fd_sc_hd__and2_1
XANTENNA__10912__B1 _10757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13954_ _13954_/A _06411_/X vssd1 vssd1 vccd1 vccd1 _14082_/Z sky130_fd_sc_hd__ebufn_8
X_12905_ _12961_/CLK _12905_/D vssd1 vssd1 vccd1 vccd1 _14032_/A sky130_fd_sc_hd__dfxtp_2
X_13885_ _13885_/A _06598_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[14] sky130_fd_sc_hd__ebufn_8
XFILLER_47_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12836_ _12842_/CLK _12836_/D vssd1 vssd1 vccd1 vccd1 _12836_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ _12768_/CLK _12767_/D vssd1 vssd1 vccd1 vccd1 _12767_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10747__A _13775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11718_ _11718_/A vssd1 vssd1 vccd1 vccd1 _12855_/D sky130_fd_sc_hd__clkbuf_1
X_12698_ _12704_/CLK _12698_/D vssd1 vssd1 vccd1 vccd1 _12698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11649_ _11649_/A _11649_/B _11649_/C _11649_/D vssd1 vssd1 vccd1 vccd1 _11688_/B
+ sky130_fd_sc_hd__and4_1
Xinput11 peripheralBus_address[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
Xinput22 peripheralBus_address[7] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07494__C _07496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ _08744_/X _08747_/X _08752_/X _08754_/X _08748_/X _08859_/X vssd1 vssd1 vccd1
+ vccd1 _08860_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07811_ _07923_/A vssd1 vssd1 vccd1 vccd1 _07910_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08791_ _10876_/D _12637_/Q _12638_/Q _12639_/Q _08742_/X _08743_/X vssd1 vssd1 vccd1
+ vccd1 _08791_/X sky130_fd_sc_hd__mux4_2
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07742_ _07742_/A _07753_/B _07748_/C vssd1 vssd1 vccd1 vccd1 _07743_/A sky130_fd_sc_hd__or3_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07673_ _07673_/A vssd1 vssd1 vccd1 vccd1 _07673_/X sky130_fd_sc_hd__clkbuf_1
X_09412_ _09422_/A _09412_/B vssd1 vssd1 vccd1 vccd1 _09413_/A sky130_fd_sc_hd__and2_1
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06624_ _06624_/A vssd1 vssd1 vccd1 vccd1 _06624_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09511__A _09638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _13391_/A _09346_/C _09343_/C _09343_/D vssd1 vssd1 vccd1 vccd1 _09352_/D
+ sky130_fd_sc_hd__and4_1
X_06555_ _06555_/A vssd1 vssd1 vccd1 vccd1 _06555_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09274_ _09284_/D _09276_/C _09206_/X vssd1 vssd1 vccd1 vccd1 _09274_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06486_ _06494_/A _06486_/B _06486_/C vssd1 vssd1 vccd1 vccd1 _06487_/A sky130_fd_sc_hd__or3_1
XFILLER_148_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08225_ _08225_/A _08235_/B _08225_/C vssd1 vssd1 vccd1 vccd1 _08226_/A sky130_fd_sc_hd__or3_1
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07966__A _08004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08156_ _08184_/A _08182_/B _08164_/C vssd1 vssd1 vccd1 vccd1 _08157_/A sky130_fd_sc_hd__or3_1
X_07107_ _07120_/A vssd1 vssd1 vccd1 vccd1 _07118_/B sky130_fd_sc_hd__clkbuf_1
X_08087_ _08101_/A _08101_/B _08087_/C vssd1 vssd1 vccd1 vccd1 _08088_/A sky130_fd_sc_hd__or3_1
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07038_ _07038_/A vssd1 vssd1 vccd1 vccd1 _07038_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11000__B _13944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08989_ _12820_/Q vssd1 vssd1 vccd1 vccd1 _11625_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10951_ _13809_/A _12663_/Q _10955_/S vssd1 vssd1 vccd1 vccd1 _10952_/B sky130_fd_sc_hd__mux2_1
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ _13670_/A _07172_/X vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_8
X_10882_ _10909_/A _10909_/B _10798_/X vssd1 vssd1 vccd1 vccd1 _10883_/B sky130_fd_sc_hd__o21ai_1
XFILLER_43_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12621_ _12646_/CLK _12621_/D vssd1 vssd1 vccd1 vccd1 _12621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _12554_/CLK _12552_/D vssd1 vssd1 vccd1 vccd1 _13680_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11503_ _11680_/A _11503_/B _11503_/C vssd1 vssd1 vccd1 vccd1 _11520_/A sky130_fd_sc_hd__and3_1
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12483_ _12505_/CLK _12483_/D vssd1 vssd1 vccd1 vccd1 _12483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_11434_ _13911_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11434_/X sky130_fd_sc_hd__or2_1
X_13310__466 vssd1 vssd1 vccd1 vccd1 _13310__466/HI _14047_/A sky130_fd_sc_hd__conb_1
XFILLER_137_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_100_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _12404_/CLK sky130_fd_sc_hd__clkbuf_16
X_11365_ _11377_/A _11365_/B vssd1 vssd1 vccd1 vccd1 _11366_/A sky130_fd_sc_hd__and2_1
XFILLER_113_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10316_ _10316_/A vssd1 vssd1 vccd1 vccd1 _12506_/D sky130_fd_sc_hd__clkbuf_1
X_14084_ _14084_/A _08051_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
X_11296_ _10648_/X _11284_/X _11295_/X _11293_/X vssd1 vssd1 vccd1 vccd1 _12747_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10247_ _10688_/C vssd1 vssd1 vccd1 vccd1 _10693_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_140_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10178_ _10191_/A _10178_/B vssd1 vssd1 vccd1 vccd1 _10179_/A sky130_fd_sc_hd__and2_1
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204__360 vssd1 vssd1 vccd1 vccd1 _13204__360/HI _13827_/A sky130_fd_sc_hd__conb_1
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13937_ _13937_/A _06452_/X vssd1 vssd1 vccd1 vccd1 _14065_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13868_ _13868_/A _06647_/X vssd1 vssd1 vccd1 vccd1 _14028_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06955__A _06955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ _12820_/CLK _12819_/D vssd1 vssd1 vccd1 vccd1 _12819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13799_ _13799_/A _06840_/X vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_43_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06340_ _06346_/A _06349_/B _06349_/C vssd1 vssd1 vccd1 vccd1 _06341_/A sky130_fd_sc_hd__or3_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06271_ input5/X vssd1 vssd1 vccd1 vccd1 _11789_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__13788__A _13788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08010_ _08010_/A _08020_/B _08016_/C vssd1 vssd1 vccd1 vccd1 _08011_/A sky130_fd_sc_hd__or3_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ _13595_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09961_/X sky130_fd_sc_hd__or2_1
XFILLER_143_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08912_ _13969_/A vssd1 vssd1 vccd1 vccd1 _09068_/A sky130_fd_sc_hd__clkbuf_1
X_09892_ _10256_/A vssd1 vssd1 vccd1 vccd1 _09892_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater88_A _14028_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__A _09633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08843_ _10162_/B vssd1 vssd1 vccd1 vccd1 _13748_/A sky130_fd_sc_hd__buf_6
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08640__S1 _08576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08774_ _12643_/Q _12644_/Q _12645_/Q _12646_/Q _08766_/X _08767_/X vssd1 vssd1 vccd1
+ vccd1 _08774_/X sky130_fd_sc_hd__mux4_2
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ _07725_/A vssd1 vssd1 vccd1 vccd1 _07725_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07656_ _07739_/A _07863_/B _07739_/C vssd1 vssd1 vccd1 vccd1 _07657_/A sky130_fd_sc_hd__or3_1
XFILLER_80_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06607_ _06607_/A vssd1 vssd1 vccd1 vccd1 _06607_/X sky130_fd_sc_hd__clkbuf_1
X_13253__409 vssd1 vssd1 vccd1 vccd1 _13253__409/HI _13924_/A sky130_fd_sc_hd__conb_1
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07587_ _07615_/A vssd1 vssd1 vccd1 vccd1 _07598_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_34_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09326_ _09324_/X _09372_/B _09326_/C vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__and3b_1
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06538_ _06556_/A _06540_/B _06540_/C vssd1 vssd1 vccd1 vccd1 _06539_/A sky130_fd_sc_hd__or3_1
XFILLER_139_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09257_ _09257_/A _09257_/B vssd1 vssd1 vccd1 vccd1 _12242_/D sky130_fd_sc_hd__nor2_1
X_06469_ _06523_/A vssd1 vssd1 vccd1 vccd1 _06481_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08208_ _08212_/A _08208_/B _08212_/C vssd1 vssd1 vccd1 vccd1 _08209_/A sky130_fd_sc_hd__or3_1
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ _09186_/X _09130_/X _09187_/X _09141_/X vssd1 vssd1 vccd1 vccd1 _12225_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08139_ _08139_/A vssd1 vssd1 vccd1 vccd1 _08139_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11649__C _11649_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11150_ _11127_/Y _11133_/X _11149_/Y _13953_/A vssd1 vssd1 vccd1 vccd1 _11151_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13147__303 vssd1 vssd1 vccd1 vccd1 _13147__303/HI _13704_/A sky130_fd_sc_hd__conb_1
XFILLER_122_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10101_ _10101_/A _10101_/B _10101_/C _10101_/D vssd1 vssd1 vccd1 vccd1 _10112_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_68_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11081_ _13841_/A _12696_/Q _11151_/B vssd1 vssd1 vccd1 vccd1 _11082_/B sky130_fd_sc_hd__mux2_1
XFILLER_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10032_ _10112_/A _10053_/B vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__and2_1
XANTENNA__10879__C1 _10749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input17_A peripheralBus_address[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11983_ _12920_/Q _14063_/A _11995_/S vssd1 vssd1 vccd1 vccd1 _11984_/B sky130_fd_sc_hd__mux2_1
XFILLER_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08839__A2 _08765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__S0 _08368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13722_ _13722_/A _07036_/X vssd1 vssd1 vccd1 vccd1 _13978_/Z sky130_fd_sc_hd__ebufn_8
X_10934_ _12660_/Q _10935_/B vssd1 vssd1 vccd1 vccd1 _10936_/B sky130_fd_sc_hd__or2_1
XFILLER_90_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09151__A _09623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ _13653_/A _07217_/X vssd1 vssd1 vccd1 vccd1 _13973_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_44_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ _10865_/A _10865_/B _10865_/C _10865_/D vssd1 vssd1 vccd1 vccd1 _10866_/D
+ sky130_fd_sc_hd__and4_1
X_12604_ _12813_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__dfxtp_2
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _13584_/A _07409_/X vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_8
X_10796_ _10800_/B _10812_/B _10796_/C vssd1 vssd1 vccd1 vccd1 _10797_/A sky130_fd_sc_hd__and3b_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _12550_/CLK _12535_/D vssd1 vssd1 vccd1 vccd1 _12535_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11071__A2 _11055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13401__A _13401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12466_ _12467_/CLK _12466_/D vssd1 vssd1 vccd1 vccd1 _12466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11417_ _11430_/A vssd1 vssd1 vccd1 vccd1 _11417_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12397_ _12414_/CLK _12397_/D vssd1 vssd1 vccd1 vccd1 _13525_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11348_ _11361_/A _11348_/B vssd1 vssd1 vccd1 vccd1 _11349_/A sky130_fd_sc_hd__and2_1
XFILLER_98_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14067_ _14067_/A _08003_/X vssd1 vssd1 vccd1 vccd1 _14067_/Z sky130_fd_sc_hd__ebufn_8
X_11279_ _11279_/A _11279_/B _11279_/C vssd1 vssd1 vccd1 vccd1 _11279_/Y sky130_fd_sc_hd__nor3_1
XFILLER_140_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12087__A1 _10670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07510_ _07517_/A _07517_/B _07510_/C vssd1 vssd1 vccd1 vccd1 _07511_/A sky130_fd_sc_hd__or3_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08490_ _08486_/X _08489_/X _08528_/S vssd1 vssd1 vccd1 vccd1 _11705_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07441_ _07441_/A vssd1 vssd1 vccd1 vccd1 _07441_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07372_ _07382_/A _07377_/B _07374_/C vssd1 vssd1 vccd1 vccd1 _07373_/A sky130_fd_sc_hd__or3_1
X_09111_ _13628_/Z vssd1 vssd1 vccd1 vccd1 _11064_/A sky130_fd_sc_hd__buf_4
X_06323_ _06333_/A _06323_/B _06323_/C vssd1 vssd1 vccd1 vccd1 _06324_/A sky130_fd_sc_hd__or3_1
XFILLER_148_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09042_ _08932_/X _08933_/X _09015_/X _09041_/X _08924_/X _08925_/X vssd1 vssd1 vccd1
+ vccd1 _09042_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08405__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07947__C _08349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08861__S1 _08808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09944_ _14037_/Z _13589_/A _09953_/S vssd1 vssd1 vccd1 vccd1 _09945_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10670__A _10670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _11412_/B _09875_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _09915_/B sky130_fd_sc_hd__nor3_4
XANTENNA_input9_A peripheralBus_address[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08140__A _11283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _13778_/A vssd1 vssd1 vccd1 vccd1 _08826_/X sky130_fd_sc_hd__buf_2
XFILLER_161_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12078__A1 _11170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ _12642_/Q _12643_/Q _12644_/Q _12645_/Q _08745_/X _08746_/X vssd1 vssd1 vccd1
+ vccd1 _08757_/X sky130_fd_sc_hd__mux4_2
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _07714_/A _07710_/B _07719_/C vssd1 vssd1 vccd1 vccd1 _07709_/A sky130_fd_sc_hd__or3_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _09398_/B vssd1 vssd1 vccd1 vccd1 _13560_/A sky130_fd_sc_hd__buf_4
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _07644_/A _07641_/B _07649_/C vssd1 vssd1 vccd1 vccd1 _07640_/A sky130_fd_sc_hd__or3_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10650_ _10650_/A vssd1 vssd1 vccd1 vccd1 _10650_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11589__B1 _11540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ _09309_/A vssd1 vssd1 vccd1 vccd1 _12255_/D sky130_fd_sc_hd__clkbuf_1
X_10581_ _13718_/A _12574_/Q _10584_/S vssd1 vssd1 vccd1 vccd1 _10582_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12320_ _12320_/CLK _12320_/D vssd1 vssd1 vccd1 vccd1 _12320_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07857__C _07995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08315__A _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ _12251_/CLK _12251_/D vssd1 vssd1 vccd1 vccd1 _12251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11202_ _11254_/S vssd1 vssd1 vccd1 vccd1 _11281_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_107_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12182_ _12195_/A vssd1 vssd1 vccd1 vccd1 _12182_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11133_ _11128_/Y _11129_/X _11130_/Y _11131_/X _11132_/Y vssd1 vssd1 vccd1 vccd1
+ _11133_/X sky130_fd_sc_hd__o221a_1
XFILLER_122_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09146__A _09146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ _11064_/A vssd1 vssd1 vccd1 vccd1 _11064_/X sky130_fd_sc_hd__buf_6
XFILLER_95_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08604__S1 _08603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _10015_/A vssd1 vssd1 vccd1 vccd1 _12432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12069__A1 _10645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11966_ _11978_/A _11966_/B vssd1 vssd1 vccd1 vccd1 _11967_/A sky130_fd_sc_hd__and2_1
X_13275__431 vssd1 vssd1 vccd1 vccd1 _13275__431/HI _13966_/A sky130_fd_sc_hd__conb_1
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10917_ _10915_/X _10917_/B _10917_/C vssd1 vssd1 vccd1 vccd1 _10918_/A sky130_fd_sc_hd__and3b_1
XFILLER_72_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13705_ _13705_/A _07077_/X vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11897_ _11897_/A vssd1 vssd1 vccd1 vccd1 _12901_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13636_ _13636_/A _07264_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
X_10848_ _10875_/B _10875_/C _10848_/C vssd1 vssd1 vccd1 vccd1 _10854_/C sky130_fd_sc_hd__and3_1
XFILLER_158_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13316__472 vssd1 vssd1 vccd1 vccd1 _13316__472/HI _14053_/A sky130_fd_sc_hd__conb_1
X_13567_ _13567_/A _07451_/X vssd1 vssd1 vccd1 vccd1 _14111_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_12_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10779_ _12623_/Q vssd1 vssd1 vccd1 vccd1 _10865_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_158_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12518_ _12522_/CLK _12518_/D vssd1 vssd1 vccd1 vccd1 _13647_/A sky130_fd_sc_hd__dfxtp_1
X_13498_ _13498_/A _07627_/X vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_8
X_12449_ _12457_/CLK _12449_/D vssd1 vssd1 vccd1 vccd1 _12449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _14119_/A _08260_/X vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__ebufn_8
X_07990_ _07990_/A vssd1 vssd1 vccd1 vccd1 _07990_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06941_ _06948_/A _06941_/B vssd1 vssd1 vccd1 vccd1 _06942_/A sky130_fd_sc_hd__or2_1
X_09660_ _09669_/A _09660_/B vssd1 vssd1 vccd1 vccd1 _09661_/A sky130_fd_sc_hd__and2_1
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06872_ _06900_/A vssd1 vssd1 vccd1 vccd1 _06884_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_55_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08611_ _12435_/Q vssd1 vssd1 vccd1 vccd1 _10029_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09591_ _12321_/Q _13564_/A vssd1 vssd1 vccd1 vccd1 _09591_/Y sky130_fd_sc_hd__xnor2_1
X_08542_ _12272_/Q vssd1 vssd1 vccd1 vccd1 _09388_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08473_ _11705_/A vssd1 vssd1 vccd1 vccd1 _13363_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07424_ _07424_/A vssd1 vssd1 vccd1 vccd1 _07424_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07355_ _07355_/A vssd1 vssd1 vccd1 vccd1 _07355_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10665__A _10665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06306_ _09125_/A vssd1 vssd1 vccd1 vccd1 _06361_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07286_ _07292_/A _07289_/B _07286_/C vssd1 vssd1 vccd1 vccd1 _07287_/A sky130_fd_sc_hd__or3_1
XANTENNA__08135__A _08135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09025_ _08969_/X _08972_/X _08970_/X _08975_/X _09024_/X _09013_/X vssd1 vssd1 vccd1
+ vccd1 _09025_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11496__A _13979_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _09982_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _09927_/X sky130_fd_sc_hd__or2_1
XFILLER_120_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09858_ _09858_/A _09858_/B _09858_/C _09858_/D vssd1 vssd1 vccd1 vccd1 _09869_/A
+ sky130_fd_sc_hd__or4_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08809_ _10864_/A _10874_/C _10874_/B _12632_/Q _08807_/X _08808_/X vssd1 vssd1 vccd1
+ vccd1 _08809_/X sky130_fd_sc_hd__mux4_2
XFILLER_45_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09789_ hold2/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09789_/X sky130_fd_sc_hd__or2_1
XFILLER_105_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13259__415 vssd1 vssd1 vccd1 vccd1 _13259__415/HI _13930_/A sky130_fd_sc_hd__conb_1
XFILLER_39_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _09636_/A _14007_/A _11823_/S vssd1 vssd1 vccd1 vccd1 _11821_/B sky130_fd_sc_hd__mux2_1
XFILLER_61_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11757_/A _11751_/B vssd1 vssd1 vccd1 vccd1 _11752_/A sky130_fd_sc_hd__and2_1
XFILLER_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_80_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _12625_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ input27/X vssd1 vssd1 vccd1 vccd1 _10720_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11680_/X _11682_/B _11682_/C vssd1 vssd1 vccd1 vccd1 _11683_/A sky130_fd_sc_hd__and3b_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13421_/A _07836_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
X_10633_ _10633_/A _10633_/B _10633_/C vssd1 vssd1 vccd1 vccd1 _10633_/Y sky130_fd_sc_hd__nor3_1
XFILLER_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10564_ _10567_/A _10564_/B vssd1 vssd1 vccd1 vccd1 _10565_/A sky130_fd_sc_hd__and2_1
X_12303_ _12331_/CLK _12303_/D vssd1 vssd1 vccd1 vccd1 _13434_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10495_ _12549_/Q _13758_/A vssd1 vssd1 vccd1 vccd1 _10499_/A sky130_fd_sc_hd__xor2_1
XFILLER_154_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12234_ _12289_/CLK _12234_/D vssd1 vssd1 vccd1 vccd1 _12234_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10537__A1 _09773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08825__S1 _08808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12165_ _12967_/Q _13373_/A vssd1 vssd1 vccd1 vccd1 _12166_/D sky130_fd_sc_hd__xor2_1
XFILLER_122_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater119_A peripheralBus_data[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11116_ _11204_/A _11116_/B vssd1 vssd1 vccd1 vccd1 _11117_/A sky130_fd_sc_hd__and2_1
XFILLER_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12096_ _14076_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__or2_1
XFILLER_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11047_ _13814_/A _11051_/B vssd1 vssd1 vccd1 vccd1 _11047_/X sky130_fd_sc_hd__or2_1
XANTENNA__11498__C1 _11497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 peripheralBus_address[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output48_A _13952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09002__S1 _08968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11949_ _11962_/A _11949_/B vssd1 vssd1 vccd1 vccd1 _11950_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_71_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _12533_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _13619_/A _07311_/X vssd1 vssd1 vccd1 vccd1 _14099_/Z sky130_fd_sc_hd__ebufn_8
X_13052__208 vssd1 vssd1 vccd1 vccd1 _13052__208/HI _13511_/A sky130_fd_sc_hd__conb_1
X_07140_ _07152_/A _07145_/B _07142_/C vssd1 vssd1 vccd1 vccd1 _07141_/A sky130_fd_sc_hd__or3_1
XFILLER_118_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07071_ _07079_/A _07076_/B _07073_/C vssd1 vssd1 vccd1 vccd1 _07072_/A sky130_fd_sc_hd__or3_1
XFILLER_145_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10528__A1 _10394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07973_ _08075_/A _08075_/B _07977_/C vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__or3_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09712_ _09800_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09713_/A sky130_fd_sc_hd__and2_1
XFILLER_101_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06924_ _06924_/A vssd1 vssd1 vccd1 vccd1 _06924_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater70_A peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ _13465_/A _09640_/X _09642_/X _09634_/X vssd1 vssd1 vccd1 vccd1 _12335_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06855_ _06863_/A _06857_/B _06857_/C vssd1 vssd1 vccd1 vccd1 _06856_/A sky130_fd_sc_hd__or3_1
XANTENNA__07960__C _07962_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09574_ _09574_/A vssd1 vssd1 vccd1 vccd1 _12320_/D sky130_fd_sc_hd__clkbuf_1
X_06786_ _06788_/A _06793_/B _06793_/C vssd1 vssd1 vccd1 vccd1 _06787_/A sky130_fd_sc_hd__or3_1
XFILLER_83_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _08525_/A vssd1 vssd1 vccd1 vccd1 _09146_/A sky130_fd_sc_hd__buf_2
XFILLER_24_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07034__A _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_62_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _12811_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_60_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ _12255_/Q vssd1 vssd1 vccd1 vccd1 _09330_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__07969__A _08089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06873__A _07248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07407_ _08084_/A vssd1 vssd1 vccd1 vccd1 _07840_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12205__A1 _10670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ _12250_/Q vssd1 vssd1 vccd1 vccd1 _09321_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10395__A _10409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07338_ _07406_/A vssd1 vssd1 vccd1 vccd1 _07393_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_75_clk_A _12555_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11003__B _13936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ _07279_/A _07276_/B _07273_/C vssd1 vssd1 vccd1 vccd1 _07270_/A sky130_fd_sc_hd__or3_1
X_09008_ _11649_/A _11657_/C _11657_/B _11661_/B _08946_/X _08947_/X vssd1 vssd1 vccd1
+ vccd1 _09008_/X sky130_fd_sc_hd__mux4_2
X_10280_ _13625_/A _10291_/B vssd1 vssd1 vccd1 vccd1 _10280_/X sky130_fd_sc_hd__or2_1
XANTENNA__10519__A1 _09750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10842__B _10917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09137__A1 _09124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13970_ _13970_/A _06368_/X vssd1 vssd1 vccd1 vccd1 _14066_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA_clkbuf_leaf_13_clk_A _12217_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09424__A _11408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ _12923_/CLK _12921_/D vssd1 vssd1 vccd1 vccd1 _12921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08991__S0 _08911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ _12853_/CLK _12852_/D vssd1 vssd1 vccd1 vccd1 _12852_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _11816_/A _11803_/B vssd1 vssd1 vccd1 vccd1 _11804_/A sky130_fd_sc_hd__and2_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12786_/CLK _12783_/D vssd1 vssd1 vccd1 vccd1 _13909_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_28_clk_A _12759_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _12853_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07879__A _07892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11734_ _11740_/A _11734_/B vssd1 vssd1 vccd1 vccd1 _11735_/A sky130_fd_sc_hd__and2_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06783__A _06809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _11665_/A _11667_/B vssd1 vssd1 vccd1 vccd1 _12843_/D sky130_fd_sc_hd__nor2_1
XFILLER_159_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_clk clkbuf_4_7_0_clk/A vssd1 vssd1 vccd1 vccd1 _12555_/CLK sky130_fd_sc_hd__clkbuf_2
X_13404_ _13404_/A _07974_/X vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_8
X_10616_ _12580_/Q _13756_/A vssd1 vssd1 vccd1 vccd1 _10616_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11596_ _11632_/B _11590_/A _11632_/A vssd1 vssd1 vccd1 vccd1 _11597_/C sky130_fd_sc_hd__a21o_1
XFILLER_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10547_ _10288_/X _10538_/X _10546_/X _10536_/X vssd1 vssd1 vccd1 vccd1 _12564_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10478_ _10478_/A vssd1 vssd1 vccd1 vccd1 _12548_/D sky130_fd_sc_hd__clkbuf_1
X_12217_ _12217_/CLK _12217_/D vssd1 vssd1 vccd1 vccd1 _13394_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11183__A1 _10670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ _12966_/Q _14108_/A _12151_/S vssd1 vssd1 vccd1 vccd1 _12149_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11864__A _11898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12079_ _14069_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12079_/X sky130_fd_sc_hd__or2_1
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06640_ _11156_/B vssd1 vssd1 vccd1 vccd1 _08184_/B sky130_fd_sc_hd__buf_6
XFILLER_65_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06571_ _06599_/A vssd1 vssd1 vccd1 vccd1 _06584_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _12589_/CLK sky130_fd_sc_hd__clkbuf_16
X_08310_ _08310_/A vssd1 vssd1 vccd1 vccd1 _08310_/X sky130_fd_sc_hd__clkbuf_1
X_09290_ _09330_/D _09292_/C _09392_/A vssd1 vssd1 vccd1 vccd1 _09290_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12995__151 vssd1 vssd1 vccd1 vccd1 _12995__151/HI _13406_/A sky130_fd_sc_hd__conb_1
X_08241_ _08351_/A vssd1 vssd1 vccd1 vccd1 _08251_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__11104__A _11124_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ _08174_/A _08174_/B _08184_/C vssd1 vssd1 vccd1 vccd1 _08173_/A sky130_fd_sc_hd__or3_1
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07123_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07135_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10943__A _13980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09509__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07054_ _07054_/A vssd1 vssd1 vccd1 vccd1 _07054_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11174__A1 _11170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13180__336 vssd1 vssd1 vccd1 vccd1 _13180__336/HI _13773_/A sky130_fd_sc_hd__conb_1
X_07956_ _07962_/A _07962_/B _07993_/C vssd1 vssd1 vccd1 vccd1 _07957_/A sky130_fd_sc_hd__or3_1
X_06907_ _08168_/A _06916_/B vssd1 vssd1 vccd1 vccd1 _06908_/A sky130_fd_sc_hd__or2_1
X_07887_ _07887_/A vssd1 vssd1 vccd1 vccd1 _07887_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09626_ _13459_/A _09613_/X _09625_/X _09621_/X vssd1 vssd1 vccd1 vccd1 _12329_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06838_ _06879_/A vssd1 vssd1 vccd1 vccd1 _06850_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13221__377 vssd1 vssd1 vccd1 vccd1 _13221__377/HI _13860_/A sky130_fd_sc_hd__conb_1
XFILLER_71_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09557_ _09557_/A vssd1 vssd1 vccd1 vccd1 _12315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06769_ _06832_/A vssd1 vssd1 vccd1 vccd1 _06780_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _12724_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08508_ _08430_/X _08431_/X _08482_/X _08507_/X _08492_/X _08449_/X vssd1 vssd1 vccd1
+ vccd1 _08508_/X sky130_fd_sc_hd__mux4_1
X_09488_ _11160_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _09488_/X sky130_fd_sc_hd__or2_1
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08439_ _09316_/C _12236_/Q _09317_/C _09258_/D _08417_/X _08418_/X vssd1 vssd1 vccd1
+ vccd1 _08439_/X sky130_fd_sc_hd__mux4_2
X_13074__230 vssd1 vssd1 vccd1 vccd1 _13074__230/HI _13549_/A sky130_fd_sc_hd__conb_1
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11450_ _13917_/A _11450_/B vssd1 vssd1 vccd1 vccd1 _11450_/X sky130_fd_sc_hd__or2_1
XANTENNA__11937__A0 _09623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10401_ _09763_/X _10395_/X _10400_/X _10398_/X vssd1 vssd1 vccd1 vccd1 _12524_/D
+ sky130_fd_sc_hd__o211a_1
X_11381_ _13918_/A _12775_/Q _11381_/S vssd1 vssd1 vccd1 vccd1 _11382_/B sky130_fd_sc_hd__mux2_1
X_13115__271 vssd1 vssd1 vccd1 vccd1 _13115__271/HI _13640_/A sky130_fd_sc_hd__conb_1
XFILLER_125_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ _10332_/A _10332_/B vssd1 vssd1 vccd1 vccd1 _10333_/A sky130_fd_sc_hd__and2_1
XANTENNA__08323__A _08335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ _09756_/X _10249_/X _10262_/X _10256_/X vssd1 vssd1 vccd1 vccd1 _12489_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12002_ _12002_/A vssd1 vssd1 vccd1 vccd1 _12925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10194_ _13622_/A _12475_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _10195_/B sky130_fd_sc_hd__mux2_1
XFILLER_87_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09154__A _14067_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13953_ _13953_/A _06413_/X vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__ebufn_8
X_12904_ _12904_/CLK _12904_/D vssd1 vssd1 vccd1 vccd1 _14031_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13884_ _13884_/A _06601_/X vssd1 vssd1 vccd1 vccd1 _14012_/Z sky130_fd_sc_hd__ebufn_8
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _12835_/CLK _12835_/D vssd1 vssd1 vccd1 vccd1 _12835_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk _12881_/CLK vssd1 vssd1 vccd1 vccd1 _12775_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13404__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09601__B _13558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12786_/CLK _12766_/D vssd1 vssd1 vccd1 vccd1 _12766_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11723_/A _11717_/B vssd1 vssd1 vccd1 vccd1 _11718_/A sky130_fd_sc_hd__and2_1
X_12697_ _12704_/CLK _12697_/D vssd1 vssd1 vccd1 vccd1 _12697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11648_ _11648_/A vssd1 vssd1 vccd1 vccd1 _12838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 peripheralBus_address[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 peripheralBus_address[8] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
X_11579_ _13967_/A _11639_/B _11632_/D _11649_/C vssd1 vssd1 vccd1 vccd1 _11602_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07810_ _07810_/A vssd1 vssd1 vccd1 vccd1 _07810_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08790_ _12632_/Q _12633_/Q _12634_/Q _10870_/A _08785_/X _08786_/X vssd1 vssd1 vccd1
+ vccd1 _08790_/X sky130_fd_sc_hd__mux4_2
XANTENNA__06688__A _06688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07741_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07753_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_65_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07672_ _07672_/A _07683_/B _07678_/C vssd1 vssd1 vccd1 vccd1 _07673_/A sky130_fd_sc_hd__or3_1
X_09411_ _13425_/A _12277_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _09412_/B sky130_fd_sc_hd__mux2_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06623_ _06625_/A _06630_/B _06630_/C vssd1 vssd1 vccd1 vccd1 _06624_/A sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_17_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _12952_/CLK sky130_fd_sc_hd__clkbuf_16
X_13058__214 vssd1 vssd1 vccd1 vccd1 _13058__214/HI _13517_/A sky130_fd_sc_hd__conb_1
X_09342_ _12261_/Q vssd1 vssd1 vccd1 vccd1 _09352_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_06554_ _06556_/A _06561_/B _06561_/C vssd1 vssd1 vccd1 vccd1 _06555_/A sky130_fd_sc_hd__or3_1
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09273_ _09321_/D vssd1 vssd1 vccd1 vccd1 _09284_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_06485_ _06485_/A vssd1 vssd1 vccd1 vccd1 _06485_/X sky130_fd_sc_hd__clkbuf_1
X_08224_ _08263_/A vssd1 vssd1 vccd1 vccd1 _08235_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_21_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08155_ _08155_/A vssd1 vssd1 vccd1 vccd1 _08155_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07106_ _07106_/A vssd1 vssd1 vccd1 vccd1 _07106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08086_ _08086_/A vssd1 vssd1 vccd1 vccd1 _08086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07037_ _07043_/A _07043_/B vssd1 vssd1 vccd1 vccd1 _07038_/A sky130_fd_sc_hd__or2_1
XFILLER_161_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07982__A _08004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08988_ _12819_/Q vssd1 vssd1 vccd1 vccd1 _11625_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07939_ _07951_/A _07945_/B _07945_/C vssd1 vssd1 vccd1 vccd1 _07940_/A sky130_fd_sc_hd__or3_1
XFILLER_113_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10950_ _10950_/A vssd1 vssd1 vccd1 vccd1 _12662_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09609_ _09586_/Y _09592_/X _09608_/Y _13569_/A vssd1 vssd1 vccd1 vccd1 _09610_/C
+ sky130_fd_sc_hd__a31o_1
X_10881_ _10881_/A _10881_/B _10881_/C vssd1 vssd1 vccd1 vccd1 _10909_/B sky130_fd_sc_hd__and3_1
XFILLER_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12620_ _12660_/CLK _12620_/D vssd1 vssd1 vccd1 vccd1 _12620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07222__A _07533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ _12565_/CLK _12551_/D vssd1 vssd1 vccd1 vccd1 _13679_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11502_ _13976_/A _13975_/A _11501_/X vssd1 vssd1 vccd1 vccd1 _11503_/C sky130_fd_sc_hd__or3b_1
XANTENNA__10830__B1 _10803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12482_ _12505_/CLK _12482_/D vssd1 vssd1 vccd1 vccd1 _12482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11433_ _10662_/X _11425_/X _11432_/X _11430_/X vssd1 vssd1 vccd1 vccd1 _12784_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11398__B _13947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11364_ _13913_/A _12770_/Q _11373_/S vssd1 vssd1 vccd1 vccd1 _11365_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10315_ _10315_/A _10315_/B vssd1 vssd1 vccd1 vccd1 _10316_/A sky130_fd_sc_hd__and2_1
XFILLER_98_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14083_ _14083_/A _08048_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11295_ _13874_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11295_/X sky130_fd_sc_hd__or2_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07892__A _07892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10246_ input7/X _11789_/C _11789_/D input5/X vssd1 vssd1 vccd1 vccd1 _10688_/C sky130_fd_sc_hd__or4b_4
XFILLER_112_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater101_A peripheralBus_data[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ _13617_/A _12470_/Q _10180_/S vssd1 vssd1 vccd1 vccd1 _10178_/B sky130_fd_sc_hd__mux2_1
XFILLER_121_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13936_ _13936_/A _06454_/X vssd1 vssd1 vccd1 vccd1 _14064_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_35_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output30_A _13788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__A _11154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13867_ _13867_/A _06650_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
X_12818_ _12829_/CLK _12818_/D vssd1 vssd1 vccd1 vccd1 _12818_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08228__A _08228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13798_ _13798_/A _06842_/X vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11074__A0 _13839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12768_/CLK _12749_/D vssd1 vssd1 vccd1 vccd1 _13876_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06270_ _08364_/A vssd1 vssd1 vccd1 vccd1 _07827_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09960_ _09186_/X _09921_/X _09958_/X _09959_/X vssd1 vssd1 vccd1 vccd1 _12418_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_6_clk _12917_/CLK vssd1 vssd1 vccd1 vccd1 _12919_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ _09067_/A vssd1 vssd1 vccd1 vccd1 _08911_/X sky130_fd_sc_hd__buf_4
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _10667_/A vssd1 vssd1 vccd1 vccd1 _10256_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10940__B _11384_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _08839_/X _08841_/X _08863_/S vssd1 vssd1 vccd1 vccd1 _10162_/B sky130_fd_sc_hd__mux2_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _12639_/Q _12640_/Q _12641_/Q _12642_/Q _08766_/X _08767_/X vssd1 vssd1 vccd1
+ vccd1 _08773_/X sky130_fd_sc_hd__mux4_2
XFILLER_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07724_ _07727_/A _07724_/B _07732_/C vssd1 vssd1 vccd1 vccd1 _07725_/A sky130_fd_sc_hd__or3_1
XFILLER_38_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09522__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ _07655_/A vssd1 vssd1 vccd1 vccd1 _07655_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11771__B _13362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10668__A _11039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ _06610_/A _06616_/B _06616_/C vssd1 vssd1 vccd1 vccd1 _06607_/A sky130_fd_sc_hd__or3_1
XFILLER_53_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07586_ _07586_/A vssd1 vssd1 vccd1 vccd1 _07586_/X sky130_fd_sc_hd__clkbuf_1
X_13292__448 vssd1 vssd1 vccd1 vccd1 _13292__448/HI _13997_/A sky130_fd_sc_hd__conb_1
XFILLER_80_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09325_ _09329_/A _09312_/B _09328_/A vssd1 vssd1 vccd1 vccd1 _09326_/C sky130_fd_sc_hd__a21o_1
X_06537_ _06599_/A vssd1 vssd1 vccd1 vccd1 _06556_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13979__A _13979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ _09316_/B _09256_/B vssd1 vssd1 vccd1 vccd1 _09257_/B sky130_fd_sc_hd__and2_1
X_06468_ _06688_/A vssd1 vssd1 vccd1 vccd1 _06523_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13333__489 vssd1 vssd1 vccd1 vccd1 _13333__489/HI _14086_/A sky130_fd_sc_hd__conb_1
X_08207_ _08207_/A vssd1 vssd1 vccd1 vccd1 _08207_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11499__A _14012_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09187_ _13402_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__or2_1
X_06399_ _06399_/A vssd1 vssd1 vccd1 vccd1 _06399_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08138_ _08148_/A _08189_/B _08138_/C vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__or3_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08069_ _08069_/A vssd1 vssd1 vccd1 vccd1 _08069_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13186__342 vssd1 vssd1 vccd1 vccd1 _13186__342/HI _13793_/A sky130_fd_sc_hd__conb_1
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10100_ _10100_/A _10100_/B _10100_/C _10100_/D vssd1 vssd1 vccd1 vccd1 _10101_/D
+ sky130_fd_sc_hd__and4_1
X_11080_ _11206_/A vssd1 vssd1 vccd1 vccd1 _11095_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08536__A2 _08427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ _10101_/C vssd1 vssd1 vccd1 vccd1 _10053_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13227__383 vssd1 vssd1 vccd1 vccd1 _13227__383/HI _13866_/A sky130_fd_sc_hd__conb_1
XFILLER_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11982_ _12033_/S vssd1 vssd1 vccd1 vccd1 _11995_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08395__S1 _08370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ _13721_/A _07038_/X vssd1 vssd1 vccd1 vccd1 _14105_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_17_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10933_ _10933_/A _10935_/B vssd1 vssd1 vccd1 vccd1 _12659_/D sky130_fd_sc_hd__nor2_1
XFILLER_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09249__B1 _09248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ _10864_/A _10864_/B _10864_/C _10864_/D vssd1 vssd1 vccd1 vccd1 _10866_/C
+ sky130_fd_sc_hd__and4_1
X_13652_ _13652_/A _07221_/X vssd1 vssd1 vccd1 vccd1 _14100_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _12813_/CLK _12603_/D vssd1 vssd1 vccd1 vccd1 _13778_/A sky130_fd_sc_hd__dfxtp_2
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _13583_/A _08076_/X vssd1 vssd1 vccd1 vccd1 _13775_/Z sky130_fd_sc_hd__ebufn_8
X_10795_ _10863_/B _10795_/B vssd1 vssd1 vccd1 vccd1 _10796_/C sky130_fd_sc_hd__or2_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09578__S _09582_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12550_/CLK _12534_/D vssd1 vssd1 vccd1 vccd1 _12534_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12465_ _12467_/CLK _12465_/D vssd1 vssd1 vccd1 vccd1 _12465_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11202__A _11254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ _13904_/A _11423_/B vssd1 vssd1 vccd1 vccd1 _11416_/X sky130_fd_sc_hd__or2_1
X_12396_ _12418_/CLK _12396_/D vssd1 vssd1 vccd1 vccd1 _13524_/A sky130_fd_sc_hd__dfxtp_1
X_11347_ _13908_/A _12765_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _11348_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11278_ _11278_/A _11278_/B _11278_/C _11278_/D vssd1 vssd1 vccd1 vccd1 _11279_/C
+ sky130_fd_sc_hd__or4_1
X_14066_ _14066_/A _08001_/X vssd1 vssd1 vccd1 vccd1 _14066_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10229_ _12474_/Q _13749_/A vssd1 vssd1 vccd1 vccd1 _10232_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09326__B _09372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13919_ _13919_/A _06504_/X vssd1 vssd1 vccd1 vccd1 _14079_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07440_ _07442_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07441_/A sky130_fd_sc_hd__or2_1
XFILLER_62_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13020__176 vssd1 vssd1 vccd1 vccd1 _13020__176/HI _13447_/A sky130_fd_sc_hd__conb_1
X_07371_ _07371_/A vssd1 vssd1 vccd1 vccd1 _07382_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09110_ _09092_/X _09100_/X _09104_/X _09109_/X vssd1 vssd1 vccd1 vccd1 _12210_/D
+ sky130_fd_sc_hd__o211a_1
X_06322_ _06361_/A vssd1 vssd1 vccd1 vccd1 _06333_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_31_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09041_ _12843_/Q _12844_/Q _12845_/Q _12846_/Q _08946_/X _08947_/X vssd1 vssd1 vccd1
+ vccd1 _09041_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09517__A _11189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09943_ _11490_/A vssd1 vssd1 vccd1 vccd1 _10700_/A sky130_fd_sc_hd__buf_2
XANTENNA__11766__B _13368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09176__C1 _09939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _09902_/A vssd1 vssd1 vccd1 vccd1 _09874_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08825_ _10909_/A _12646_/Q _10908_/B _10908_/A _08807_/X _08808_/X vssd1 vssd1 vccd1
+ vccd1 _08825_/X sky130_fd_sc_hd__mux4_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08756_ _12638_/Q _12639_/Q _10876_/B _12641_/Q _08742_/X _08743_/X vssd1 vssd1 vccd1
+ vccd1 _08756_/X sky130_fd_sc_hd__mux4_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _07763_/A vssd1 vssd1 vccd1 vccd1 _07719_/C sky130_fd_sc_hd__clkbuf_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08687_ _08684_/X _08686_/X _08712_/S vssd1 vssd1 vccd1 vccd1 _09398_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07638_ _07693_/A vssd1 vssd1 vccd1 vccd1 _07649_/C sky130_fd_sc_hd__clkbuf_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07569_ _07569_/A vssd1 vssd1 vccd1 vccd1 _07569_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09308_ _09312_/B _09372_/B _09308_/C vssd1 vssd1 vccd1 vccd1 _09309_/A sky130_fd_sc_hd__and3b_1
XFILLER_70_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10580_ _10580_/A vssd1 vssd1 vccd1 vccd1 _12573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10261__A1 _09753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09239_ _09258_/D vssd1 vssd1 vccd1 vccd1 _09317_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12250_ _12251_/CLK _12250_/D vssd1 vssd1 vccd1 vccd1 _12250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11201_ _13978_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11254_/S sky130_fd_sc_hd__and2_4
XFILLER_5_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12181_ _11153_/X _09100_/X _12180_/X _12097_/X vssd1 vssd1 vccd1 vccd1 _12970_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11132_ _12705_/Q _13946_/A vssd1 vssd1 vccd1 vccd1 _11132_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_162_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11063_ _11061_/X _11055_/X _11062_/X _11053_/X vssd1 vssd1 vccd1 vccd1 _12690_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08050__B _08110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10014_ _10160_/A _10014_/B vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__and2_1
XFILLER_135_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11965_ _14106_/Z _14042_/A _11974_/S vssd1 vssd1 vccd1 vccd1 _11966_/B sky130_fd_sc_hd__mux2_1
XFILLER_151_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13704_ _13704_/A _07080_/X vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _10885_/A _10915_/C _10921_/C vssd1 vssd1 vccd1 vccd1 _10917_/C sky130_fd_sc_hd__a21o_1
XFILLER_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11896_ _11927_/A _11896_/B vssd1 vssd1 vccd1 vccd1 _11897_/A sky130_fd_sc_hd__and2_1
X_13635_ _13635_/A _07267_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10847_ _10847_/A _10847_/B vssd1 vssd1 vccd1 vccd1 _12638_/D sky130_fd_sc_hd__nor2_1
XFILLER_158_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13566_ _13566_/A _07453_/X vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ _10778_/A vssd1 vssd1 vccd1 vccd1 _12622_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07410__A _09918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12517_ _12517_/CLK _12517_/D vssd1 vssd1 vccd1 vccd1 _13761_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_157_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13497_ _13497_/A _07631_/X vssd1 vssd1 vccd1 vccd1 _13625_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_157_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ _12451_/CLK _12448_/D vssd1 vssd1 vccd1 vccd1 _12448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12379_ _12386_/CLK _12379_/D vssd1 vssd1 vccd1 vccd1 _12379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14118_ _14118_/A _08258_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[23] sky130_fd_sc_hd__ebufn_8
XFILLER_141_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08241__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10490__B _13753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06940_ _06940_/A vssd1 vssd1 vccd1 vccd1 _06940_/X sky130_fd_sc_hd__clkbuf_1
X_14049_ _14049_/A _07912_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_79_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06871_ _06871_/A vssd1 vssd1 vccd1 vccd1 _06871_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08610_ _10021_/D _12432_/Q _10021_/B _10024_/B _08575_/X _08576_/X vssd1 vssd1 vccd1
+ vccd1 _08610_/X sky130_fd_sc_hd__mux4_2
X_09590_ _12309_/Q _09851_/B vssd1 vssd1 vccd1 vccd1 _09590_/X sky130_fd_sc_hd__and2_1
XANTENNA__06696__A _06722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08541_ _08447_/X _08452_/X _08455_/X _08458_/X _08467_/X _09157_/A vssd1 vssd1 vccd1
+ vccd1 _08541_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08472_ _08468_/X _08471_/X _13396_/A vssd1 vssd1 vccd1 vccd1 _11705_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07423_ _07430_/A _07423_/B vssd1 vssd1 vccd1 vccd1 _07424_/A sky130_fd_sc_hd__or2_1
XANTENNA__10946__A _10952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07354_ _07356_/A _07364_/B _07361_/C vssd1 vssd1 vccd1 vccd1 _07355_/A sky130_fd_sc_hd__or3_1
XANTENNA__07958__C _07962_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07320__A _09918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06305_ _11457_/A vssd1 vssd1 vccd1 vccd1 _09125_/A sky130_fd_sc_hd__buf_6
X_07285_ _07285_/A vssd1 vssd1 vccd1 vccd1 _07285_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08135__B _08189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ _13971_/A vssd1 vssd1 vccd1 vccd1 _09024_/X sky130_fd_sc_hd__buf_2
XFILLER_163_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09926_ _09963_/B vssd1 vssd1 vccd1 vccd1 _09958_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_86_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _12388_/Q _13565_/A vssd1 vssd1 vccd1 vccd1 _09858_/D sky130_fd_sc_hd__xor2_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08808_ _08887_/A vssd1 vssd1 vccd1 vccd1 _08808_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09788_ _09116_/X _09776_/X _09787_/X _09781_/X vssd1 vssd1 vccd1 vccd1 _12372_/D
+ sky130_fd_sc_hd__o211a_1
X_13298__454 vssd1 vssd1 vccd1 vccd1 _13298__454/HI _14019_/A sky130_fd_sc_hd__conb_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08739_ _08886_/A vssd1 vssd1 vccd1 vccd1 _08739_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _12865_/Q _14010_/A _11760_/S vssd1 vssd1 vccd1 vccd1 _11751_/B sky130_fd_sc_hd__mux2_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13339__495 vssd1 vssd1 vccd1 vccd1 _13339__495/HI _14092_/A sky130_fd_sc_hd__conb_1
X_10701_ _10701_/A vssd1 vssd1 vccd1 vccd1 _12602_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11681_ _11658_/A _11680_/C _11687_/C vssd1 vssd1 vccd1 vccd1 _11682_/C sky130_fd_sc_hd__a21o_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13420_/A _07834_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10632_ _10632_/A _10632_/B _10632_/C _10632_/D vssd1 vssd1 vccd1 vccd1 _10633_/C
+ sky130_fd_sc_hd__or4_1
XANTENNA__08326__A _08338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10563_ _13713_/A _12569_/Q _10635_/B vssd1 vssd1 vccd1 vccd1 _10564_/B sky130_fd_sc_hd__mux2_1
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12302_ _12331_/CLK _12302_/D vssd1 vssd1 vccd1 vccd1 _13433_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _10494_/A _10494_/B _10494_/C _10494_/D vssd1 vssd1 vccd1 vccd1 _10505_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12233_ _12289_/CLK _12233_/D vssd1 vssd1 vccd1 vccd1 _12233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12164_ _12963_/Q _13369_/A vssd1 vssd1 vccd1 vccd1 _12166_/C sky130_fd_sc_hd__xor2_1
XFILLER_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _13851_/A _12706_/Q _11118_/S vssd1 vssd1 vccd1 vccd1 _11116_/B sky130_fd_sc_hd__mux2_1
XFILLER_150_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12095_ _11061_/X _12088_/X _12094_/X _12084_/X vssd1 vssd1 vccd1 vccd1 _12949_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11046_ _10659_/X _11041_/X _11045_/X _11039_/X vssd1 vssd1 vccd1 vccd1 _12684_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09604__B _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11948_ _09631_/A _14037_/A _11957_/S vssd1 vssd1 vccd1 vccd1 _11949_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09620__A _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ _11886_/A _11879_/B vssd1 vssd1 vccd1 vccd1 _11880_/A sky130_fd_sc_hd__and2_1
X_13618_ _13618_/A _07313_/X vssd1 vssd1 vccd1 vccd1 _14098_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10485__B _10613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13091__247 vssd1 vssd1 vccd1 vccd1 _13091__247/HI _13600_/A sky130_fd_sc_hd__conb_1
X_13549_ _13549_/A _07491_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07070_ _07070_/A vssd1 vssd1 vccd1 vccd1 _07070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132__288 vssd1 vssd1 vccd1 vccd1 _13132__288/HI _13673_/A sky130_fd_sc_hd__conb_1
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07972_ _07972_/A vssd1 vssd1 vccd1 vccd1 _07972_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09711_ hold2/A _12356_/Q _09711_/S vssd1 vssd1 vccd1 vccd1 _09712_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11489__A0 _13976_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06923_ _06923_/A _06929_/B vssd1 vssd1 vccd1 vccd1 _06924_/A sky130_fd_sc_hd__or2_1
XFILLER_28_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09642_ _11184_/A _09653_/B vssd1 vssd1 vccd1 vccd1 _09642_/X sky130_fd_sc_hd__or2_1
X_06854_ _06854_/A vssd1 vssd1 vccd1 vccd1 _06854_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13026__182 vssd1 vssd1 vccd1 vccd1 _13026__182/HI _13453_/A sky130_fd_sc_hd__conb_1
XANTENNA_repeater63_A _13623_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06785_ _06785_/A vssd1 vssd1 vccd1 vccd1 _06785_/X sky130_fd_sc_hd__clkbuf_1
X_09573_ _09579_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09574_/A sky130_fd_sc_hd__and2_1
XFILLER_35_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _08524_/A vssd1 vssd1 vccd1 vccd1 _09140_/A sky130_fd_sc_hd__buf_2
XFILLER_35_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09530__A _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ _09330_/C _12252_/Q _09329_/B _09320_/D _08373_/X _08374_/X vssd1 vssd1 vccd1
+ vccd1 _08455_/X sky130_fd_sc_hd__mux4_2
XANTENNA__07969__B _07969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07406_ _07406_/A vssd1 vssd1 vccd1 vccd1 _08084_/A sky130_fd_sc_hd__buf_2
XFILLER_149_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08386_ _09322_/D _12245_/Q _12246_/Q _12247_/Q _08376_/X _08377_/X vssd1 vssd1 vccd1
+ vccd1 _08386_/X sky130_fd_sc_hd__mux4_2
XFILLER_136_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07337_ _07337_/A vssd1 vssd1 vccd1 vccd1 _07337_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07985__A _07999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ _07281_/A vssd1 vssd1 vccd1 vccd1 _07279_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09007_ _12841_/Q vssd1 vssd1 vccd1 vccd1 _11661_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07199_ _07199_/A vssd1 vssd1 vccd1 vccd1 _07199_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11300__A _11325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10924__C1 _10895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09909_ _13531_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09909_/X sky130_fd_sc_hd__or2_1
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12920_ _12923_/CLK _12920_/D vssd1 vssd1 vccd1 vccd1 _12920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _12853_/CLK _12851_/D vssd1 vssd1 vccd1 vccd1 _12851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08991__S1 _08913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11802_ _09623_/A _14002_/A _11805_/S vssd1 vssd1 vccd1 vccd1 _11803_/B sky130_fd_sc_hd__mux2_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12782_/CLK _12782_/D vssd1 vssd1 vccd1 vccd1 _13908_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _12860_/Q _14005_/A _11743_/S vssd1 vssd1 vccd1 vccd1 _11734_/B sky130_fd_sc_hd__mux2_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11677_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11667_/B sky130_fd_sc_hd__and2_1
X_13403_ _13403_/A _07963_/X vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__ebufn_8
X_10615_ _12568_/Q _13744_/A vssd1 vssd1 vccd1 vccd1 _10615_/Y sky130_fd_sc_hd__nor2_1
X_11595_ _11595_/A _11642_/A vssd1 vssd1 vccd1 vccd1 _11595_/X sky130_fd_sc_hd__and2_1
XFILLER_155_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10546_ _13692_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10546_/X sky130_fd_sc_hd__or2_1
XFILLER_6_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater131_A _14106_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10477_ _10477_/A _10477_/B vssd1 vssd1 vccd1 vccd1 _10478_/A sky130_fd_sc_hd__and2_1
XFILLER_136_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12216_ _12903_/CLK _12216_/D vssd1 vssd1 vccd1 vccd1 _13393_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12147_ _12147_/A vssd1 vssd1 vccd1 vccd1 _12965_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09615__A _09655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12078_ _11170_/X _12075_/X _12077_/X _12071_/X vssd1 vssd1 vccd1 vccd1 _12942_/D
+ sky130_fd_sc_hd__o211a_1
X_11029_ _11070_/B vssd1 vssd1 vccd1 vccd1 _11038_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06570_ _06570_/A vssd1 vssd1 vccd1 vccd1 _06570_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08240_ _08240_/A vssd1 vssd1 vccd1 vccd1 _08251_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08171_ _08228_/A vssd1 vssd1 vccd1 vccd1 _08184_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07122_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07122_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07053_ _07055_/A _07055_/B vssd1 vssd1 vccd1 vccd1 _07054_/A sky130_fd_sc_hd__or2_1
XFILLER_161_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11774__B _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ _07955_/A vssd1 vssd1 vccd1 vccd1 _07955_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__07971__C _07977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06906_ _06955_/A vssd1 vssd1 vccd1 vccd1 _06916_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_55_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07886_ _07894_/A _07890_/B _07890_/C vssd1 vssd1 vccd1 vccd1 _07887_/A sky130_fd_sc_hd__or3_1
XFILLER_56_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07045__A _07045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ _09625_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09625_/X sky130_fd_sc_hd__or2_1
XFILLER_83_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10685__A1 _10548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06837_ _06837_/A vssd1 vssd1 vccd1 vccd1 _06837_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11790__A _11790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _09563_/A _09556_/B vssd1 vssd1 vccd1 vccd1 _09557_/A sky130_fd_sc_hd__and2_1
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06768_ _07406_/A vssd1 vssd1 vccd1 vccd1 _06832_/A sky130_fd_sc_hd__clkbuf_2
X_08507_ _09362_/A _09368_/A _12268_/Q _12269_/Q _08417_/X _08418_/X vssd1 vssd1 vccd1
+ vccd1 _08507_/X sky130_fd_sc_hd__mux4_1
X_09487_ _13423_/A _09483_/X _09486_/X _09192_/X vssd1 vssd1 vccd1 vccd1 _12292_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06699_ _06701_/A _06706_/B _06706_/C vssd1 vssd1 vccd1 vccd1 _06700_/A sky130_fd_sc_hd__or3_1
X_08438_ _12237_/Q vssd1 vssd1 vccd1 vccd1 _09317_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11014__B _13947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08369_ _13393_/A vssd1 vssd1 vccd1 vccd1 _08525_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10400_ _13653_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10400_/X sky130_fd_sc_hd__or2_1
X_11380_ _11801_/A vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__buf_2
XFILLER_125_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10331_ _13657_/A _12511_/Q _10342_/S vssd1 vssd1 vccd1 vccd1 _10332_/B sky130_fd_sc_hd__mux2_1
XFILLER_118_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10262_ _13619_/A _10262_/B vssd1 vssd1 vccd1 vccd1 _10262_/X sky130_fd_sc_hd__or2_1
XFILLER_152_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ _12013_/A _12001_/B vssd1 vssd1 vccd1 vccd1 _12002_/A sky130_fd_sc_hd__and2_1
X_10193_ _10317_/A vssd1 vssd1 vccd1 vccd1 _10208_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13952_ _13952_/A _06417_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[17] sky130_fd_sc_hd__ebufn_8
XANTENNA__11322__C1 _11319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12903_ _12903_/CLK _12903_/D vssd1 vssd1 vccd1 vccd1 _13377_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__10676__A1 _10408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13883_ _13883_/A _06603_/X vssd1 vssd1 vccd1 vccd1 _13979_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12834_ _12842_/CLK _12834_/D vssd1 vssd1 vccd1 vccd1 _12834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13354__510 vssd1 vssd1 vccd1 vccd1 _13354__510/HI _14123_/A sky130_fd_sc_hd__conb_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12768_/CLK _12765_/D vssd1 vssd1 vccd1 vccd1 _12765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _12855_/Q _14000_/A _11726_/S vssd1 vssd1 vccd1 vccd1 _11717_/B sky130_fd_sc_hd__mux2_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12704_/CLK _12696_/D vssd1 vssd1 vccd1 vccd1 _12696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11647_ _11672_/A _11682_/B _11647_/C vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__and3b_1
Xinput13 peripheralBus_address[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput24 peripheralBus_address[9] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11578_ _11632_/D _11643_/B _11577_/Y vssd1 vssd1 vccd1 vccd1 _12823_/D sky130_fd_sc_hd__a21oi_1
XFILLER_116_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10529_ _13685_/A _10535_/B vssd1 vssd1 vccd1 vccd1 _10529_/X sky130_fd_sc_hd__or2_1
XFILLER_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07740_ _07740_/A vssd1 vssd1 vccd1 vccd1 _07740_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_74_clk_A _12555_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07671_ _07698_/A vssd1 vssd1 vccd1 vccd1 _07683_/B sky130_fd_sc_hd__clkbuf_1
X_09410_ _09410_/A vssd1 vssd1 vccd1 vccd1 _12276_/D sky130_fd_sc_hd__clkbuf_1
X_06622_ _06622_/A vssd1 vssd1 vccd1 vccd1 _06622_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13097__253 vssd1 vssd1 vccd1 vccd1 _13097__253/HI _13606_/A sky130_fd_sc_hd__conb_1
X_09341_ _09341_/A _09344_/B _09263_/X vssd1 vssd1 vccd1 vccd1 _12260_/D sky130_fd_sc_hd__nor3b_1
X_06553_ _06553_/A vssd1 vssd1 vccd1 vccd1 _06553_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_89_clk_A _12438_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07312__B _07317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ _09272_/A vssd1 vssd1 vccd1 vccd1 _12245_/D sky130_fd_sc_hd__clkbuf_1
X_06484_ _06494_/A _06486_/B _06486_/C vssd1 vssd1 vccd1 vccd1 _06485_/A sky130_fd_sc_hd__or3_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08223_ _08223_/A vssd1 vssd1 vccd1 vccd1 _08223_/X sky130_fd_sc_hd__clkbuf_1
X_13138__294 vssd1 vssd1 vccd1 vccd1 _13138__294/HI _13695_/A sky130_fd_sc_hd__conb_1
XANTENNA__10954__A _10971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A _12217_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11769__B _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ _08184_/A _08182_/B _08164_/C vssd1 vssd1 vccd1 vccd1 _08155_/A sky130_fd_sc_hd__or3_1
X_07105_ _07108_/A _07105_/B _07115_/C vssd1 vssd1 vccd1 vccd1 _07106_/A sky130_fd_sc_hd__or3_1
X_08085_ _08101_/A _08101_/B _08087_/C vssd1 vssd1 vccd1 vccd1 _08086_/A sky130_fd_sc_hd__or3_1
XFILLER_106_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07036_ _07036_/A vssd1 vssd1 vccd1 vccd1 _07036_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08987_ _11626_/C _11571_/D _12816_/Q _11627_/B _08911_/X _08913_/X vssd1 vssd1 vccd1
+ vccd1 _08987_/X sky130_fd_sc_hd__mux4_2
XFILLER_130_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_5_0_clk clkbuf_4_5_0_clk/A vssd1 vssd1 vccd1 vccd1 _12438_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_29_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07938_ _07999_/A vssd1 vssd1 vccd1 vccd1 _07951_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10658__A1 _10394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__B _13941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ _07869_/A vssd1 vssd1 vccd1 vccd1 _07869_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ _09608_/A _09608_/B _09608_/C vssd1 vssd1 vccd1 vccd1 _09608_/Y sky130_fd_sc_hd__nor3_1
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10880_ _10909_/A _10881_/A _10880_/C _10880_/D vssd1 vssd1 vccd1 vccd1 _10922_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09539_ _09546_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09540_/A sky130_fd_sc_hd__and2_1
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _12550_/CLK _12550_/D vssd1 vssd1 vccd1 vccd1 _13760_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11501_ _10939_/B _10939_/C _10939_/D _10938_/A _13973_/A _13974_/A vssd1 vssd1 vccd1
+ vccd1 _11501_/X sky130_fd_sc_hd__mux4_1
XFILLER_157_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ _12505_/CLK _12481_/D vssd1 vssd1 vccd1 vccd1 _12481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11432_ _13910_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11432_/X sky130_fd_sc_hd__or2_1
XFILLER_164_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11363_ _11363_/A vssd1 vssd1 vccd1 vccd1 _11377_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10314_ _13652_/A _12506_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10315_/B sky130_fd_sc_hd__mux2_1
X_14082_ _14082_/A _08045_/X vssd1 vssd1 vccd1 vccd1 _14082_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_106_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11294_ _10645_/X _11284_/X _11291_/X _11293_/X vssd1 vssd1 vccd1 vccd1 _12746_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10245_ _13762_/A _10244_/Y _10180_/S _09959_/X vssd1 vssd1 vccd1 vccd1 _12484_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09165__A _09631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ _10317_/A vssd1 vssd1 vccd1 vccd1 _10191_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13935_ _13935_/A _07846_/X vssd1 vssd1 vccd1 vccd1 _14063_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08711__A0 _08568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13866_ _13866_/A _06652_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
XFILLER_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07413__A _08168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12817_ _12829_/CLK _12817_/D vssd1 vssd1 vccd1 vccd1 _12817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13797_ _13797_/A _06844_/X vssd1 vssd1 vccd1 vccd1 _14117_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_97_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12782_/CLK _12748_/D vssd1 vssd1 vccd1 vccd1 _13875_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12679_ _12682_/CLK _12679_/D vssd1 vssd1 vccd1 vccd1 _13808_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10493__B _13757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08910_ _13968_/A vssd1 vssd1 vccd1 vccd1 _09067_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09890_ _13524_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09890_/X sky130_fd_sc_hd__or2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08772_/X _08774_/X _08773_/X _08840_/X _08876_/A _08838_/X vssd1 vssd1 vccd1
+ vccd1 _08841_/X sky130_fd_sc_hd__mux4_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10014__A _10160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07307__B _07317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ _12635_/Q _12636_/Q _12637_/Q _12638_/Q _08766_/X _08767_/X vssd1 vssd1 vccd1
+ vccd1 _08772_/X sky130_fd_sc_hd__mux4_2
XFILLER_111_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11837__A0 _14012_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07723_ _07723_/A vssd1 vssd1 vccd1 vccd1 _07723_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10949__A _10952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07654_ _07659_/A _07654_/B _07664_/C vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__or3_1
XFILLER_26_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06605_ _06633_/A vssd1 vssd1 vccd1 vccd1 _06616_/C sky130_fd_sc_hd__clkbuf_1
X_07585_ _07588_/A _07585_/B _07593_/C vssd1 vssd1 vccd1 vccd1 _07586_/A sky130_fd_sc_hd__or3_1
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08138__B _08189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _09347_/A _09336_/B _09336_/C vssd1 vssd1 vccd1 vccd1 _09324_/X sky130_fd_sc_hd__and3_1
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06536_ _06688_/A vssd1 vssd1 vccd1 vccd1 _06599_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09255_ _09316_/B _09256_/B _09248_/X vssd1 vssd1 vccd1 vccd1 _09257_/A sky130_fd_sc_hd__o21ai_1
XFILLER_21_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06467_ _06467_/A vssd1 vssd1 vccd1 vccd1 _06467_/X sky130_fd_sc_hd__clkbuf_1
X_08206_ _08212_/A _08208_/B _08212_/C vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__or3_1
XFILLER_154_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06398_ _06403_/A _06400_/B vssd1 vssd1 vccd1 vccd1 _06399_/A sky130_fd_sc_hd__or2_1
X_09186_ _11189_/A vssd1 vssd1 vccd1 vccd1 _09186_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__13995__A _13995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08137_ _08150_/A vssd1 vssd1 vccd1 vccd1 _08148_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07993__A _07997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ _08081_/A _08077_/B _08070_/C vssd1 vssd1 vccd1 vccd1 _08069_/A sky130_fd_sc_hd__or3_1
XFILLER_161_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07019_ _07019_/A _07019_/B vssd1 vssd1 vccd1 vccd1 _07020_/A sky130_fd_sc_hd__or2_1
XANTENNA__09194__A0 _11706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10030_ _10030_/A _10030_/B _10030_/C _10030_/D vssd1 vssd1 vccd1 vccd1 _10101_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__06402__A _07845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09041__S0 _08946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _13402_/A _12103_/B vssd1 vssd1 vccd1 vccd1 _12033_/S sky130_fd_sc_hd__nand2_4
XFILLER_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13720_ _13720_/A _07040_/X vssd1 vssd1 vccd1 vccd1 _13976_/Z sky130_fd_sc_hd__ebufn_8
X_10932_ _12659_/Q _10932_/B vssd1 vssd1 vccd1 vccd1 _10935_/B sky130_fd_sc_hd__and2_1
XANTENNA__07233__A _08177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13651_ _13651_/A _07225_/X vssd1 vssd1 vccd1 vccd1 _14099_/Z sky130_fd_sc_hd__ebufn_8
X_10863_ _10863_/A _10863_/B _10863_/C _10863_/D vssd1 vssd1 vccd1 vccd1 _10866_/B
+ sky130_fd_sc_hd__and4_1
X_12602_ _12652_/CLK _12602_/D vssd1 vssd1 vccd1 vccd1 _13777_/A sky130_fd_sc_hd__dfxtp_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13582_/A _07414_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
X_10794_ _10863_/B _10865_/A _10794_/C vssd1 vssd1 vccd1 vccd1 _10800_/B sky130_fd_sc_hd__and3_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _12533_/CLK _12533_/D vssd1 vssd1 vccd1 vccd1 _13662_/A sky130_fd_sc_hd__dfxtp_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12464_ _12467_/CLK _12464_/D vssd1 vssd1 vccd1 vccd1 _12464_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08064__A _08064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11415_ _11153_/X _11411_/X _11414_/X _11319_/X vssd1 vssd1 vccd1 vccd1 _12777_/D
+ sky130_fd_sc_hd__o211a_1
X_12395_ _12404_/CLK _12395_/D vssd1 vssd1 vccd1 vccd1 _13523_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_125_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11346_ _11363_/A vssd1 vssd1 vccd1 vccd1 _11361_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14065_ _14065_/A _07998_/X vssd1 vssd1 vccd1 vccd1 _14065_/Z sky130_fd_sc_hd__ebufn_8
X_11277_ _12731_/Q _13939_/A vssd1 vssd1 vccd1 vccd1 _11278_/D sky130_fd_sc_hd__xor2_1
XANTENNA__07408__A _07822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10228_ _12478_/Q _13753_/A vssd1 vssd1 vccd1 vccd1 _10232_/A sky130_fd_sc_hd__xor2_1
XFILLER_67_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06312__A _06462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10159_ _12467_/Q _10159_/B vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__xor2_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09623__A _09623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13918_ _13918_/A _06506_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
XFILLER_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10488__B _13756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13849_ _13849_/A _06700_/X vssd1 vssd1 vccd1 vccd1 _14009_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07370_ _07370_/A vssd1 vssd1 vccd1 vccd1 _07370_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06982__A _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06321_ _06321_/A vssd1 vssd1 vccd1 vccd1 _06321_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09040_ _08920_/X _08923_/X _08930_/X _08931_/X _08952_/X _08925_/X vssd1 vssd1 vccd1
+ vccd1 _09040_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09942_ _09160_/X _09921_/X _09941_/X _09916_/X vssd1 vssd1 vccd1 vccd1 _12412_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater93_A peripheralBus_data[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _11412_/B _09873_/B _10637_/B vssd1 vssd1 vccd1 vccd1 _09902_/A sky130_fd_sc_hd__or3_4
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _12648_/Q vssd1 vssd1 vccd1 vccd1 _10908_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11782__B _13367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08755_ _12640_/Q vssd1 vssd1 vccd1 vccd1 _10876_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _09484_/B vssd1 vssd1 vccd1 vccd1 _07763_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300__456 vssd1 vssd1 vccd1 vccd1 _13300__456/HI _14021_/A sky130_fd_sc_hd__conb_1
X_08686_ _08593_/X _08595_/X _08659_/X _08685_/X _08678_/X _08647_/X vssd1 vssd1 vccd1
+ vccd1 _08686_/X sky130_fd_sc_hd__mux4_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07637_ _09484_/B vssd1 vssd1 vccd1 vccd1 _07693_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07988__A _08022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ _07575_/A _08103_/B _07580_/C vssd1 vssd1 vccd1 vccd1 _07569_/A sky130_fd_sc_hd__or3_1
XANTENNA__06892__A _09125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09307_ _09330_/B _09306_/C _09330_/A vssd1 vssd1 vccd1 vccd1 _09308_/C sky130_fd_sc_hd__a21o_1
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06519_ _06521_/A _06526_/B _06526_/C vssd1 vssd1 vccd1 vccd1 _06520_/A sky130_fd_sc_hd__or3_1
X_07499_ _07553_/A vssd1 vssd1 vccd1 vccd1 _07510_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_09238_ _09242_/C _09238_/B vssd1 vssd1 vccd1 vccd1 _12237_/D sky130_fd_sc_hd__nor2_1
XFILLER_154_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ _09633_/A vssd1 vssd1 vccd1 vccd1 _10662_/A sky130_fd_sc_hd__buf_4
XFILLER_135_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _10552_/X _11185_/A _11199_/X _11195_/X vssd1 vssd1 vccd1 vccd1 _12726_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12180_ _14095_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__or2_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _12695_/Q _11388_/B vssd1 vssd1 vccd1 vccd1 _11131_/X sky130_fd_sc_hd__and2_1
XANTENNA__12134__A _12134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11062_ _13819_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11062_/X sky130_fd_sc_hd__or2_1
XFILLER_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10013_ _10021_/C _10016_/C vssd1 vssd1 vccd1 vccd1 _10014_/B sky130_fd_sc_hd__xor2_1
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input22_A peripheralBus_address[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11964_ _11998_/A vssd1 vssd1 vccd1 vccd1 _11978_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08059__A _08072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043__199 vssd1 vssd1 vccd1 vccd1 _13043__199/HI _13486_/A sky130_fd_sc_hd__conb_1
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13703_ _13703_/A _07085_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
X_10915_ _10915_/A _10921_/C _10915_/C vssd1 vssd1 vccd1 vccd1 _10915_/X sky130_fd_sc_hd__and3_1
XFILLER_72_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11895_ _12901_/Q _14045_/A _11895_/S vssd1 vssd1 vccd1 vccd1 _11896_/B sky130_fd_sc_hd__mux2_1
X_13634_ _13634_/A _07270_/X vssd1 vssd1 vccd1 vccd1 _13666_/Z sky130_fd_sc_hd__ebufn_8
X_10846_ _10875_/C _10848_/C _10781_/X vssd1 vssd1 vccd1 vccd1 _10847_/B sky130_fd_sc_hd__o21ai_1
XFILLER_158_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13565_ _13565_/A _07455_/X vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__ebufn_8
X_10777_ _10780_/B _10812_/B _10777_/C vssd1 vssd1 vccd1 vccd1 _10778_/A sky130_fd_sc_hd__and3b_1
XFILLER_9_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12516_ _12583_/CLK _12516_/D vssd1 vssd1 vccd1 vccd1 _12516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13496_ _13496_/A _07634_/X vssd1 vssd1 vccd1 vccd1 _14104_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_145_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12447_ _12451_/CLK _12447_/D vssd1 vssd1 vccd1 vccd1 _12447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09618__A _11160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12378_ _12386_/CLK _12378_/D vssd1 vssd1 vccd1 vccd1 _12378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _14117_/A _08256_/X vssd1 vssd1 vccd1 vccd1 _14117_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_125_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11329_ _11381_/S vssd1 vssd1 vccd1 vccd1 _11408_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14048_ _14048_/A _07909_/X vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_140_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06870_ _06877_/A _06870_/B _06870_/C vssd1 vssd1 vccd1 vccd1 _06871_/A sky130_fd_sc_hd__or3_1
XANTENNA__06977__A _07417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08540_ _11708_/C vssd1 vssd1 vccd1 vccd1 _13373_/A sky130_fd_sc_hd__buf_4
XFILLER_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08471_ _08388_/X _08389_/X _08390_/X _08469_/X _08479_/A _08470_/X vssd1 vssd1 vccd1
+ vccd1 _08471_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09881__A1 _09139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__B _10146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07422_ _07422_/A vssd1 vssd1 vccd1 vccd1 _07422_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07353_ _07393_/A vssd1 vssd1 vccd1 vccd1 _07364_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06304_ _06304_/A vssd1 vssd1 vccd1 vccd1 _06304_/X sky130_fd_sc_hd__clkbuf_1
X_07284_ _07292_/A _07289_/B _07286_/C vssd1 vssd1 vccd1 vccd1 _07285_/A sky130_fd_sc_hd__or3_1
X_09023_ _10938_/B vssd1 vssd1 vccd1 vccd1 _13940_/A sky130_fd_sc_hd__buf_6
XFILLER_148_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09528__A _09846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11777__B _13374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09925_ _09925_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _09963_/B sky130_fd_sc_hd__and2_1
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _12377_/Q _13554_/A vssd1 vssd1 vccd1 vccd1 _09858_/C sky130_fd_sc_hd__xor2_1
XANTENNA__10703__A0 _14098_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06887__A _07090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08807_ _08886_/A vssd1 vssd1 vccd1 vccd1 _08807_/X sky130_fd_sc_hd__buf_4
XFILLER_100_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09787_ _13501_/A _09787_/B vssd1 vssd1 vccd1 vccd1 _09787_/X sky130_fd_sc_hd__or2_1
XFILLER_85_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06999_ _07007_/A _07007_/B vssd1 vssd1 vccd1 vccd1 _07000_/A sky130_fd_sc_hd__or2_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _12620_/Q vssd1 vssd1 vccd1 vccd1 _10773_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11017__B _13940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _09396_/C vssd1 vssd1 vccd1 vccd1 _13557_/A sky130_fd_sc_hd__buf_6
XFILLER_14_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _10700_/A _10700_/B vssd1 vssd1 vccd1 vccd1 _10701_/A sky130_fd_sc_hd__or2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11680_/A _11687_/C _11680_/C vssd1 vssd1 vccd1 vccd1 _11680_/X sky130_fd_sc_hd__and3_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10856__B _10917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ _12567_/Q _13743_/A vssd1 vssd1 vccd1 vccd1 _10632_/D sky130_fd_sc_hd__xor2_1
XFILLER_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11431__A1 _10659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10562_ _10562_/A vssd1 vssd1 vccd1 vccd1 _12568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ _12301_/CLK _12301_/D vssd1 vssd1 vccd1 vccd1 _13432_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10872__A _10872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10493_ _12548_/Q _13757_/A vssd1 vssd1 vccd1 vccd1 _10494_/D sky130_fd_sc_hd__xor2_1
X_12232_ _12301_/CLK _12232_/D vssd1 vssd1 vccd1 vccd1 _12232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _12959_/Q _13365_/A vssd1 vssd1 vccd1 vccd1 _12166_/B sky130_fd_sc_hd__xor2_1
XFILLER_107_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11114_ _11206_/A vssd1 vssd1 vccd1 vccd1 _11204_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12094_ _14075_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12094_/X sky130_fd_sc_hd__or2_1
XFILLER_1_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11045_ _13813_/A _11051_/B vssd1 vssd1 vccd1 vccd1 _11045_/X sky130_fd_sc_hd__or2_1
XANTENNA__11498__A1 _13979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09173__A _09636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10112__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11947_ _11998_/A vssd1 vssd1 vccd1 vccd1 _11962_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11878_ _12896_/Q _14040_/A _11878_/S vssd1 vssd1 vccd1 vccd1 _11879_/B sky130_fd_sc_hd__mux2_1
X_13617_ _13617_/A _07315_/X vssd1 vssd1 vccd1 vccd1 _14033_/Z sky130_fd_sc_hd__ebufn_8
X_10829_ _12634_/Q vssd1 vssd1 vccd1 vccd1 _10870_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11422__A1 _10648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13548_ _13548_/A _07495_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_9_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13479_ _13479_/A _07677_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11597__B _11604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07971_ _07983_/A _07971_/B _07977_/C vssd1 vssd1 vccd1 vccd1 _07972_/A sky130_fd_sc_hd__or3_1
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09710_ _09710_/A vssd1 vssd1 vccd1 vccd1 _12355_/D sky130_fd_sc_hd__clkbuf_1
X_06922_ _06922_/A vssd1 vssd1 vccd1 vccd1 _06922_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09641_ _09655_/B vssd1 vssd1 vccd1 vccd1 _09653_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06853_ _06863_/A _06857_/B _06857_/C vssd1 vssd1 vccd1 vccd1 _06854_/A sky130_fd_sc_hd__or3_1
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09572_ _13467_/A _12320_/Q _09575_/S vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__mux2_1
X_06784_ _06788_/A _06793_/B _06793_/C vssd1 vssd1 vccd1 vccd1 _06785_/A sky130_fd_sc_hd__or3_1
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08523_ _12271_/Q vssd1 vssd1 vccd1 vccd1 _09382_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08454_ _12253_/Q vssd1 vssd1 vccd1 vccd1 _09329_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07405_ _07405_/A vssd1 vssd1 vccd1 vccd1 _07405_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08385_ _12244_/Q vssd1 vssd1 vccd1 vccd1 _09322_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07336_ _07342_/A _07336_/B _07347_/C vssd1 vssd1 vccd1 vccd1 _07337_/A sky130_fd_sc_hd__or3_1
XFILLER_149_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07267_ _07267_/A vssd1 vssd1 vccd1 vccd1 _07267_/X sky130_fd_sc_hd__clkbuf_1
X_09006_ _12840_/Q vssd1 vssd1 vccd1 vccd1 _11657_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07198_ _07206_/A _07203_/B _07200_/C vssd1 vssd1 vccd1 vccd1 _07199_/A sky130_fd_sc_hd__or3_1
XFILLER_105_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13265__421 vssd1 vssd1 vccd1 vccd1 _13265__421/HI _13956_/A sky130_fd_sc_hd__conb_1
XFILLER_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09908_ _09186_/X _09902_/X _09907_/X _09905_/X vssd1 vssd1 vccd1 vccd1 _12402_/D
+ sky130_fd_sc_hd__o211a_1
X_13306__462 vssd1 vssd1 vccd1 vccd1 _13306__462/HI _14027_/A sky130_fd_sc_hd__conb_1
XFILLER_86_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09839_ _09839_/A vssd1 vssd1 vccd1 vccd1 _12387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12850_ _12850_/CLK _12850_/D vssd1 vssd1 vccd1 vccd1 _12850_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _11801_/A vssd1 vssd1 vccd1 vccd1 _11816_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _12782_/CLK _12781_/D vssd1 vssd1 vccd1 vccd1 _13907_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11732_/A vssd1 vssd1 vccd1 vccd1 _12859_/D sky130_fd_sc_hd__clkbuf_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11677_/A _11664_/B _11576_/X vssd1 vssd1 vccd1 vccd1 _11665_/A sky130_fd_sc_hd__o21ai_1
XFILLER_14_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13402_ _13402_/A _07853_/X vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_8
X_10614_ _12568_/Q _10614_/B vssd1 vssd1 vccd1 vccd1 _10614_/X sky130_fd_sc_hd__and2_1
X_11594_ _11632_/A _11632_/B _11631_/C _11631_/D vssd1 vssd1 vccd1 vccd1 _11642_/A
+ sky130_fd_sc_hd__and4_1
X_10545_ _10285_/X _10538_/X _10544_/X _10536_/X vssd1 vssd1 vccd1 vccd1 _12563_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09168__A _14070_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08072__A _08072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10476_ _13693_/A _12548_/Q _10480_/S vssd1 vssd1 vccd1 vccd1 _10477_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12215_ _12295_/CLK _12215_/D vssd1 vssd1 vccd1 vccd1 _13392_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_142_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10107__A _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater124_A _14108_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12146_ _12149_/A _12146_/B vssd1 vssd1 vccd1 vccd1 _12147_/A sky130_fd_sc_hd__and2_1
XANTENNA__10391__A1 _09753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12077_ _14068_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12077_/X sky130_fd_sc_hd__or2_1
XFILLER_96_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output53_A _13378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ _11412_/A _11028_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _11070_/B sky130_fd_sc_hd__nor3_4
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12041__B _13362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09631__A _09631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12979_ _12980_/CLK _12979_/D vssd1 vssd1 vccd1 vccd1 _14104_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10496__B _13755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07151__A _07205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08170_ _09125_/B vssd1 vssd1 vccd1 vccd1 _08228_/A sky130_fd_sc_hd__buf_2
XFILLER_146_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07121_ _07121_/A _07131_/B _07128_/C vssd1 vssd1 vccd1 vccd1 _07122_/A sky130_fd_sc_hd__or3_1
XFILLER_118_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13249__405 vssd1 vssd1 vccd1 vccd1 _13249__405/HI _13920_/A sky130_fd_sc_hd__conb_1
X_07052_ _07052_/A vssd1 vssd1 vccd1 vccd1 _07052_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07954_ _07983_/A _07971_/B _07962_/C vssd1 vssd1 vccd1 vccd1 _07955_/A sky130_fd_sc_hd__or3_1
X_06905_ _10512_/B vssd1 vssd1 vccd1 vccd1 _06955_/A sky130_fd_sc_hd__buf_2
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07885_ _07885_/A vssd1 vssd1 vccd1 vccd1 _07885_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09624_ _13458_/A _09613_/X _09623_/X _09621_/X vssd1 vssd1 vccd1 vccd1 _12328_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06836_ _06836_/A _06843_/B _06843_/C vssd1 vssd1 vccd1 vccd1 _06837_/A sky130_fd_sc_hd__or3_1
X_09555_ _13462_/A _12315_/Q _09558_/S vssd1 vssd1 vccd1 vccd1 _09556_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11790__B _11924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06767_ _07603_/A vssd1 vssd1 vccd1 vccd1 _07406_/A sky130_fd_sc_hd__buf_4
XFILLER_71_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08506_ _08421_/X _08423_/X _08427_/X _08428_/X _08448_/X _08449_/X vssd1 vssd1 vccd1
+ vccd1 _08506_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09486_ _11153_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__or2_1
X_06698_ _06698_/A vssd1 vssd1 vccd1 vccd1 _06698_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ _09210_/A _09315_/D _12233_/Q _09316_/D _08417_/X _08418_/X vssd1 vssd1 vccd1
+ vccd1 _08437_/X sky130_fd_sc_hd__mux4_2
XFILLER_12_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08368_ _08524_/A vssd1 vssd1 vccd1 vccd1 _08368_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07319_ input7/X _11789_/C _07319_/C input5/X vssd1 vssd1 vccd1 vccd1 _09918_/B sky130_fd_sc_hd__or4b_4
XFILLER_127_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_112_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _12289_/CLK sky130_fd_sc_hd__clkbuf_16
X_08299_ _08364_/C vssd1 vssd1 vccd1 vccd1 _08309_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_109_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10330_ _10330_/A vssd1 vssd1 vccd1 vccd1 _12510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06405__A _07861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ _09753_/X _10249_/X _10260_/X _10256_/X vssd1 vssd1 vccd1 vccd1 _12488_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12000_ _12925_/Q _14068_/A _12012_/S vssd1 vssd1 vccd1 vccd1 _12001_/B sky130_fd_sc_hd__mux2_1
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10192_ _10192_/A vssd1 vssd1 vccd1 vccd1 _12474_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11570__B1 _11569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07236__A _11790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13951_ _13951_/A _06420_/X vssd1 vssd1 vccd1 vccd1 _13983_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11981__A _13402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ _12919_/CLK _12902_/D vssd1 vssd1 vccd1 vccd1 _12902_/Q sky130_fd_sc_hd__dfxtp_1
X_13882_ _13882_/A _06607_/X vssd1 vssd1 vccd1 vccd1 _13978_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_62_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12833_ _12835_/CLK _12833_/D vssd1 vssd1 vccd1 vccd1 _12833_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12768_/CLK _12764_/D vssd1 vssd1 vccd1 vccd1 _12764_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08067__A _08067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11715_ _11715_/A vssd1 vssd1 vccd1 vccd1 _12854_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12699_/CLK _12695_/D vssd1 vssd1 vccd1 vccd1 _12695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11646_ _11649_/B _11649_/C _11649_/D _11649_/A vssd1 vssd1 vccd1 vccd1 _11647_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 peripheralBus_address[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
Xinput25 peripheralBus_oe vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_4
X_11577_ _11632_/D _11643_/B _11576_/X vssd1 vssd1 vccd1 vccd1 _11577_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10528_ _10394_/X _10525_/X _10527_/X _10523_/X vssd1 vssd1 vccd1 vccd1 _12556_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12036__B _13368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10459_ _10480_/S vssd1 vssd1 vccd1 vccd1 _10473_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_97_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12129_ _12132_/A _12129_/B vssd1 vssd1 vccd1 vccd1 _12130_/A sky130_fd_sc_hd__and2_1
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07670_ _07670_/A vssd1 vssd1 vccd1 vccd1 _07670_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06985__A _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06621_ _06625_/A _06630_/B _06630_/C vssd1 vssd1 vccd1 vccd1 _06622_/A sky130_fd_sc_hd__or3_1
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09340_ _09370_/A _09346_/C _09363_/A vssd1 vssd1 vccd1 vccd1 _09344_/B sky130_fd_sc_hd__and3_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06552_ _06729_/A _07323_/B _06561_/C vssd1 vssd1 vccd1 vccd1 _06553_/A sky130_fd_sc_hd__or3_1
X_09271_ _09276_/C _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09272_/A sky130_fd_sc_hd__and3b_1
XFILLER_61_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06483_ _06523_/A vssd1 vssd1 vccd1 vccd1 _06494_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08222_ _08225_/A _08222_/B _08225_/C vssd1 vssd1 vccd1 vccd1 _08223_/A sky130_fd_sc_hd__or3_1
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08153_ _08153_/A vssd1 vssd1 vccd1 vccd1 _08164_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_119_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07104_ _07162_/A vssd1 vssd1 vccd1 vccd1 _07115_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08084_ _08084_/A vssd1 vssd1 vccd1 vccd1 _08101_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_134_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07035_ _07043_/A _07043_/B vssd1 vssd1 vccd1 vccd1 _07036_/A sky130_fd_sc_hd__or2_1
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08986_ _12817_/Q vssd1 vssd1 vccd1 vccd1 _11627_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07937_ _07937_/A vssd1 vssd1 vccd1 vccd1 _07937_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07868_ _07868_/A _07877_/B _07877_/C vssd1 vssd1 vccd1 vccd1 _07869_/A sky130_fd_sc_hd__or3_1
XFILLER_28_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09607_ _09607_/A _09607_/B _09607_/C _09607_/D vssd1 vssd1 vccd1 vccd1 _09608_/C
+ sky130_fd_sc_hd__or4_1
X_06819_ _06983_/B vssd1 vssd1 vccd1 vccd1 _07248_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07799_ _07809_/A _07806_/B _07801_/C vssd1 vssd1 vccd1 vccd1 _07800_/A sky130_fd_sc_hd__or3_1
X_09538_ _13457_/A _12310_/Q _09610_/B vssd1 vssd1 vccd1 vccd1 _09539_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09469_ _12275_/Q _13551_/A vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__xnor2_1
XFILLER_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11500_ _13980_/A _11459_/A _11499_/X _11497_/X vssd1 vssd1 vccd1 vccd1 _12806_/D
+ sky130_fd_sc_hd__o211a_1
X_12480_ _12522_/CLK _12480_/D vssd1 vssd1 vccd1 vccd1 _12480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _10659_/X _11425_/X _11429_/X _11430_/X vssd1 vssd1 vccd1 vccd1 _12783_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11041__A _11055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__B1 _09978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11362_ _11362_/A vssd1 vssd1 vccd1 vccd1 _12769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10313_ _10313_/A vssd1 vssd1 vccd1 vccd1 _12505_/D sky130_fd_sc_hd__clkbuf_1
X_14081_ _14081_/A _08043_/X vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ _11430_/A vssd1 vssd1 vccd1 vccd1 _11293_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10244_ _10244_/A _10244_/B vssd1 vssd1 vccd1 vccd1 _10244_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10175_ _10988_/A vssd1 vssd1 vccd1 vccd1 _10317_/A sky130_fd_sc_hd__clkbuf_2
X_12985__141 vssd1 vssd1 vccd1 vccd1 _12985__141/HI _13382_/A sky130_fd_sc_hd__conb_1
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13934_ _13934_/A _06461_/X vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09181__A _13625_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13865_ _13865_/A _06656_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[26] sky130_fd_sc_hd__ebufn_8
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09612__C _10637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11216__A _11254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12816_ _12820_/CLK _12816_/D vssd1 vssd1 vccd1 vccd1 _12816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13796_ _13796_/A _06849_/X vssd1 vssd1 vccd1 vccd1 _13988_/Z sky130_fd_sc_hd__ebufn_8
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12782_/CLK _12747_/D vssd1 vssd1 vccd1 vccd1 _13874_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _12682_/CLK _12678_/D vssd1 vssd1 vccd1 vccd1 _13807_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_147_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13170__326 vssd1 vssd1 vccd1 vccd1 _13170__326/HI _13763_/A sky130_fd_sc_hd__conb_1
XFILLER_147_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11629_ _11640_/B _11640_/C vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__and2_1
XFILLER_156_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08244__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13211__367 vssd1 vssd1 vccd1 vccd1 _13211__367/HI _13834_/A sky130_fd_sc_hd__conb_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _10908_/B _12648_/Q _12649_/Q _12650_/Q _08739_/X _08740_/X vssd1 vssd1 vccd1
+ vccd1 _08840_/X sky130_fd_sc_hd__mux4_2
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064__220 vssd1 vssd1 vccd1 vccd1 _13064__220/HI _13539_/A sky130_fd_sc_hd__conb_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _12631_/Q _12632_/Q _12633_/Q _12634_/Q _08766_/X _08767_/X vssd1 vssd1 vccd1
+ vccd1 _08771_/X sky130_fd_sc_hd__mux4_2
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07722_ _07727_/A _07724_/B _07732_/C vssd1 vssd1 vccd1 vccd1 _07723_/A sky130_fd_sc_hd__or3_1
XFILLER_27_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09091__A _14107_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07604__A _07923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13105__261 vssd1 vssd1 vccd1 vccd1 _13105__261/HI _13614_/A sky130_fd_sc_hd__conb_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07653_ _07653_/A vssd1 vssd1 vccd1 vccd1 _07653_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06604_ _06604_/A vssd1 vssd1 vccd1 vccd1 _06616_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_80_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07323__B _07323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07584_ _07584_/A vssd1 vssd1 vccd1 vccd1 _07584_/X sky130_fd_sc_hd__clkbuf_1
X_09323_ _09323_/A _09323_/B _09323_/C _09323_/D vssd1 vssd1 vccd1 vccd1 _09336_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_40_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06535_ _06535_/A vssd1 vssd1 vccd1 vccd1 _06535_/X sky130_fd_sc_hd__clkbuf_1
X_09254_ _09254_/A _09256_/B vssd1 vssd1 vccd1 vccd1 _12241_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08561__S0 _08559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06466_ _06729_/A _07827_/B _06472_/C vssd1 vssd1 vccd1 vccd1 _06467_/A sky130_fd_sc_hd__or3_1
XANTENNA__07977__C _07977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08205_ _08205_/A vssd1 vssd1 vccd1 vccd1 _08205_/X sky130_fd_sc_hd__clkbuf_1
X_09185_ _13626_/Z vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__buf_4
X_06397_ _06397_/A vssd1 vssd1 vccd1 vccd1 _06397_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08136_ _08136_/A vssd1 vssd1 vccd1 vccd1 _08136_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07993__B _08062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _08067_/A vssd1 vssd1 vccd1 vccd1 _08081_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07018_ _07018_/A vssd1 vssd1 vccd1 vccd1 _07018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08170__A _09125_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08969_ _12813_/Q _12814_/Q _11571_/D _12816_/Q _08967_/X _08968_/X vssd1 vssd1 vccd1
+ vccd1 _08969_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11980_ _11998_/A vssd1 vssd1 vccd1 vccd1 _11996_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09041__S1 _08947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ _12659_/Q _10932_/B _10757_/X vssd1 vssd1 vccd1 vccd1 _10933_/A sky130_fd_sc_hd__o21ai_1
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13650_ _13650_/A _07227_/X vssd1 vssd1 vccd1 vccd1 _14098_/Z sky130_fd_sc_hd__ebufn_8
X_10862_ _10874_/A vssd1 vssd1 vccd1 vccd1 _10862_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12802_/CLK _12601_/D vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__dfxtp_4
X_13581_ _13581_/A _07416_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10793_ _10793_/A vssd1 vssd1 vccd1 vccd1 _12625_/D sky130_fd_sc_hd__clkbuf_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08552__S0 _08549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12532_ _12583_/CLK _12532_/D vssd1 vssd1 vccd1 vccd1 _13661_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12463_ _12467_/CLK _12463_/D vssd1 vssd1 vccd1 vccd1 _12463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11414_ _13903_/A _11423_/B vssd1 vssd1 vccd1 vccd1 _11414_/X sky130_fd_sc_hd__or2_1
X_12394_ _12404_/CLK _12394_/D vssd1 vssd1 vccd1 vccd1 _13522_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_73_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11345_ _11345_/A vssd1 vssd1 vccd1 vccd1 _12764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14064_ _14064_/A _07996_/X vssd1 vssd1 vccd1 vccd1 _14064_/Z sky130_fd_sc_hd__ebufn_8
X_11276_ _12735_/Q _13943_/A vssd1 vssd1 vccd1 vccd1 _11278_/C sky130_fd_sc_hd__xor2_1
X_13048__204 vssd1 vssd1 vccd1 vccd1 _13048__204/HI _13507_/A sky130_fd_sc_hd__conb_1
XANTENNA__08080__A _11026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11516__B1 _11515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10227_ _10227_/A _10227_/B _10227_/C _10226_/Y vssd1 vssd1 vccd1 vccd1 _10244_/A
+ sky130_fd_sc_hd__or4b_1
XANTENNA_clkbuf_leaf_88_clk_A _12438_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07408__B _07840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10158_ _10158_/A vssd1 vssd1 vccd1 vccd1 _12466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10089_ _10089_/A _10089_/B _10089_/C vssd1 vssd1 vccd1 vccd1 _10094_/B sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_11_clk_A _12917_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08696__A0 _08628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13917_ _13917_/A _06508_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[14] sky130_fd_sc_hd__ebufn_8
X_13848_ _13848_/A _06702_/X vssd1 vssd1 vccd1 vccd1 _13976_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_26_clk_A _12881_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13779_ _13779_/A _06895_/X vssd1 vssd1 vccd1 vccd1 _14099_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__08543__S0 _09140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06320_ _06320_/A _06323_/B _06323_/C vssd1 vssd1 vccd1 vccd1 _06321_/A sky130_fd_sc_hd__or3_1
XFILLER_148_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_clk clkbuf_4_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09941_ _09941_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _09941_/X sky130_fd_sc_hd__or2_1
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09176__A1 _10665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _09872_/A vssd1 vssd1 vccd1 vccd1 _12390_/D sky130_fd_sc_hd__clkbuf_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater86_A _14033_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08823_ _12645_/Q vssd1 vssd1 vccd1 vccd1 _10909_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08754_ _12634_/Q _12635_/Q _10876_/D _12637_/Q _08742_/X _08743_/X vssd1 vssd1 vccd1
+ vccd1 _08754_/X sky130_fd_sc_hd__mux4_2
XFILLER_73_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _07705_/A vssd1 vssd1 vccd1 vccd1 _07705_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _10130_/B _12459_/Q _12460_/Q _12461_/Q _08549_/X _08551_/X vssd1 vssd1 vccd1
+ vccd1 _08685_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_92_clk _12438_/CLK vssd1 vssd1 vccd1 vccd1 _12418_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _07636_/A vssd1 vssd1 vccd1 vccd1 _07636_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07567_ _07623_/A vssd1 vssd1 vccd1 vccd1 _07580_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__10695__A _10872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09306_ _09330_/A _09330_/B _09306_/C vssd1 vssd1 vccd1 vccd1 _09312_/B sky130_fd_sc_hd__and3_1
XFILLER_110_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06518_ _06518_/A vssd1 vssd1 vccd1 vccd1 _06518_/X sky130_fd_sc_hd__clkbuf_1
X_07498_ _09875_/B vssd1 vssd1 vccd1 vccd1 _07553_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09237_ _09317_/C _09234_/A _09236_/X vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__o21ai_1
X_06449_ _06451_/A _06449_/B vssd1 vssd1 vccd1 vccd1 _06450_/A sky130_fd_sc_hd__or2_1
XFILLER_154_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09168_ _14070_/Z vssd1 vssd1 vccd1 vccd1 _09633_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_147_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08119_ _08119_/A vssd1 vssd1 vccd1 vccd1 _08119_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09099_ _09102_/A _12060_/A _12059_/B _12062_/B vssd1 vssd1 vccd1 vccd1 _12195_/A
+ sky130_fd_sc_hd__or4_2
X_11130_ _12695_/Q _13936_/A vssd1 vssd1 vccd1 vccd1 _11130_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09167__A1 _10659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11061_ _11061_/A vssd1 vssd1 vccd1 vccd1 _11061_/X sky130_fd_sc_hd__buf_6
XFILLER_135_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07228__B _07231_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10012_ _10012_/A vssd1 vssd1 vccd1 vccd1 _12431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A peripheralBus_address[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11963_ _11963_/A vssd1 vssd1 vccd1 vccd1 _12914_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_83_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _12659_/CLK sky130_fd_sc_hd__clkbuf_16
X_13702_ _13702_/A _07087_/X vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__ebufn_8
X_10914_ _10914_/A _10915_/C vssd1 vssd1 vccd1 vccd1 _12653_/D sky130_fd_sc_hd__nor2_1
X_11894_ _11894_/A vssd1 vssd1 vccd1 vccd1 _12900_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10101__C _10101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13633_ _13633_/A _07272_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
X_10845_ _10875_/C _10848_/C vssd1 vssd1 vccd1 vccd1 _10847_/A sky130_fd_sc_hd__and2_1
X_13564_ _13564_/A _07458_/X vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_8
X_10776_ _10865_/D _10785_/D vssd1 vssd1 vccd1 vccd1 _10777_/C sky130_fd_sc_hd__or2_1
XFILLER_157_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12515_ _12515_/CLK _12515_/D vssd1 vssd1 vccd1 vccd1 _12515_/Q sky130_fd_sc_hd__dfxtp_1
X_13495_ _13495_/A _07636_/X vssd1 vssd1 vccd1 vccd1 _13623_/Z sky130_fd_sc_hd__ebufn_8
X_12446_ _12451_/CLK _12446_/D vssd1 vssd1 vccd1 vccd1 _12446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12377_ _12377_/CLK _12377_/D vssd1 vssd1 vccd1 vccd1 _12377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11328_ _13977_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11381_/S sky130_fd_sc_hd__and2_4
XANTENNA__07419__A _07480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14116_ _14116_/A _08252_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[21] sky130_fd_sc_hd__ebufn_8
XFILLER_114_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12044__B _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282__438 vssd1 vssd1 vccd1 vccd1 _13282__438/HI _13987_/A sky130_fd_sc_hd__conb_1
XANTENNA__09158__A1 _10652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11259_ _12740_/Q _11386_/B vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__and2_1
X_14047_ _14047_/A _07904_/X vssd1 vssd1 vccd1 vccd1 _14111_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__09634__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10712__A1 _10394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13323__479 vssd1 vssd1 vccd1 vccd1 _13323__479/HI _14060_/A sky130_fd_sc_hd__conb_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07154__A _07533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_clk _12555_/CLK vssd1 vssd1 vccd1 vccd1 _12522_/CLK sky130_fd_sc_hd__clkbuf_16
X_08470_ _13395_/A vssd1 vssd1 vccd1 vccd1 _08470_/X sky130_fd_sc_hd__buf_2
XFILLER_63_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176__332 vssd1 vssd1 vccd1 vccd1 _13176__332/HI _13769_/A sky130_fd_sc_hd__conb_1
XFILLER_51_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07421_ _07430_/A _07423_/B vssd1 vssd1 vccd1 vccd1 _07422_/A sky130_fd_sc_hd__or2_1
XANTENNA__08516__S0 _08417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07352_ _07352_/A vssd1 vssd1 vccd1 vccd1 _07352_/X sky130_fd_sc_hd__clkbuf_1
X_06303_ _06303_/A _06308_/B _06308_/C vssd1 vssd1 vccd1 vccd1 _06304_/A sky130_fd_sc_hd__or3_1
X_13217__373 vssd1 vssd1 vccd1 vccd1 _13217__373/HI _13856_/A sky130_fd_sc_hd__conb_1
X_07283_ _07283_/A vssd1 vssd1 vccd1 vccd1 _07283_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09022_ _09019_/X _09021_/X _09043_/S vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__mux2_2
XFILLER_163_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09149__A1 _10645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09924_ _10107_/A vssd1 vssd1 vccd1 vccd1 _09982_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09544__A _09582_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _12380_/Q _13557_/A vssd1 vssd1 vccd1 vccd1 _09858_/B sky130_fd_sc_hd__xor2_1
XANTENNA_input7_A peripheralBus_address[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08806_ _12631_/Q vssd1 vssd1 vccd1 vccd1 _10874_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06998_ _07979_/B vssd1 vssd1 vccd1 vccd1 _07007_/B sky130_fd_sc_hd__clkbuf_1
X_09786_ _09112_/X _09776_/X _09785_/X _09781_/X vssd1 vssd1 vccd1 vccd1 _12371_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07064__A _08035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08737_ _12618_/Q vssd1 vssd1 vccd1 vccd1 _10773_/D sky130_fd_sc_hd__clkbuf_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _12634_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_clk_A clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07999__A _07999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _08664_/X _08667_/X _08682_/S vssd1 vssd1 vccd1 vccd1 _09396_/C sky130_fd_sc_hd__mux2_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07619_ _07630_/A _07626_/B _07621_/C vssd1 vssd1 vccd1 vccd1 _07620_/A sky130_fd_sc_hd__or3_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08599_ _09397_/B vssd1 vssd1 vccd1 vccd1 _09851_/B sky130_fd_sc_hd__buf_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08507__S0 _08417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ _12572_/Q _13748_/A vssd1 vssd1 vccd1 vccd1 _10632_/C sky130_fd_sc_hd__xor2_1
XFILLER_14_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10561_ _10567_/A _10561_/B vssd1 vssd1 vccd1 vccd1 _10562_/A sky130_fd_sc_hd__and2_1
XFILLER_155_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12300_ _12301_/CLK _12300_/D vssd1 vssd1 vccd1 vccd1 _13431_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10492_ _12537_/Q _13746_/A vssd1 vssd1 vccd1 vccd1 _10494_/C sky130_fd_sc_hd__xor2_1
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ _12301_/CLK _12231_/D vssd1 vssd1 vccd1 vccd1 _12231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12162_ _12956_/Q _13362_/A vssd1 vssd1 vccd1 vccd1 _12166_/A sky130_fd_sc_hd__xor2_1
X_11113_ _11113_/A vssd1 vssd1 vccd1 vccd1 _12705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13010__166 vssd1 vssd1 vccd1 vccd1 _13010__166/HI _13421_/A sky130_fd_sc_hd__conb_1
X_12093_ _11189_/X _12088_/X _12092_/X _12084_/X vssd1 vssd1 vccd1 vccd1 _12948_/D
+ sky130_fd_sc_hd__o211a_1
X_11044_ _10394_/X _11041_/X _11043_/X _11039_/X vssd1 vssd1 vccd1 vccd1 _12683_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _12850_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11946_ _11946_/A vssd1 vssd1 vccd1 vccd1 _12909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11877_ _11877_/A vssd1 vssd1 vccd1 vccd1 _12895_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11224__A _11363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13616_ _13616_/A _07318_/X vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_60_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10828_ _10828_/A _10828_/B vssd1 vssd1 vccd1 vccd1 _12633_/D sky130_fd_sc_hd__nor2_1
XFILLER_158_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12039__B _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13547_ _13547_/A _07497_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
X_10759_ _10863_/D _10774_/B _10758_/Y vssd1 vssd1 vccd1 vccd1 _12618_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__09629__A _11170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13478_ _13478_/A _07679_/X vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_161_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12429_ _12617_/CLK _12429_/D vssd1 vssd1 vccd1 vccd1 _12429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07149__A _11924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07970_ _07970_/A vssd1 vssd1 vccd1 vccd1 _07970_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09364__A _09379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ _06923_/A _06929_/B vssd1 vssd1 vccd1 vccd1 _06922_/A sky130_fd_sc_hd__or2_1
XFILLER_67_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09640_ _09640_/A vssd1 vssd1 vccd1 vccd1 _09640_/X sky130_fd_sc_hd__clkbuf_2
X_06852_ _06879_/A vssd1 vssd1 vccd1 vccd1 _06863_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__08985__S0 _08941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ _09571_/A vssd1 vssd1 vccd1 vccd1 _12319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06783_ _06809_/A vssd1 vssd1 vccd1 vccd1 _06793_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _12800_/CLK sky130_fd_sc_hd__clkbuf_16
X_08522_ _08381_/X _08386_/X _08388_/X _08389_/X _08448_/X _08517_/X vssd1 vssd1 vccd1
+ vccd1 _08522_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08453_ _12251_/Q vssd1 vssd1 vccd1 vccd1 _09330_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07404_ _07822_/A _07404_/B _07496_/C vssd1 vssd1 vccd1 vccd1 _07405_/A sky130_fd_sc_hd__or3_1
XANTENNA__07331__B _07336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08384_ _08371_/X _08375_/X _08378_/X _08381_/X _08382_/X _08383_/X vssd1 vssd1 vccd1
+ vccd1 _08384_/X sky130_fd_sc_hd__mux4_1
X_07335_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07347_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_136_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07266_ _07266_/A _07276_/B _07273_/C vssd1 vssd1 vccd1 vccd1 _07267_/A sky130_fd_sc_hd__or3_1
XFILLER_136_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09005_ _12839_/Q vssd1 vssd1 vccd1 vccd1 _11657_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_07197_ _07197_/A vssd1 vssd1 vccd1 vccd1 _07197_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__07059__A _08266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10924__A1 _10872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09790__A1 _09120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06898__A _07328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09907_ _13530_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09907_/X sky130_fd_sc_hd__or2_1
XFILLER_59_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09838_ _10173_/A _09838_/B vssd1 vssd1 vccd1 vccd1 _09839_/A sky130_fd_sc_hd__and2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06410__B _06412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11028__B _11028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09769_ _09767_/X _09759_/X _09768_/X _09765_/X vssd1 vssd1 vccd1 vccd1 _12365_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _12726_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _11800_/A vssd1 vssd1 vccd1 vccd1 _12873_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09721__B _13561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12780_/CLK _12780_/D vssd1 vssd1 vccd1 vccd1 _13906_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11740_/A _11731_/B vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__and2_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11662_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _12842_/D sky130_fd_sc_hd__nor2_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _13401_/A _07851_/X vssd1 vssd1 vccd1 vccd1 _14105_/Z sky130_fd_sc_hd__ebufn_8
X_10613_ _12578_/Q _10613_/B vssd1 vssd1 vccd1 vccd1 _10613_/X sky130_fd_sc_hd__and2_1
X_11593_ _11632_/B _11590_/A _11592_/Y vssd1 vssd1 vccd1 vccd1 _12827_/D sky130_fd_sc_hd__a21oi_1
XFILLER_155_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08900__S0 _10697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ _13691_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10544_/X sky130_fd_sc_hd__or2_1
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10475_ _10475_/A vssd1 vssd1 vccd1 vccd1 _12547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12214_ _12295_/CLK _12214_/D vssd1 vssd1 vccd1 vccd1 _13391_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_123_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12145_ _12965_/Q _14107_/A _12151_/S vssd1 vssd1 vccd1 vccd1 _12146_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater117_A _14079_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12076_ _12101_/B vssd1 vssd1 vccd1 vccd1 _12086_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_111_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11027_ _11055_/A vssd1 vssd1 vccd1 vccd1 _11027_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10123__A _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output46_A _13762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk _12759_/CLK vssd1 vssd1 vccd1 vccd1 _12753_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ _12980_/CLK _12978_/D vssd1 vssd1 vccd1 vccd1 _14103_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07432__A _07468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11929_ _11929_/A vssd1 vssd1 vccd1 vccd1 _11998_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07120_ _07120_/A vssd1 vssd1 vccd1 vccd1 _07131_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09359__A _09380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08263__A _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13288__444 vssd1 vssd1 vccd1 vccd1 _13288__444/HI _13993_/A sky130_fd_sc_hd__conb_1
X_07051_ _07055_/A _07055_/B vssd1 vssd1 vccd1 vccd1 _07052_/A sky130_fd_sc_hd__or2_1
XANTENNA__11401__B _13940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11159__A1 _11153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09772__A1 _09770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13329__485 vssd1 vssd1 vccd1 vccd1 _13329__485/HI _14082_/A sky130_fd_sc_hd__conb_1
XFILLER_102_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09094__A _11924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07953_ _07999_/A vssd1 vssd1 vccd1 vccd1 _07983_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06904_ _06913_/A vssd1 vssd1 vccd1 vccd1 _08168_/A sky130_fd_sc_hd__clkbuf_4
X_07884_ _07894_/A _07890_/B _07890_/C vssd1 vssd1 vccd1 vccd1 _07885_/A sky130_fd_sc_hd__or3_1
XFILLER_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09623_ _09623_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09623_/X sky130_fd_sc_hd__or2_1
XFILLER_83_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06835_ _06835_/A vssd1 vssd1 vccd1 vccd1 _06835_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09554_ _09554_/A vssd1 vssd1 vccd1 vccd1 _12314_/D sky130_fd_sc_hd__clkbuf_1
X_06766_ _06766_/A vssd1 vssd1 vccd1 vccd1 _06766_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08505_ _11707_/B vssd1 vssd1 vccd1 vccd1 _13368_/A sky130_fd_sc_hd__buf_4
X_09485_ _09526_/B vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__clkbuf_1
X_06697_ _06701_/A _06706_/B _06706_/C vssd1 vssd1 vccd1 vccd1 _06698_/A sky130_fd_sc_hd__or3_1
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08436_ _12234_/Q vssd1 vssd1 vccd1 vccd1 _09316_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_08367_ _13392_/A vssd1 vssd1 vccd1 vccd1 _08524_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07318_ _07318_/A vssd1 vssd1 vccd1 vccd1 _07318_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09269__A _09269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ _08298_/A vssd1 vssd1 vccd1 vccd1 _08298_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07249_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07260_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_137_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ _13618_/A _10262_/B vssd1 vssd1 vccd1 vccd1 _10260_/X sky130_fd_sc_hd__or2_1
XFILLER_152_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09716__B _13562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _10191_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10192_/A sky130_fd_sc_hd__and2_1
XFILLER_133_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11039__A _11039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13950_ _13950_/A _06422_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
XFILLER_47_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13081__237 vssd1 vssd1 vccd1 vccd1 _13081__237/HI _13576_/A sky130_fd_sc_hd__conb_1
XANTENNA__11322__A1 _11064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12901_ _12918_/CLK _12901_/D vssd1 vssd1 vccd1 vccd1 _12901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13881_ _13881_/A _06609_/X vssd1 vssd1 vccd1 vccd1 _14009_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _12835_/CLK _12832_/D vssd1 vssd1 vccd1 vccd1 _12832_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10074__B1_N _10160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13122__278 vssd1 vssd1 vccd1 vccd1 _13122__278/HI _13663_/A sky130_fd_sc_hd__conb_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07252__A _07291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_1_0_clk_A clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12776_/CLK _12763_/D vssd1 vssd1 vccd1 vccd1 _12763_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11723_/A _11714_/B vssd1 vssd1 vccd1 vccd1 _11715_/A sky130_fd_sc_hd__and2_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12699_/CLK _12694_/D vssd1 vssd1 vccd1 vccd1 _12694_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _11649_/A _11649_/B _11645_/C _11645_/D vssd1 vssd1 vccd1 vccd1 _11672_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput15 peripheralBus_address[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09451__A0 _13437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput26 peripheralBus_we vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__08083__A _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11576_ _11576_/A vssd1 vssd1 vccd1 vccd1 _11576_/X sky130_fd_sc_hd__buf_2
XFILLER_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10527_ _13684_/A _10535_/B vssd1 vssd1 vccd1 vccd1 _10527_/X sky130_fd_sc_hd__or2_1
X_13016__172 vssd1 vssd1 vccd1 vccd1 _13016__172/HI _13443_/A sky130_fd_sc_hd__conb_1
XFILLER_143_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10458_ _10458_/A vssd1 vssd1 vccd1 vccd1 _12542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10389_ _09750_/X _10379_/X _10388_/X _10383_/X vssd1 vssd1 vccd1 vccd1 _12520_/D
+ sky130_fd_sc_hd__o211a_1
X_12128_ _12960_/Q _14102_/A _12135_/S vssd1 vssd1 vccd1 vccd1 _12129_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12052__B _13367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ _12059_/A _12059_/B vssd1 vssd1 vccd1 vccd1 _12059_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09642__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06620_ _06633_/A vssd1 vssd1 vccd1 vccd1 _06630_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11077__A0 _13840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06551_ _08182_/B vssd1 vssd1 vccd1 vccd1 _06561_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09270_ _09347_/A _09328_/C _09334_/C _09328_/B vssd1 vssd1 vccd1 vccd1 _09271_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10824__B1 _10781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06482_ _06482_/A vssd1 vssd1 vccd1 vccd1 _06482_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08221_ _08221_/A vssd1 vssd1 vccd1 vccd1 _08221_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_159_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08152_ _08152_/A vssd1 vssd1 vccd1 vccd1 _08152_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_158_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07103_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07162_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11131__B _11388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08083_ _10693_/A vssd1 vssd1 vccd1 vccd1 _08101_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_clk _12917_/CLK vssd1 vssd1 vccd1 vccd1 _12961_/CLK sky130_fd_sc_hd__clkbuf_16
X_07034_ _10637_/A vssd1 vssd1 vccd1 vccd1 _07043_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_161_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08985_ _11518_/A _12811_/Q _12812_/Q _11626_/D _08941_/X _08942_/X vssd1 vssd1 vccd1
+ vccd1 _08985_/X sky130_fd_sc_hd__mux4_1
X_07936_ _07936_/A _07945_/B _07945_/C vssd1 vssd1 vccd1 vccd1 _07937_/A sky130_fd_sc_hd__or3_1
XFILLER_102_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11304__A1 _10659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07867_ _07920_/A vssd1 vssd1 vccd1 vccd1 _07877_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09606_ _12312_/Q _13555_/A vssd1 vssd1 vccd1 vccd1 _09607_/D sky130_fd_sc_hd__xor2_1
XFILLER_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06818_ _06818_/A vssd1 vssd1 vccd1 vccd1 _06818_/X sky130_fd_sc_hd__clkbuf_1
X_07798_ _07798_/A vssd1 vssd1 vccd1 vccd1 _07809_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08168__A _08168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09537_ _09537_/A vssd1 vssd1 vccd1 vccd1 _12309_/D sky130_fd_sc_hd__clkbuf_1
X_06749_ _06760_/A _06751_/B _06751_/C vssd1 vssd1 vccd1 vccd1 _06750_/A sky130_fd_sc_hd__or3_1
XFILLER_52_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10815__B1 _10803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09468_ _09468_/A _09468_/B _09468_/C _09468_/D vssd1 vssd1 vccd1 vccd1 _09479_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08419_ _09210_/B _09210_/A _12232_/Q _12233_/Q _08417_/X _08418_/X vssd1 vssd1 vccd1
+ vccd1 _08419_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09399_ _09399_/A _09399_/B _09399_/C _09399_/D vssd1 vssd1 vccd1 vccd1 _09400_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_11_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11430_ _11430_/A vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _11361_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11362_/A sky130_fd_sc_hd__and2_1
XFILLER_165_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10312_ _10315_/A _10312_/B vssd1 vssd1 vccd1 vccd1 _10313_/A sky130_fd_sc_hd__and2_1
XFILLER_152_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14080_ _14080_/A _08040_/X vssd1 vssd1 vccd1 vccd1 _14112_/Z sky130_fd_sc_hd__ebufn_8
X_11292_ _11443_/A vssd1 vssd1 vccd1 vccd1 _11430_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10243_ _10243_/A _10243_/B _10243_/C vssd1 vssd1 vccd1 vccd1 _10244_/B sky130_fd_sc_hd__or3_1
XFILLER_106_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10174_ _10174_/A vssd1 vssd1 vccd1 vccd1 _12469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13933_ _13933_/A _06465_/X vssd1 vssd1 vccd1 vccd1 _14125_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_86_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13864_ _13864_/A _06658_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[25] sky130_fd_sc_hd__ebufn_8
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12815_ _12829_/CLK _12815_/D vssd1 vssd1 vccd1 vccd1 _12815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13795_ _13795_/A _06851_/X vssd1 vssd1 vccd1 vccd1 _13987_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _12782_/CLK _12746_/D vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _12687_/CLK _12677_/D vssd1 vssd1 vccd1 vccd1 _13954_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11628_ _11628_/A _11628_/B _11628_/C _11628_/D vssd1 vssd1 vccd1 vccd1 _11645_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06326__A _07045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12047__B _13374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11559_ _11627_/A _11558_/C _11625_/B vssd1 vssd1 vccd1 vccd1 _11560_/C sky130_fd_sc_hd__a21o_1
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _08763_/X _08764_/X _08765_/X _08768_/X _08850_/A _08769_/X vssd1 vssd1 vccd1
+ vccd1 _08770_/X sky130_fd_sc_hd__mux4_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07721_ _07763_/A vssd1 vssd1 vccd1 vccd1 _07732_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07652_ _07659_/A _07654_/B _07664_/C vssd1 vssd1 vccd1 vccd1 _07653_/A sky130_fd_sc_hd__or3_1
XFILLER_38_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06603_ _06603_/A vssd1 vssd1 vccd1 vccd1 _06603_/X sky130_fd_sc_hd__clkbuf_1
X_07583_ _07588_/A _07585_/B _07593_/C vssd1 vssd1 vccd1 vccd1 _07584_/A sky130_fd_sc_hd__or3_1
XANTENNA__07323__C _08089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09322_ _09322_/A _09322_/B _09328_/B _09322_/D vssd1 vssd1 vccd1 vccd1 _09323_/D
+ sky130_fd_sc_hd__and4_1
X_06534_ _06534_/A _06540_/B _06540_/C vssd1 vssd1 vccd1 vccd1 _06535_/A sky130_fd_sc_hd__or3_1
XFILLER_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10273__A1 _09767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08561__S1 _08560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09253_ _09315_/A _09315_/B _09253_/C vssd1 vssd1 vccd1 vccd1 _09256_/B sky130_fd_sc_hd__and3_1
X_06465_ _06465_/A vssd1 vssd1 vccd1 vccd1 _06465_/X sky130_fd_sc_hd__clkbuf_1
X_08204_ _08212_/A _08208_/B _08212_/C vssd1 vssd1 vccd1 vccd1 _08205_/A sky130_fd_sc_hd__or3_1
X_09184_ _09182_/X _09130_/X _09183_/X _09141_/X vssd1 vssd1 vccd1 vccd1 _12224_/D
+ sky130_fd_sc_hd__o211a_1
X_06396_ _06403_/A _06400_/B vssd1 vssd1 vccd1 vccd1 _06397_/A sky130_fd_sc_hd__or2_1
XFILLER_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08135_ _08135_/A _08189_/B _08138_/C vssd1 vssd1 vccd1 vccd1 _08136_/A sky130_fd_sc_hd__or3_1
XFILLER_135_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08066_ _08066_/A vssd1 vssd1 vccd1 vccd1 _08066_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07993__C _07993_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ _07019_/A _07019_/B vssd1 vssd1 vccd1 vccd1 _07018_/A sky130_fd_sc_hd__or2_1
X_13344__500 vssd1 vssd1 vccd1 vccd1 _13344__500/HI _14113_/A sky130_fd_sc_hd__conb_1
XFILLER_162_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08968_ _09068_/A vssd1 vssd1 vccd1 vccd1 _08968_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07919_ _11154_/B vssd1 vssd1 vccd1 vccd1 _07931_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08899_ _12657_/Q vssd1 vssd1 vccd1 vccd1 _10928_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10930_ _12658_/Q _10927_/A _10929_/Y _10749_/X vssd1 vssd1 vccd1 vccd1 _12658_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10861_ _10861_/A vssd1 vssd1 vccd1 vccd1 _12642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12802_/CLK _12600_/D vssd1 vssd1 vccd1 vccd1 _13775_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_140_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13580_ _13580_/A _07418_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13193__349 vssd1 vssd1 vccd1 vccd1 _13193__349/HI _13800_/A sky130_fd_sc_hd__conb_1
X_10792_ _10795_/B _10812_/B _10792_/C vssd1 vssd1 vccd1 vccd1 _10793_/A sky130_fd_sc_hd__and3b_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08552__S1 _08551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12531_ _12583_/CLK _12531_/D vssd1 vssd1 vccd1 vccd1 _13660_/A sky130_fd_sc_hd__dfxtp_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11052__A _11443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12462_ _12467_/CLK _12462_/D vssd1 vssd1 vccd1 vccd1 _12462_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11213__A0 _13874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09957__A1 _09182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ _11452_/B vssd1 vssd1 vccd1 vccd1 _11423_/B sky130_fd_sc_hd__clkbuf_1
X_12393_ _12400_/CLK _12393_/D vssd1 vssd1 vccd1 vccd1 _13521_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11344_ _11344_/A _11344_/B vssd1 vssd1 vccd1 vccd1 _11345_/A sky130_fd_sc_hd__and2_1
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14063_ _14063_/A _08183_/X vssd1 vssd1 vccd1 vccd1 _14063_/Z sky130_fd_sc_hd__ebufn_8
X_11275_ _12727_/Q _13935_/A vssd1 vssd1 vccd1 vccd1 _11278_/B sky130_fd_sc_hd__xor2_1
X_13087__243 vssd1 vssd1 vccd1 vccd1 _13087__243/HI _13582_/A sky130_fd_sc_hd__conb_1
XFILLER_152_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10226_ _12469_/Q _13744_/A vssd1 vssd1 vccd1 vccd1 _10226_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_140_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07408__C _07496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10157_ _10159_/B _10157_/B _10157_/C vssd1 vssd1 vccd1 vccd1 _10158_/A sky130_fd_sc_hd__and3b_1
X_13128__284 vssd1 vssd1 vccd1 vccd1 _13128__284/HI _13669_/A sky130_fd_sc_hd__conb_1
XFILLER_94_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10088_ _10098_/C _10099_/C _10088_/C _10088_/D vssd1 vssd1 vccd1 vccd1 _10089_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13916_ _13916_/A _06511_/X vssd1 vssd1 vccd1 vccd1 _14012_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__09920__A _09937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13847_ _13847_/A _06705_/X vssd1 vssd1 vccd1 vccd1 _14007_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13778_ _13778_/A _06897_/X vssd1 vssd1 vccd1 vccd1 _14098_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12729_ _12776_/CLK _12729_/D vssd1 vssd1 vccd1 vccd1 _12729_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08543__S1 _09146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09940_ _09940_/A vssd1 vssd1 vccd1 vccd1 _12411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _11151_/A _09871_/B _09871_/C vssd1 vssd1 vccd1 vccd1 _09872_/A sky130_fd_sc_hd__and3_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08822_ _10876_/A _10875_/A _10874_/A _10881_/A _08807_/X _08808_/X vssd1 vssd1 vccd1
+ vccd1 _08822_/X sky130_fd_sc_hd__mux4_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07615__A _07615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater79_A _14034_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08753_ _12636_/Q vssd1 vssd1 vccd1 vccd1 _10876_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09333__C1 _09263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07704_ _07714_/A _07710_/B _07704_/C vssd1 vssd1 vccd1 vccd1 _07705_/A sky130_fd_sc_hd__or3_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08684_ _08580_/X _08582_/X _08588_/X _08591_/X _08678_/X _08647_/X vssd1 vssd1 vccd1
+ vccd1 _08684_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07635_ _07644_/A _07641_/B _07635_/C vssd1 vssd1 vccd1 vccd1 _07636_/A sky130_fd_sc_hd__or3_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07566_ _09484_/B vssd1 vssd1 vccd1 vccd1 _07623_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09305_ _09330_/B _09306_/C _09304_/Y vssd1 vssd1 vccd1 vccd1 _12254_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__07350__A _07403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06517_ _06521_/A _06526_/B _06526_/C vssd1 vssd1 vccd1 vccd1 _06518_/A sky130_fd_sc_hd__or3_1
X_07497_ _07497_/A vssd1 vssd1 vccd1 vccd1 _07497_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09236_ _09271_/C vssd1 vssd1 vccd1 vccd1 _09236_/X sky130_fd_sc_hd__clkbuf_4
X_06448_ _06448_/A vssd1 vssd1 vccd1 vccd1 _06448_/X sky130_fd_sc_hd__clkbuf_1
X_09167_ _10659_/A _09145_/X _09166_/X _09148_/X vssd1 vssd1 vccd1 vccd1 _12220_/D
+ sky130_fd_sc_hd__a211o_1
X_06379_ _07480_/A vssd1 vssd1 vccd1 vccd1 _08338_/A sky130_fd_sc_hd__clkbuf_4
X_08118_ _08122_/A _08128_/B _08122_/C vssd1 vssd1 vccd1 vccd1 _08119_/A sky130_fd_sc_hd__or3_1
XFILLER_162_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_0_0_clk_A clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09098_ _11789_/A _11789_/B _11789_/C _11789_/D vssd1 vssd1 vccd1 vccd1 _12062_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_119_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08049_ _11283_/B vssd1 vssd1 vccd1 vccd1 _08110_/B sky130_fd_sc_hd__buf_2
XFILLER_135_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11060_ _10414_/X _11055_/X _11059_/X _11053_/X vssd1 vssd1 vccd1 vccd1 _12689_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10011_ _10016_/C _10146_/A _10011_/C vssd1 vssd1 vccd1 vccd1 _10012_/A sky130_fd_sc_hd__and3b_1
XFILLER_76_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09724__B _13565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11962_ _11962_/A _11962_/B vssd1 vssd1 vccd1 vccd1 _11963_/A sky130_fd_sc_hd__and2_1
XFILLER_84_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09740__A _11283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ _13701_/A _07089_/X vssd1 vssd1 vccd1 vccd1 _14117_/Z sky130_fd_sc_hd__ebufn_8
X_10913_ _10922_/A _10922_/B _10922_/C vssd1 vssd1 vccd1 vccd1 _10915_/C sky130_fd_sc_hd__and3_1
XFILLER_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11893_ _11927_/A _11893_/B vssd1 vssd1 vccd1 vccd1 _11894_/A sky130_fd_sc_hd__and2_1
XFILLER_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13632_ _13632_/A _07274_/X vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ _12638_/Q vssd1 vssd1 vccd1 vccd1 _10875_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08356__A _08358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_11_0_clk_A clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13563_ _13563_/A _07460_/X vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__ebufn_8
X_10775_ _10803_/A vssd1 vssd1 vccd1 vccd1 _10812_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12514_ _12583_/CLK _12514_/D vssd1 vssd1 vccd1 vccd1 _12514_/Q sky130_fd_sc_hd__dfxtp_1
X_13494_ _13494_/A _07640_/X vssd1 vssd1 vccd1 vccd1 _14102_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_9_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12445_ _12451_/CLK _12445_/D vssd1 vssd1 vccd1 vccd1 _12445_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14093__A _14093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09187__A _13402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ _12377_/CLK _12376_/D vssd1 vssd1 vccd1 vccd1 _12376_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08091__A _08186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14115_ _14115_/A _08249_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[20] sky130_fd_sc_hd__ebufn_8
X_11327_ _11363_/A vssd1 vssd1 vccd1 vccd1 _11344_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14046_ _14046_/A _07902_/X vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__ebufn_8
X_11258_ _12740_/Q _13948_/A vssd1 vssd1 vccd1 vccd1 _11258_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13437__A _13437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ _10209_/A vssd1 vssd1 vccd1 vccd1 _12479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11189_ _11189_/A vssd1 vssd1 vccd1 vccd1 _11189_/X sky130_fd_sc_hd__buf_6
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12060__B _12062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07420_ _07468_/A vssd1 vssd1 vccd1 vccd1 _07430_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08266__A _08266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11404__B _13939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08516__S1 _08418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07351_ _07356_/A _07351_/B _07361_/C vssd1 vssd1 vccd1 vccd1 _07352_/A sky130_fd_sc_hd__or3_1
XFILLER_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06302_ _06302_/A vssd1 vssd1 vccd1 vccd1 _06302_/X sky130_fd_sc_hd__clkbuf_1
X_07282_ _07292_/A _07289_/B _07286_/C vssd1 vssd1 vccd1 vccd1 _07283_/A sky130_fd_sc_hd__or3_1
XFILLER_164_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09021_ _08957_/X _08960_/X _08959_/X _09020_/X _09057_/A _09013_/X vssd1 vssd1 vccd1
+ vccd1 _09021_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09923_ _10112_/A vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__buf_2
XFILLER_104_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _12384_/Q _13561_/A vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__xor2_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _12625_/Q _10863_/B _10863_/A _12628_/Q _08733_/X _08735_/X vssd1 vssd1 vccd1
+ vccd1 _08805_/X sky130_fd_sc_hd__mux4_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ _13500_/A _09787_/B vssd1 vssd1 vccd1 vccd1 _09785_/X sky130_fd_sc_hd__or2_1
X_06997_ _07033_/A vssd1 vssd1 vccd1 vccd1 _07007_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_39_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08736_ _12614_/Q _10806_/C _10806_/B _12617_/Q _08733_/X _08735_/X vssd1 vssd1 vccd1
+ vccd1 _08736_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08667_ _08615_/X _08619_/X _08617_/X _08666_/X _08663_/X _08652_/X vssd1 vssd1 vccd1
+ vccd1 _08667_/X sky130_fd_sc_hd__mux4_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07618_ _07661_/A vssd1 vssd1 vccd1 vccd1 _07630_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09609__B1 _13569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _08585_/X _08596_/X _08682_/S vssd1 vssd1 vccd1 vccd1 _09397_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08176__A _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08507__S1 _08418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _07558_/A _07558_/B _07551_/C vssd1 vssd1 vccd1 vccd1 _07550_/A sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_87_clk_A _12438_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06408__B _06412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10560_ _13712_/A _12568_/Q _10635_/B vssd1 vssd1 vccd1 vccd1 _10561_/B sky130_fd_sc_hd__mux2_1
X_09219_ _09224_/C _09219_/B vssd1 vssd1 vccd1 vccd1 _12232_/D sky130_fd_sc_hd__nor2_1
XFILLER_10_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09719__B _13564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ _12540_/Q _13749_/A vssd1 vssd1 vccd1 vccd1 _10494_/B sky130_fd_sc_hd__xor2_1
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10872__C _10881_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ _12301_/CLK _12230_/D vssd1 vssd1 vccd1 vccd1 _12230_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_10_clk_A _12217_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12161_ _12161_/A _12161_/B _12161_/C _12161_/D vssd1 vssd1 vccd1 vccd1 _12178_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_146_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11112_ _11112_/A _11112_/B vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__and2_1
X_12092_ _14074_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12092_/X sky130_fd_sc_hd__or2_1
XFILLER_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11043_ _13812_/A _11051_/B vssd1 vssd1 vccd1 vccd1 _11043_/X sky130_fd_sc_hd__or2_1
XFILLER_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08443__S0 _08368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_clk clkbuf_4_3_0_clk/A vssd1 vssd1 vccd1 vccd1 _12217_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_29_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13199__355 vssd1 vssd1 vccd1 vccd1 _13199__355/HI _13806_/A sky130_fd_sc_hd__conb_1
XFILLER_57_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11945_ _11945_/A _11945_/B vssd1 vssd1 vccd1 vccd1 _11946_/A sky130_fd_sc_hd__and2_1
XFILLER_55_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11876_ _11886_/A _11876_/B vssd1 vssd1 vccd1 vccd1 _11877_/A sky130_fd_sc_hd__and2_1
XANTENNA__11407__B1 _13951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13615_ _13615_/A _07994_/X vssd1 vssd1 vccd1 vccd1 _13775_/Z sky130_fd_sc_hd__ebufn_8
X_10827_ _10869_/C _10825_/A _10781_/X vssd1 vssd1 vccd1 vccd1 _10828_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13546_ _13546_/A _07501_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
X_10758_ _10863_/D _10774_/B _10757_/X vssd1 vssd1 vccd1 vccd1 _10758_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13477_ _13477_/A _07682_/X vssd1 vssd1 vccd1 vccd1 _13765_/Z sky130_fd_sc_hd__ebufn_8
X_10689_ _10706_/A vssd1 vssd1 vccd1 vccd1 _10703_/S sky130_fd_sc_hd__clkbuf_4
X_12428_ _12617_/CLK _12428_/D vssd1 vssd1 vccd1 vccd1 _12428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12359_ _12367_/CLK _12359_/D vssd1 vssd1 vccd1 vccd1 _13488_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14029_ _14029_/A _08192_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
X_06920_ _06920_/A vssd1 vssd1 vccd1 vccd1 _06920_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__12071__A _12084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07165__A _07205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06851_ _06851_/A vssd1 vssd1 vccd1 vccd1 _06851_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08985__S1 _08942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09570_ _09579_/A _09570_/B vssd1 vssd1 vccd1 vccd1 _09571_/A sky130_fd_sc_hd__and2_1
XFILLER_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06782_ _06832_/A vssd1 vssd1 vccd1 vccd1 _06793_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__09380__A _09380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08521_ _11707_/D vssd1 vssd1 vccd1 vccd1 _13370_/A sky130_fd_sc_hd__buf_4
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08452_ _09321_/C _12248_/Q _09322_/A _09321_/B _08445_/X _08446_/X vssd1 vssd1 vccd1
+ vccd1 _08452_/X sky130_fd_sc_hd__mux4_2
X_07403_ _07403_/A vssd1 vssd1 vccd1 vccd1 _07496_/C sky130_fd_sc_hd__buf_2
XFILLER_51_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11134__B _13945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ _13395_/A vssd1 vssd1 vccd1 vccd1 _08383_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07331__C _07739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07334_ _07334_/A vssd1 vssd1 vccd1 vccd1 _07334_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07265_ _07291_/A vssd1 vssd1 vccd1 vccd1 _07276_/B sky130_fd_sc_hd__clkbuf_1
X_09004_ _11641_/A _12835_/Q _11639_/A _12837_/Q _08946_/X _08947_/X vssd1 vssd1 vccd1
+ vccd1 _09004_/X sky130_fd_sc_hd__mux4_2
XFILLER_164_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07196_ _07206_/A _07203_/B _07200_/C vssd1 vssd1 vccd1 vccd1 _07197_/A sky130_fd_sc_hd__or3_1
XFILLER_129_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13033__189 vssd1 vssd1 vccd1 vccd1 _13033__189/HI _13476_/A sky130_fd_sc_hd__conb_1
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09790__A2 _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09906_ _09182_/X _09902_/X _09904_/X _09905_/X vssd1 vssd1 vccd1 vccd1 _12401_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07075__A _07090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ _13532_/A _12387_/Q _09837_/S vssd1 vssd1 vccd1 vccd1 _09838_/B sky130_fd_sc_hd__mux2_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08750__A0 _08736_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11028__C _11156_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ _13494_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09768_/X sky130_fd_sc_hd__or2_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _08612_/X _08615_/X _08614_/X _08617_/X _08663_/X _08670_/X vssd1 vssd1 vccd1
+ vccd1 _08719_/X sky130_fd_sc_hd__mux4_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09699_ _09705_/A _09699_/B vssd1 vssd1 vccd1 vccd1 _09700_/A sky130_fd_sc_hd__and2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _12859_/Q _14004_/A _11743_/S vssd1 vssd1 vccd1 vccd1 _11731_/B sky130_fd_sc_hd__mux2_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11677_/B _11661_/B _11661_/C vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__and3_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _13400_/A _07849_/X vssd1 vssd1 vccd1 vccd1 _14104_/Z sky130_fd_sc_hd__ebufn_8
X_10612_ _12578_/Q _13754_/A vssd1 vssd1 vccd1 vccd1 _10612_/Y sky130_fd_sc_hd__nor2_1
X_11592_ _11632_/B _11590_/A _11505_/B vssd1 vssd1 vccd1 vccd1 _11592_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10543_ _10414_/X _10538_/X _10542_/X _10536_/X vssd1 vssd1 vccd1 vccd1 _12562_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10474_ _10477_/A _10474_/B vssd1 vssd1 vccd1 vccd1 _10475_/A sky130_fd_sc_hd__and2_1
X_12213_ _12968_/CLK _12213_/D vssd1 vssd1 vccd1 vccd1 _14110_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12144_ _12144_/A vssd1 vssd1 vccd1 vccd1 _12964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12075_ _12088_/A vssd1 vssd1 vccd1 vccd1 _12075_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11026_ _11410_/A _11026_/B _11410_/C vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__or3_4
XFILLER_64_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07713__A _07892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output39_A _13594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12977_ _12980_/CLK _12977_/D vssd1 vssd1 vccd1 vccd1 _14102_/A sky130_fd_sc_hd__dfxtp_1
X_11928_ _11928_/A vssd1 vssd1 vccd1 vccd1 _12904_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11859_ _11869_/A _11859_/B vssd1 vssd1 vccd1 vccd1 _11860_/A sky130_fd_sc_hd__and2_1
XFILLER_33_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13529_ _13529_/A _07546_/X vssd1 vssd1 vccd1 vccd1 _13625_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07050_ _07050_/A vssd1 vssd1 vccd1 vccd1 _07050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11564__C1 _11515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07952_ _07952_/A vssd1 vssd1 vccd1 vccd1 _07952_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10119__B1 _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06903_ _06903_/A vssd1 vssd1 vccd1 vccd1 _06903_/X sky130_fd_sc_hd__clkbuf_1
X_07883_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07894_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09622_ _13457_/A _09613_/X _09620_/X _09621_/X vssd1 vssd1 vccd1 vccd1 _12327_/D
+ sky130_fd_sc_hd__o211a_1
X_06834_ _06836_/A _06843_/B _06843_/C vssd1 vssd1 vccd1 vccd1 _06835_/A sky130_fd_sc_hd__or3_1
XFILLER_56_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater61_A _14072_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09553_ _09563_/A _09553_/B vssd1 vssd1 vccd1 vccd1 _09554_/A sky130_fd_sc_hd__and2_1
X_06765_ _06775_/A _06765_/B _06765_/C vssd1 vssd1 vccd1 vccd1 _06766_/A sky130_fd_sc_hd__or3_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08504_ _08500_/X _08503_/X _08528_/S vssd1 vssd1 vccd1 vccd1 _11707_/B sky130_fd_sc_hd__mux2_1
X_09484_ _09484_/A _09484_/B _12062_/A vssd1 vssd1 vccd1 vccd1 _09526_/B sky130_fd_sc_hd__or3_2
X_06696_ _06722_/A vssd1 vssd1 vccd1 vccd1 _06706_/C sky130_fd_sc_hd__clkbuf_1
X_08435_ _12232_/Q vssd1 vssd1 vccd1 vccd1 _09315_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13360__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08366_ _12231_/Q vssd1 vssd1 vccd1 vccd1 _09210_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07317_ _07490_/A _07317_/B _07993_/C vssd1 vssd1 vccd1 vccd1 _07318_/A sky130_fd_sc_hd__or3_1
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08297_ _08300_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08298_/A sky130_fd_sc_hd__or2_1
XANTENNA__08894__S0 _10697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07248_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07302_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07179_ _07205_/A vssd1 vssd1 vccd1 vccd1 _07190_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09285__A _13391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ _13621_/A _12474_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__mux2_1
XFILLER_132_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12900_ _12919_/CLK _12900_/D vssd1 vssd1 vccd1 vccd1 _12900_/Q sky130_fd_sc_hd__dfxtp_1
X_13880_ _13880_/A _06611_/X vssd1 vssd1 vccd1 vccd1 _13976_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__09732__B _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07533__A _07533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12831_ _12835_/CLK _12831_/D vssd1 vssd1 vccd1 vccd1 _12831_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11055__A _11055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12776_/CLK _12762_/D vssd1 vssd1 vccd1 vccd1 _12762_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _12854_/Q _13999_/A _11726_/S vssd1 vssd1 vccd1 vccd1 _11714_/B sky130_fd_sc_hd__mux2_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12710_/CLK _12693_/D vssd1 vssd1 vccd1 vccd1 _13822_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11649_/B _11634_/X _11643_/Y _11515_/X vssd1 vssd1 vccd1 vccd1 _12837_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08364__A _08364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput16 peripheralBus_address[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
X_11575_ _11639_/C vssd1 vssd1 vccd1 vccd1 _11632_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput27 rst vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_6
X_10526_ _10553_/B vssd1 vssd1 vccd1 vccd1 _10535_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10457_ _10461_/A _10457_/B vssd1 vssd1 vccd1 vccd1 _10458_/A sky130_fd_sc_hd__and2_1
XFILLER_123_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10388_ _13649_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10388_/X sky130_fd_sc_hd__or2_1
XANTENNA__06612__A _06688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ _12127_/A vssd1 vssd1 vccd1 vccd1 _12959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09923__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ _13376_/A _12057_/Y _11711_/B _09404_/A _13402_/A vssd1 vssd1 vccd1 vccd1
+ _12936_/D sky130_fd_sc_hd__o2111a_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11009_ _12667_/Q _13941_/A vssd1 vssd1 vccd1 vccd1 _11011_/C sky130_fd_sc_hd__xor2_1
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06550_ _11285_/B vssd1 vssd1 vccd1 vccd1 _08182_/B sky130_fd_sc_hd__clkbuf_2
X_13255__411 vssd1 vssd1 vccd1 vccd1 _13255__411/HI _13926_/A sky130_fd_sc_hd__conb_1
XFILLER_61_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06481_ _06481_/A _06486_/B _06486_/C vssd1 vssd1 vccd1 vccd1 _06482_/A sky130_fd_sc_hd__or3_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08220_ _08225_/A _08222_/B _08225_/C vssd1 vssd1 vccd1 vccd1 _08221_/A sky130_fd_sc_hd__or3_1
XFILLER_60_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11412__B _11412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08151_ _08184_/A _08151_/B _08151_/C vssd1 vssd1 vccd1 vccd1 _08152_/A sky130_fd_sc_hd__or3_1
X_07102_ _07102_/A vssd1 vssd1 vccd1 vccd1 _07102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08082_ _08082_/A vssd1 vssd1 vccd1 vccd1 _08082_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07033_ _07033_/A vssd1 vssd1 vccd1 vccd1 _07043_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__08628__S0 _08549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08984_ _12813_/Q vssd1 vssd1 vccd1 vccd1 _11626_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07935_ _08004_/A vssd1 vssd1 vccd1 vccd1 _07945_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07866_ _08166_/A vssd1 vssd1 vccd1 vccd1 _07920_/A sky130_fd_sc_hd__clkbuf_4
X_09605_ _12316_/Q _13559_/A vssd1 vssd1 vccd1 vccd1 _09607_/C sky130_fd_sc_hd__xor2_1
XANTENNA__07353__A _07393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06817_ _07827_/A _07323_/B _07969_/B vssd1 vssd1 vccd1 vccd1 _06818_/A sky130_fd_sc_hd__or3_1
X_07797_ _07797_/A vssd1 vssd1 vccd1 vccd1 _07797_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09536_ _09546_/A _09536_/B vssd1 vssd1 vccd1 vccd1 _09537_/A sky130_fd_sc_hd__and2_1
XFILLER_71_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06748_ _06748_/A vssd1 vssd1 vccd1 vccd1 _06760_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09467_ _09467_/A _09467_/B _09467_/C _09467_/D vssd1 vssd1 vccd1 vccd1 _09468_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_52_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06679_ _06679_/A vssd1 vssd1 vccd1 vccd1 _06679_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08418_ _08525_/A vssd1 vssd1 vccd1 vccd1 _08418_/X sky130_fd_sc_hd__buf_2
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09398_ _09398_/A _09398_/B _09398_/C _09848_/B vssd1 vssd1 vccd1 vccd1 _09400_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039__195 vssd1 vssd1 vccd1 vccd1 _13039__195/HI _13482_/A sky130_fd_sc_hd__conb_1
X_08349_ _08349_/A _08349_/B vssd1 vssd1 vccd1 vccd1 _08350_/A sky130_fd_sc_hd__or2_1
XFILLER_165_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11360_ _13912_/A _12769_/Q _11373_/S vssd1 vssd1 vccd1 vccd1 _11361_/B sky130_fd_sc_hd__mux2_1
XFILLER_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10311_ _13651_/A _12505_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10312_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09727__B _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ _13873_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11291_/X sky130_fd_sc_hd__or2_1
XFILLER_152_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10242_ _10242_/A _10242_/B _10242_/C _10242_/D vssd1 vssd1 vccd1 vccd1 _10243_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10173_ _10173_/A _10173_/B vssd1 vssd1 vccd1 vccd1 _10174_/A sky130_fd_sc_hd__and2_1
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09743__A _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13932_ _13932_/A _06467_/X vssd1 vssd1 vccd1 vccd1 _14028_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13863_ _13863_/A _06660_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[24] sky130_fd_sc_hd__ebufn_8
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12814_ _12823_/CLK _12814_/D vssd1 vssd1 vccd1 vccd1 _12814_/Q sky130_fd_sc_hd__dfxtp_1
X_13794_ _13794_/A _06854_/X vssd1 vssd1 vccd1 vccd1 _14082_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _12782_/CLK _12745_/D vssd1 vssd1 vccd1 vccd1 _13872_/A sky130_fd_sc_hd__dfxtp_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12699_/CLK _12676_/D vssd1 vssd1 vccd1 vccd1 _12676_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11627_ _11627_/A _11627_/B _11627_/C _11627_/D vssd1 vssd1 vccd1 vccd1 _11628_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_128_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09918__A _11457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ _11625_/B _11627_/A _11558_/C vssd1 vssd1 vccd1 vccd1 _11565_/C sky130_fd_sc_hd__and3_1
XFILLER_144_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ _12062_/A vssd1 vssd1 vccd1 vccd1 _11410_/C sky130_fd_sc_hd__buf_2
XFILLER_128_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11489_ _13976_/Z _13976_/A _11489_/S vssd1 vssd1 vccd1 vccd1 _11490_/B sky130_fd_sc_hd__mux2_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09653__A _14109_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07720_ _07720_/A vssd1 vssd1 vccd1 vccd1 _07720_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11298__A1 _10652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09372__B _09372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07651_ _07693_/A vssd1 vssd1 vccd1 vccd1 _07664_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_93_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06602_ _06610_/A _06602_/B _06602_/C vssd1 vssd1 vccd1 vccd1 _06603_/A sky130_fd_sc_hd__or3_1
XFILLER_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07582_ _07623_/A vssd1 vssd1 vccd1 vccd1 _07593_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09321_ _09330_/C _09321_/B _09321_/C _09321_/D vssd1 vssd1 vccd1 vccd1 _09323_/C
+ sky130_fd_sc_hd__and4_1
X_06533_ _06533_/A vssd1 vssd1 vccd1 vccd1 _06533_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09252_ _09315_/A _09251_/B _09248_/X vssd1 vssd1 vccd1 vccd1 _09254_/A sky130_fd_sc_hd__o21ai_1
X_06464_ _06729_/A _07827_/B _06472_/C vssd1 vssd1 vccd1 vccd1 _06465_/A sky130_fd_sc_hd__or3_1
X_08203_ _08203_/A vssd1 vssd1 vccd1 vccd1 _08203_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11142__B _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09183_ _13401_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _09183_/X sky130_fd_sc_hd__or2_1
X_06395_ _06395_/A vssd1 vssd1 vccd1 vccd1 _06395_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08134_ _08134_/A vssd1 vssd1 vccd1 vccd1 _08134_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08732__A _13776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08065_ _08065_/A _08077_/B _08070_/C vssd1 vssd1 vccd1 vccd1 _08066_/A sky130_fd_sc_hd__or3_1
XFILLER_161_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07016_ _07016_/A vssd1 vssd1 vccd1 vccd1 _07016_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09026__S0 _08967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08967_ _09067_/A vssd1 vssd1 vccd1 vccd1 _08967_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07918_ _07918_/A vssd1 vssd1 vccd1 vccd1 _07918_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08898_ _08787_/X _08791_/X _08790_/X _08793_/X _08769_/X _08850_/X vssd1 vssd1 vccd1
+ vccd1 _08898_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09351__B1 _09248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07849_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07849_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _10936_/A _10860_/B _10860_/C vssd1 vssd1 vccd1 vccd1 _10861_/A sky130_fd_sc_hd__and3_1
XFILLER_140_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09519_ _11061_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09519_/X sky130_fd_sc_hd__or2_1
XFILLER_25_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07811__A _07923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09654__A1 _13469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ _10865_/A _10794_/C vssd1 vssd1 vccd1 vccd1 _10792_/C sky130_fd_sc_hd__or2_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12583_/CLK _12530_/D vssd1 vssd1 vccd1 vccd1 _13659_/A sky130_fd_sc_hd__dfxtp_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06427__A _06913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _12461_/CLK _12461_/D vssd1 vssd1 vccd1 vccd1 _12461_/Q sky130_fd_sc_hd__dfxtp_1
X_11412_ _11412_/A _11412_/B _11412_/C vssd1 vssd1 vccd1 vccd1 _11452_/B sky130_fd_sc_hd__nor3_2
XFILLER_138_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09738__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ _12400_/CLK _12392_/D vssd1 vssd1 vccd1 vccd1 _13520_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11343_ _13907_/A _12764_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _11344_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09457__B _13560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14062_ _14062_/A _07946_/X vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__ebufn_8
X_11274_ _12732_/Q _13940_/A vssd1 vssd1 vccd1 vccd1 _11278_/A sky130_fd_sc_hd__xor2_1
XFILLER_4_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10225_ _12477_/Q _13752_/A vssd1 vssd1 vccd1 vccd1 _10227_/C sky130_fd_sc_hd__xor2_1
XFILLER_133_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10156_ _10155_/B _10155_/C _12466_/Q vssd1 vssd1 vccd1 vccd1 _10157_/C sky130_fd_sc_hd__a21o_1
XFILLER_121_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11508__A _11634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ _10098_/A _10099_/A _10099_/B vssd1 vssd1 vccd1 vccd1 _10088_/D sky130_fd_sc_hd__and3_1
XANTENNA__08089__A _08089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13915_ _13915_/A _06513_/X vssd1 vssd1 vccd1 vccd1 _13979_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_74_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09893__A1 _09160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13846_ _13846_/A _06707_/X vssd1 vssd1 vccd1 vccd1 _14070_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13777_ _13777_/A _06899_/X vssd1 vssd1 vccd1 vccd1 _14097_/Z sky130_fd_sc_hd__ebufn_8
X_10989_ _11206_/A vssd1 vssd1 vccd1 vccd1 _11078_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12728_ _12743_/CLK _12728_/D vssd1 vssd1 vccd1 vccd1 _12728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ _12659_/CLK _12659_/D vssd1 vssd1 vccd1 vccd1 _12659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09648__A _10667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _09847_/Y _09853_/X _09869_/Y _13567_/A vssd1 vssd1 vccd1 vccd1 _09871_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _12644_/Q vssd1 vssd1 vccd1 vccd1 _10881_/A sky130_fd_sc_hd__clkbuf_2
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09008__S0 _08946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _10874_/C _12631_/Q _12632_/Q _12633_/Q _08742_/X _08743_/X vssd1 vssd1 vccd1
+ vccd1 _08752_/X sky130_fd_sc_hd__mux4_2
XFILLER_100_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07703_ _07703_/A vssd1 vssd1 vccd1 vccd1 _07703_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11137__B _13938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08683_ _09398_/A vssd1 vssd1 vccd1 vccd1 _13559_/A sky130_fd_sc_hd__buf_6
XFILLER_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07634_ _07634_/A vssd1 vssd1 vccd1 vccd1 _07634_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07565_ _07565_/A vssd1 vssd1 vccd1 vccd1 _07565_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09304_ _09330_/B _09306_/C _09392_/A vssd1 vssd1 vccd1 vccd1 _09304_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11153__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06516_ _07507_/A vssd1 vssd1 vccd1 vccd1 _06526_/C sky130_fd_sc_hd__clkbuf_1
X_07496_ _07504_/A _07504_/B _07496_/C vssd1 vssd1 vccd1 vccd1 _07497_/A sky130_fd_sc_hd__or3_1
XFILLER_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09235_ _09317_/C _09317_/D _09235_/C vssd1 vssd1 vccd1 vccd1 _09242_/C sky130_fd_sc_hd__and3_1
XFILLER_139_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06447_ _06451_/A _06449_/B vssd1 vssd1 vccd1 vccd1 _06448_/A sky130_fd_sc_hd__or2_1
XFILLER_22_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09166_ _13397_/A _09179_/B vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__and2_1
X_06378_ _06548_/C _07603_/A _06725_/A vssd1 vssd1 vccd1 vccd1 _07480_/A sky130_fd_sc_hd__or3_4
XFILLER_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08117_ _08117_/A vssd1 vssd1 vccd1 vccd1 _08117_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09097_ _09097_/A _09097_/B _09097_/C vssd1 vssd1 vccd1 vccd1 _11789_/D sky130_fd_sc_hd__or3_1
XFILLER_119_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08048_ _08048_/A vssd1 vssd1 vccd1 vccd1 _08048_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10010_ _10021_/D _10022_/A vssd1 vssd1 vccd1 vccd1 _10011_/C sky130_fd_sc_hd__or2_1
XFILLER_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09999_ _09997_/A _09996_/A _09994_/X vssd1 vssd1 vccd1 vccd1 _10000_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11328__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13160__316 vssd1 vssd1 vccd1 vccd1 _13160__316/HI _13733_/A sky130_fd_sc_hd__conb_1
XFILLER_28_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ peripheralBus_data[10] _14041_/A _11974_/S vssd1 vssd1 vccd1 vccd1 _11962_/B
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10912_ _10922_/A _10909_/X _10757_/X vssd1 vssd1 vccd1 vccd1 _10914_/A sky130_fd_sc_hd__o21ai_1
X_13700_ _13700_/A _07092_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13201__357 vssd1 vssd1 vccd1 vccd1 _13201__357/HI _13824_/A sky130_fd_sc_hd__conb_1
X_11892_ _12900_/Q _14044_/A _11895_/S vssd1 vssd1 vccd1 vccd1 _11893_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13631_ _13631_/A _07277_/X vssd1 vssd1 vccd1 vccd1 _14079_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10843_ _10843_/A vssd1 vssd1 vccd1 vccd1 _12637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08356__B _08358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13562_ _13562_/A _07463_/X vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_13_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10774_ _10865_/D _10774_/B _10809_/B vssd1 vssd1 vccd1 vccd1 _10780_/B sky130_fd_sc_hd__and3_1
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08075__C _08110_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ _12583_/CLK _12513_/D vssd1 vssd1 vccd1 vccd1 _12513_/Q sky130_fd_sc_hd__dfxtp_1
X_13054__210 vssd1 vssd1 vccd1 vccd1 _13054__210/HI _13513_/A sky130_fd_sc_hd__conb_1
XANTENNA__11998__A _11998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13493_ _13493_/A _07642_/X vssd1 vssd1 vccd1 vccd1 _14037_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_157_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12444_ _12451_/CLK _12444_/D vssd1 vssd1 vccd1 vccd1 _12444_/Q sky130_fd_sc_hd__dfxtp_1
X_12375_ _12377_/CLK _12375_/D vssd1 vssd1 vccd1 vccd1 _12375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14114_ _14114_/A _08247_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[19] sky130_fd_sc_hd__ebufn_8
XFILLER_99_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11326_ _10552_/X _11312_/A _11325_/X _11319_/X vssd1 vssd1 vccd1 vccd1 _12759_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14045_ _14045_/A _07900_/X vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__ebufn_8
X_11257_ _12736_/Q _13944_/A vssd1 vssd1 vccd1 vccd1 _11257_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_69_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09915__B _09915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10208_ _10208_/A _10208_/B vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__and2_1
X_11188_ _11184_/X _11185_/X _11187_/X _11180_/X vssd1 vssd1 vccd1 vccd1 _12721_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10139_ _10142_/B _10157_/B _10139_/C vssd1 vssd1 vccd1 vccd1 _10140_/A sky130_fd_sc_hd__and3b_1
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11673__A1 _11689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13829_ _13829_/A _06752_/X vssd1 vssd1 vccd1 vccd1 _14117_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07350_ _07403_/A vssd1 vssd1 vccd1 vccd1 _07361_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06301_ _06303_/A _06308_/B _06308_/C vssd1 vssd1 vccd1 vccd1 _06302_/A sky130_fd_sc_hd__or3_1
X_07281_ _07281_/A vssd1 vssd1 vccd1 vccd1 _07292_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_148_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ _11657_/B _12841_/Q _12842_/Q _12843_/Q _08918_/X _08919_/X vssd1 vssd1 vccd1
+ vccd1 _09020_/X sky130_fd_sc_hd__mux4_2
XFILLER_164_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09097__B _09097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09922_ _13583_/A vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater91_A peripheralBus_data[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09853_ _09848_/X _09849_/Y _09850_/Y _09851_/X _09852_/Y vssd1 vssd1 vccd1 vccd1
+ _09853_/X sky130_fd_sc_hd__o221a_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _12627_/Q vssd1 vssd1 vccd1 vccd1 _10863_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09784_ _09092_/X _09776_/X _09783_/X _09781_/X vssd1 vssd1 vccd1 vccd1 _12370_/D
+ sky130_fd_sc_hd__o211a_1
X_06996_ _06996_/A vssd1 vssd1 vccd1 vccd1 _06996_/X sky130_fd_sc_hd__clkbuf_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09841__A _10173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ _08887_/A vssd1 vssd1 vccd1 vccd1 _08735_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13363__A _13363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _10111_/A _10130_/D _12457_/Q _12458_/Q _08575_/X _08576_/X vssd1 vssd1 vccd1
+ vccd1 _08666_/X sky130_fd_sc_hd__mux4_2
XFILLER_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _07617_/A vssd1 vssd1 vccd1 vccd1 _07617_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08597_ _13588_/A vssd1 vssd1 vccd1 vccd1 _08682_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_42_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07548_ _08197_/A vssd1 vssd1 vccd1 vccd1 _07558_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_14_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07479_ _07479_/A vssd1 vssd1 vccd1 vccd1 _07479_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09218_ _09315_/D _09211_/X _09217_/X vssd1 vssd1 vccd1 vccd1 _09219_/B sky130_fd_sc_hd__o21ai_1
X_10490_ _12544_/Q _13753_/A vssd1 vssd1 vccd1 vccd1 _10494_/A sky130_fd_sc_hd__xor2_1
XFILLER_148_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09149_ _10645_/A _09145_/X _09146_/X _09148_/X vssd1 vssd1 vccd1 vccd1 _12216_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _12954_/Q _13360_/A vssd1 vssd1 vccd1 vccd1 _12161_/D sky130_fd_sc_hd__xor2_1
XFILLER_123_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11111_ _13850_/A _12705_/Q _11118_/S vssd1 vssd1 vccd1 vccd1 _11112_/B sky130_fd_sc_hd__mux2_1
XFILLER_162_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12091_ _11184_/X _12088_/X _12090_/X _12084_/X vssd1 vssd1 vccd1 vccd1 _12947_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11042_ _11070_/B vssd1 vssd1 vccd1 vccd1 _11051_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08443__S1 _08370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input20_A peripheralBus_address[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09470__B _13564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ peripheralBus_data[5] _14036_/A _11957_/S vssd1 vssd1 vccd1 vccd1 _11945_/B
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11505__B _11505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11875_ _12895_/Q _14039_/A _11878_/S vssd1 vssd1 vccd1 vccd1 _11876_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10826_ _10869_/C _10869_/D _10840_/C vssd1 vssd1 vccd1 vccd1 _10828_/A sky130_fd_sc_hd__and3_1
X_13614_ _13614_/A _07324_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13545_ _13545_/A _07503_/X vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_8
X_10757_ _10803_/A vssd1 vssd1 vccd1 vccd1 _10757_/X sky130_fd_sc_hd__buf_2
XANTENNA__12080__A1 _10659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11521__A _11582_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13476_ _13476_/A _07684_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
X_10688_ _11457_/A _11924_/B _10688_/C vssd1 vssd1 vccd1 vccd1 _10706_/A sky130_fd_sc_hd__or3_4
XFILLER_139_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12427_ _12659_/CLK _12427_/D vssd1 vssd1 vccd1 vccd1 _12427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12358_ _12369_/CLK _12358_/D vssd1 vssd1 vccd1 vccd1 _13487_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09926__A _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11309_ _10665_/X _11299_/X _11308_/X _11306_/X vssd1 vssd1 vccd1 vccd1 _12752_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12289_ _12289_/CLK _12289_/D vssd1 vssd1 vccd1 vccd1 _12289_/Q sky130_fd_sc_hd__dfxtp_1
X_14028_ _14028_/A _08196_/X vssd1 vssd1 vccd1 vccd1 _14028_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06850_ _06850_/A _06857_/B _06857_/C vssd1 vssd1 vccd1 vccd1 _06851_/A sky130_fd_sc_hd__or3_1
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06781_ _06781_/A vssd1 vssd1 vccd1 vccd1 _06781_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08520_ _08513_/X _08518_/X _09162_/A vssd1 vssd1 vccd1 vccd1 _11707_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08451_ _12247_/Q vssd1 vssd1 vccd1 vccd1 _09321_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07402_ _07402_/A vssd1 vssd1 vccd1 vccd1 _07402_/X sky130_fd_sc_hd__clkbuf_1
X_08382_ _13394_/A vssd1 vssd1 vccd1 vccd1 _08382_/X sky130_fd_sc_hd__buf_2
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07333_ _07342_/A _07336_/B _07739_/C vssd1 vssd1 vccd1 vccd1 _07334_/A sky130_fd_sc_hd__or3_1
XFILLER_149_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07264_ _07264_/A vssd1 vssd1 vccd1 vccd1 _07264_/X sky130_fd_sc_hd__clkbuf_1
X_09003_ _12834_/Q vssd1 vssd1 vccd1 vccd1 _11641_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07195_ _07208_/A vssd1 vssd1 vccd1 vccd1 _07206_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_117_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09836__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09905_ _10256_/A vssd1 vssd1 vccd1 vccd1 _09905_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _09836_/A vssd1 vssd1 vccd1 vccd1 _10173_/A sky130_fd_sc_hd__buf_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09767_ _10662_/A vssd1 vssd1 vccd1 vccd1 _09767_/X sky130_fd_sc_hd__buf_6
XFILLER_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06979_ _07417_/A _07969_/B vssd1 vssd1 vccd1 vccd1 _06980_/A sky130_fd_sc_hd__or2_1
XFILLER_74_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _09399_/B vssd1 vssd1 vccd1 vccd1 _13564_/A sky130_fd_sc_hd__buf_4
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _13498_/A _12352_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09699_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10510__A _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08187__A _08240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11325__B _11325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ _13588_/A vssd1 vssd1 vccd1 vccd1 _08712_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13272__428 vssd1 vssd1 vccd1 vccd1 _13272__428/HI _13963_/A sky130_fd_sc_hd__conb_1
X_11660_ _11677_/B _11659_/B _11576_/X vssd1 vssd1 vccd1 vccd1 _11662_/A sky130_fd_sc_hd__o21ai_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10611_ _12576_/Q _13752_/A vssd1 vssd1 vccd1 vccd1 _10611_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_41_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_115_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _12242_/CLK sky130_fd_sc_hd__clkbuf_16
X_11591_ _12827_/Q vssd1 vssd1 vccd1 vccd1 _11632_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10542_ _13690_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__or2_1
XFILLER_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13313__469 vssd1 vssd1 vccd1 vccd1 _13313__469/HI _14050_/A sky130_fd_sc_hd__conb_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10473_ _13692_/A _12547_/Q _10473_/S vssd1 vssd1 vccd1 vccd1 _10474_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12212_ _12968_/CLK _12212_/D vssd1 vssd1 vccd1 vccd1 _14109_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12143_ _12149_/A _12143_/B vssd1 vssd1 vccd1 vccd1 _12144_/A sky130_fd_sc_hd__and2_1
X_13166__322 vssd1 vssd1 vccd1 vccd1 _13166__322/HI _13739_/A sky130_fd_sc_hd__conb_1
XANTENNA__09465__B _13554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12074_ _10652_/A _12061_/X _12073_/X _12071_/X vssd1 vssd1 vccd1 vccd1 _12941_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11025_ _13954_/A _11023_/Y _10955_/S _11024_/X vssd1 vssd1 vccd1 vccd1 _12677_/D
+ sky130_fd_sc_hd__o211a_1
X_13207__363 vssd1 vssd1 vccd1 vccd1 _13207__363/HI _13830_/A sky130_fd_sc_hd__conb_1
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12976_ _12980_/CLK _12976_/D vssd1 vssd1 vccd1 vccd1 _14101_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11927_ _11927_/A _11927_/B vssd1 vssd1 vccd1 vccd1 _11928_/A sky130_fd_sc_hd__and2_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11858_ _12890_/Q _14034_/A _11861_/S vssd1 vssd1 vccd1 vccd1 _11859_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_106_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _12331_/CLK sky130_fd_sc_hd__clkbuf_16
X_10809_ _10866_/A _10809_/B _10809_/C _10809_/D vssd1 vssd1 vccd1 vccd1 _10880_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_158_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11789_ _11789_/A _11789_/B _11789_/C _11789_/D vssd1 vssd1 vccd1 vccd1 _11924_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_119_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13528_ _13528_/A _07550_/X vssd1 vssd1 vccd1 vccd1 _14104_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_158_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ _13459_/A _07731_/X vssd1 vssd1 vccd1 vccd1 _14035_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_154_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_71_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07951_ _07951_/A _07971_/B _07962_/C vssd1 vssd1 vccd1 vccd1 _07952_/A sky130_fd_sc_hd__or3_1
X_06902_ _07328_/A _07336_/B _07073_/C vssd1 vssd1 vccd1 vccd1 _06903_/A sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_86_clk_A _12438_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ _07882_/A vssd1 vssd1 vccd1 vccd1 _07882_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09621_ _09634_/A vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06833_ _06967_/A vssd1 vssd1 vccd1 vccd1 _06843_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_68_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09552_ _13461_/A _12314_/Q _09558_/S vssd1 vssd1 vccd1 vccd1 _09553_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06764_ _06764_/A vssd1 vssd1 vccd1 vccd1 _06764_/X sky130_fd_sc_hd__clkbuf_1
X_08503_ _08409_/X _08411_/X _08475_/X _08502_/X _08492_/X _08424_/X vssd1 vssd1 vccd1
+ vccd1 _08503_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11145__B _13935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09483_ _09513_/A vssd1 vssd1 vccd1 vccd1 _09483_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06695_ _06753_/A vssd1 vssd1 vccd1 vccd1 _06706_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08591__S0 _08556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ _11706_/C vssd1 vssd1 vccd1 vccd1 _13361_/A sky130_fd_sc_hd__buf_4
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13000__156 vssd1 vssd1 vccd1 vccd1 _13000__156/HI _13411_/A sky130_fd_sc_hd__conb_1
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ _08365_/A vssd1 vssd1 vccd1 vccd1 _08365_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10476__S _10480_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A _12881_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11161__A _13840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ _10512_/B vssd1 vssd1 vccd1 vccd1 _07993_/C sky130_fd_sc_hd__buf_2
XFILLER_165_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ _08296_/A vssd1 vssd1 vccd1 vccd1 _08296_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07247_ _07247_/A vssd1 vssd1 vccd1 vccd1 _07247_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_2_0_clk clkbuf_4_3_0_clk/A vssd1 vssd1 vccd1 vccd1 _12917_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_164_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_39_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07178_ _07178_/A vssd1 vssd1 vccd1 vccd1 _07178_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10224__B _13754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09819_ _09836_/A vssd1 vssd1 vccd1 vccd1 _09834_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10530__A1 _09763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12830_ _12835_/CLK _12830_/D vssd1 vssd1 vccd1 vccd1 _12830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12776_/CLK _12761_/D vssd1 vssd1 vccd1 vccd1 _12761_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08582__S0 _08556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13551__A _13551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11763_/S vssd1 vssd1 vccd1 vccd1 _11726_/S sky130_fd_sc_hd__buf_2
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12710_/CLK _12692_/D vssd1 vssd1 vccd1 vccd1 _13821_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11643_ _11649_/B _11643_/B _11649_/D vssd1 vssd1 vccd1 vccd1 _11643_/Y sky130_fd_sc_hd__nand3_1
XFILLER_42_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08364__B _08364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11574_ _11574_/A _11643_/B vssd1 vssd1 vccd1 vccd1 _12822_/D sky130_fd_sc_hd__nor2_1
Xinput17 peripheralBus_address[2] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10525_ _10538_/A vssd1 vssd1 vccd1 vccd1 _10525_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10456_ _13687_/A _12542_/Q _10456_/S vssd1 vssd1 vccd1 vccd1 _10457_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08380__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10387_ _10385_/X _10379_/X _10386_/X _10383_/X vssd1 vssd1 vccd1 vccd1 _12519_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_repeater122_A peripheralBus_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ _12132_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12127_/A sky130_fd_sc_hd__and2_1
XFILLER_96_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12057_ _12057_/A _12057_/B vssd1 vssd1 vccd1 vccd1 _12057_/Y sky130_fd_sc_hd__nor2_2
XFILLER_111_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11008_ _12675_/Q _13949_/A vssd1 vssd1 vccd1 vccd1 _11011_/B sky130_fd_sc_hd__xor2_1
XANTENNA_output51_A _13376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10521__A1 _09753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12959_ _12962_/CLK _12959_/D vssd1 vssd1 vccd1 vccd1 _12959_/Q sky130_fd_sc_hd__dfxtp_1
X_13294__450 vssd1 vssd1 vccd1 vccd1 _13294__450/HI _14015_/A sky130_fd_sc_hd__conb_1
XFILLER_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08573__S0 _08549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06480_ _06480_/A vssd1 vssd1 vccd1 vccd1 _06480_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08150_ _08150_/A vssd1 vssd1 vccd1 vccd1 _08184_/A sky130_fd_sc_hd__clkbuf_2
X_13335__491 vssd1 vssd1 vccd1 vccd1 _13335__491/HI _14088_/A sky130_fd_sc_hd__conb_1
XANTENNA__11412__C _11412_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07101_ _07108_/A _07105_/B _07101_/C vssd1 vssd1 vccd1 vccd1 _07102_/A sky130_fd_sc_hd__or3_1
X_08081_ _08081_/A _08113_/B _08087_/C vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__or3_1
X_07032_ _07032_/A vssd1 vssd1 vccd1 vccd1 _07032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08628__S1 _08551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ _10939_/C vssd1 vssd1 vccd1 vccd1 _13937_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_87_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07934_ _08166_/A vssd1 vssd1 vccd1 vccd1 _08004_/A sky130_fd_sc_hd__buf_2
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07865_ _07892_/A vssd1 vssd1 vccd1 vccd1 _07877_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_56_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _12313_/Q _13556_/A vssd1 vssd1 vccd1 vccd1 _09607_/B sky130_fd_sc_hd__xor2_1
XFILLER_44_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06816_ _10512_/B vssd1 vssd1 vccd1 vccd1 _07969_/B sky130_fd_sc_hd__buf_4
X_07796_ _07796_/A _07806_/B _07801_/C vssd1 vssd1 vccd1 vccd1 _07797_/A sky130_fd_sc_hd__or3_1
XFILLER_44_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09535_ _13456_/A _12309_/Q _09610_/B vssd1 vssd1 vccd1 vccd1 _09536_/B sky130_fd_sc_hd__mux2_1
X_06747_ _06747_/A vssd1 vssd1 vccd1 vccd1 _06747_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13371__A _13371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09466_ _12289_/Q _13565_/A vssd1 vssd1 vccd1 vccd1 _09467_/D sky130_fd_sc_hd__xnor2_1
X_06678_ _06686_/A _06678_/B _06678_/C vssd1 vssd1 vccd1 vccd1 _06679_/A sky130_fd_sc_hd__or3_1
XFILLER_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08417_ _08524_/A vssd1 vssd1 vccd1 vccd1 _08417_/X sky130_fd_sc_hd__clkbuf_4
X_09397_ _09397_/A _09397_/B _09397_/C _09397_/D vssd1 vssd1 vccd1 vccd1 _09400_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__08184__B _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10028__B1 _09978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ _08348_/A vssd1 vssd1 vccd1 vccd1 _08348_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08279_ _08288_/A _08285_/B vssd1 vssd1 vccd1 vccd1 _08280_/A sky130_fd_sc_hd__or2_1
XFILLER_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10310_ _10348_/S vssd1 vssd1 vccd1 vccd1 _10324_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_152_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11290_ _11160_/X _11284_/X _11289_/X _11195_/X vssd1 vssd1 vccd1 vccd1 _12745_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10241_ _12468_/Q _13743_/A vssd1 vssd1 vccd1 vccd1 _10242_/D sky130_fd_sc_hd__xor2_1
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10172_ _13616_/A _12469_/Q _10180_/S vssd1 vssd1 vccd1 vccd1 _10173_/B sky130_fd_sc_hd__mux2_1
XFILLER_160_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13931_ _13931_/A _06471_/X vssd1 vssd1 vccd1 vccd1 _13995_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13862_ _13862_/A _06663_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[23] sky130_fd_sc_hd__ebufn_8
X_13278__434 vssd1 vssd1 vccd1 vccd1 _13278__434/HI _13983_/A sky130_fd_sc_hd__conb_1
XFILLER_74_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12813_ _12813_/CLK _12813_/D vssd1 vssd1 vccd1 vccd1 _12813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13793_ _13793_/A _06856_/X vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _12780_/CLK _12744_/D vssd1 vssd1 vccd1 vccd1 _13871_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13319__475 vssd1 vssd1 vccd1 vccd1 _13319__475/HI _14056_/A sky130_fd_sc_hd__conb_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12699_/CLK _12675_/D vssd1 vssd1 vccd1 vccd1 _12675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11626_ _11626_/A _11626_/B _11626_/C _11626_/D vssd1 vssd1 vccd1 vccd1 _11628_/C
+ sky130_fd_sc_hd__and4_1
X_12992__148 vssd1 vssd1 vccd1 vccd1 _12992__148/HI _13389_/A sky130_fd_sc_hd__conb_1
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09918__B _09918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ _11557_/A vssd1 vssd1 vccd1 vccd1 _12818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10508_ _10508_/A vssd1 vssd1 vccd1 vccd1 _12550_/D sky130_fd_sc_hd__clkbuf_1
X_11488_ _11488_/A vssd1 vssd1 vccd1 vccd1 _12801_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09188__A1 _09186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10439_ _13682_/A _12537_/Q _10507_/B vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__mux2_1
XFILLER_143_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _12115_/A _12109_/B vssd1 vssd1 vccd1 vccd1 _12110_/A sky130_fd_sc_hd__and2_1
XFILLER_111_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07650_ _07650_/A vssd1 vssd1 vccd1 vccd1 _07650_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06601_ _06601_/A vssd1 vssd1 vccd1 vccd1 _06601_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07581_ _07581_/A vssd1 vssd1 vccd1 vccd1 _07581_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09320_ _09328_/A _09329_/A _09330_/A _09320_/D vssd1 vssd1 vccd1 vccd1 _09323_/B
+ sky130_fd_sc_hd__and4_1
X_06532_ _06534_/A _06540_/B _06540_/C vssd1 vssd1 vccd1 vccd1 _06533_/A sky130_fd_sc_hd__or3_1
XFILLER_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ _09251_/A _09251_/B vssd1 vssd1 vccd1 vccd1 _12240_/D sky130_fd_sc_hd__nor2_1
X_06463_ _06547_/A vssd1 vssd1 vccd1 vccd1 _07827_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08202_ _08212_/A _08208_/B _08212_/C vssd1 vssd1 vccd1 vccd1 _08203_/A sky130_fd_sc_hd__or3_1
XFILLER_21_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ _11184_/A vssd1 vssd1 vccd1 vccd1 _09182_/X sky130_fd_sc_hd__clkbuf_8
X_06394_ _06403_/A _06400_/B vssd1 vssd1 vccd1 vccd1 _06395_/A sky130_fd_sc_hd__or2_1
XFILLER_159_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13071__227 vssd1 vssd1 vccd1 vccd1 _13071__227/HI _13546_/A sky130_fd_sc_hd__conb_1
XFILLER_147_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08133_ _08135_/A _08189_/B _08138_/C vssd1 vssd1 vccd1 vccd1 _08134_/A sky130_fd_sc_hd__or3_1
XFILLER_107_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07629__A _08022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _08064_/A vssd1 vssd1 vccd1 vccd1 _08077_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_134_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13112__268 vssd1 vssd1 vccd1 vccd1 _13112__268/HI _13637_/A sky130_fd_sc_hd__conb_1
X_07015_ _07019_/A _07019_/B vssd1 vssd1 vccd1 vccd1 _07016_/A sky130_fd_sc_hd__or2_1
XFILLER_161_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09844__A _10173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10733__A1 _10288_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13366__A _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ _11518_/B _12810_/Q _12811_/Q _12812_/Q _08941_/X _08942_/X vssd1 vssd1 vccd1
+ vccd1 _08966_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09026__S1 _08968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07917_ _07921_/A _07917_/B _07917_/C vssd1 vssd1 vccd1 vccd1 _07918_/A sky130_fd_sc_hd__or3_1
XFILLER_29_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10502__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ _10165_/B vssd1 vssd1 vccd1 vccd1 _13756_/A sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_95_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _12377_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07848_ _07962_/A _07854_/B _07852_/C vssd1 vssd1 vccd1 vccd1 _07849_/A sky130_fd_sc_hd__or3_1
XFILLER_44_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13006__162 vssd1 vssd1 vccd1 vccd1 _13006__162/HI _13417_/A sky130_fd_sc_hd__conb_1
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07779_ _07782_/A _07779_/B _07787_/C vssd1 vssd1 vccd1 vccd1 _07780_/A sky130_fd_sc_hd__or3_1
XANTENNA__08537__S0 _09140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ _13434_/A _09513_/X _09517_/X _09509_/X vssd1 vssd1 vccd1 vccd1 _12303_/D
+ sky130_fd_sc_hd__o211a_1
X_10790_ _10865_/A _10865_/B _10790_/C vssd1 vssd1 vccd1 vccd1 _10795_/B sky130_fd_sc_hd__and3_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09455_/A _09449_/B vssd1 vssd1 vccd1 vccd1 _09450_/A sky130_fd_sc_hd__and2_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _12461_/CLK _12460_/D vssd1 vssd1 vccd1 vccd1 _12460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11411_ _11438_/A vssd1 vssd1 vccd1 vccd1 _11411_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12391_ _12404_/CLK _12391_/D vssd1 vssd1 vccd1 vccd1 _13519_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11342_ _11381_/S vssd1 vssd1 vccd1 vccd1 _11356_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12164__B _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11273_ _11273_/A _11273_/B _11273_/C _11273_/D vssd1 vssd1 vccd1 vccd1 _11279_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_152_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14061_ _14061_/A _07944_/X vssd1 vssd1 vccd1 vccd1 _14125_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_165_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10224_ _12479_/Q _13754_/A vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__xor2_1
XFILLER_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10155_ _12466_/Q _10155_/B _10155_/C vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__and3_1
XFILLER_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10086_ _10097_/A _10086_/B _10086_/C _10100_/A vssd1 vssd1 vccd1 vccd1 _10089_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_86_clk _12438_/CLK vssd1 vssd1 vccd1 vccd1 _12443_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08089__B _08089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13914_ _13914_/A _06518_/X vssd1 vssd1 vccd1 vccd1 _13978_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_114_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13845_ _13845_/A _06711_/X vssd1 vssd1 vccd1 vccd1 _14069_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11524__A _11680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13776_ _13776_/A _06903_/X vssd1 vssd1 vccd1 vccd1 _14096_/Z sky130_fd_sc_hd__ebufn_8
X_10988_ _10988_/A vssd1 vssd1 vccd1 vccd1 _11206_/A sky130_fd_sc_hd__buf_2
XANTENNA__06618__A _06694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12727_ _12743_/CLK _12727_/D vssd1 vssd1 vccd1 vccd1 _12727_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09929__A _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12658_ _12659_/CLK _12658_/D vssd1 vssd1 vccd1 vccd1 _12658_/Q sky130_fd_sc_hd__dfxtp_1
X_11609_ _11609_/A _11609_/B vssd1 vssd1 vccd1 vccd1 _12831_/D sky130_fd_sc_hd__nor2_1
X_12589_ _12589_/CLK _12589_/D vssd1 vssd1 vccd1 vccd1 _13716_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_10_clk _12217_/CLK vssd1 vssd1 vccd1 vccd1 _12962_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07449__A _07473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _12642_/Q vssd1 vssd1 vccd1 vccd1 _10875_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09008__S1 _08947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08751_ _12630_/Q vssd1 vssd1 vccd1 vccd1 _10874_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _12505_/CLK sky130_fd_sc_hd__clkbuf_16
X_07702_ _07714_/A _07710_/B _07704_/C vssd1 vssd1 vccd1 vccd1 _07703_/A sky130_fd_sc_hd__or3_1
X_08682_ _08679_/X _08681_/X _08682_/S vssd1 vssd1 vccd1 vccd1 _09398_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07633_ _07644_/A _07641_/B _07635_/C vssd1 vssd1 vccd1 vccd1 _07634_/A sky130_fd_sc_hd__or3_1
XFILLER_81_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07564_ _07575_/A _08103_/B _07564_/C vssd1 vssd1 vccd1 vccd1 _07565_/A sky130_fd_sc_hd__or3_1
XFILLER_41_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09303_ _09320_/D vssd1 vssd1 vccd1 vccd1 _09330_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06515_ _08210_/A vssd1 vssd1 vccd1 vccd1 _07507_/A sky130_fd_sc_hd__buf_4
XFILLER_34_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08844__A0 _08782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ _07495_/A vssd1 vssd1 vccd1 vccd1 _07495_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06446_ _06446_/A vssd1 vssd1 vccd1 vccd1 _06446_/X sky130_fd_sc_hd__clkbuf_1
X_09234_ _09234_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _12236_/D sky130_fd_sc_hd__nor2_1
XFILLER_22_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08743__A _13777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09165_ _09631_/A vssd1 vssd1 vccd1 vccd1 _10659_/A sky130_fd_sc_hd__buf_4
X_06377_ input18/X _12059_/A _06377_/C vssd1 vssd1 vccd1 vccd1 _06725_/A sky130_fd_sc_hd__or3_1
X_08116_ _08122_/A _08128_/B _08122_/C vssd1 vssd1 vccd1 vccd1 _08117_/A sky130_fd_sc_hd__or3_1
XFILLER_108_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ input19/X _09096_/B _09096_/C input18/X vssd1 vssd1 vccd1 vccd1 _12059_/B
+ sky130_fd_sc_hd__or4b_2
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08047_ _08052_/A _08047_/B _08057_/C vssd1 vssd1 vccd1 vccd1 _08048_/A sky130_fd_sc_hd__or3_1
XFILLER_135_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09998_ _10112_/A _10030_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10008_/D sky130_fd_sc_hd__and3_1
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08949_ _12818_/Q vssd1 vssd1 vccd1 vccd1 _11562_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_68_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _12517_/CLK sky130_fd_sc_hd__clkbuf_16
X_11960_ _11977_/S vssd1 vssd1 vccd1 vccd1 _11974_/S sky130_fd_sc_hd__buf_2
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07822__A _07822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ _10906_/Y _10904_/C _10910_/X vssd1 vssd1 vccd1 vccd1 _12652_/D sky130_fd_sc_hd__a21oi_1
X_13240__396 vssd1 vssd1 vccd1 vccd1 _13240__396/HI _13895_/A sky130_fd_sc_hd__conb_1
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11891_ _11891_/A vssd1 vssd1 vccd1 vccd1 _12899_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09740__C _10637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13630_ _13630_/A _07280_/X vssd1 vssd1 vccd1 vccd1 _14078_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_44_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10842_ _10848_/C _10917_/B _10842_/C vssd1 vssd1 vccd1 vccd1 _10843_/A sky130_fd_sc_hd__and3b_1
XANTENNA__12159__B _13372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__C _08360_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ _13561_/A _07465_/X vssd1 vssd1 vccd1 vccd1 _13625_/Z sky130_fd_sc_hd__ebufn_8
X_10773_ _10864_/C _10773_/B _10863_/C _10773_/D vssd1 vssd1 vccd1 vccd1 _10809_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_158_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12512_ _12517_/CLK _12512_/D vssd1 vssd1 vccd1 vccd1 _12512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13492_ _13492_/A _07645_/X vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_9_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12443_ _12443_/CLK _12443_/D vssd1 vssd1 vccd1 vccd1 _12443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11198__A1 _10548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12374_ _12377_/CLK _12374_/D vssd1 vssd1 vccd1 vccd1 _12374_/Q sky130_fd_sc_hd__dfxtp_1
X_13134__290 vssd1 vssd1 vccd1 vccd1 _13134__290/HI _13675_/A sky130_fd_sc_hd__conb_1
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14113_ _14113_/A _08245_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11325_ _13886_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11325_/X sky130_fd_sc_hd__or2_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11256_ _11256_/A vssd1 vssd1 vccd1 vccd1 _12742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14044_ _14044_/A _07898_/X vssd1 vssd1 vccd1 vccd1 _14108_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_106_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06901__A _07090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _13626_/A _12479_/Q _10214_/S vssd1 vssd1 vccd1 vccd1 _10208_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11519__A _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ _13849_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11187_/X sky130_fd_sc_hd__or2_1
XFILLER_121_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10138_ _10137_/B _10126_/D _10137_/D _10148_/C vssd1 vssd1 vccd1 vccd1 _10139_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _12829_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10069_ _10086_/B _10076_/D vssd1 vssd1 vccd1 vccd1 _10070_/C sky130_fd_sc_hd__nand2_1
XFILLER_48_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13828_ _13828_/A _06757_/X vssd1 vssd1 vccd1 vccd1 _13988_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_63_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12998__154 vssd1 vssd1 vccd1 vccd1 _12998__154/HI _13409_/A sky130_fd_sc_hd__conb_1
XFILLER_16_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13759_ _13759_/A _06945_/X vssd1 vssd1 vccd1 vccd1 _14079_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06300_ _06300_/A vssd1 vssd1 vccd1 vccd1 _06300_/X sky130_fd_sc_hd__clkbuf_1
X_07280_ _07280_/A vssd1 vssd1 vccd1 vccd1 _07280_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07179__A _07205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09394__A _09967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09921_ _09934_/S vssd1 vssd1 vccd1 vccd1 _09921_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07907__A _07920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183__339 vssd1 vssd1 vccd1 vccd1 _13183__339/HI _13790_/A sky130_fd_sc_hd__conb_1
X_09852_ _12387_/Q _13564_/A vssd1 vssd1 vccd1 vccd1 _09852_/Y sky130_fd_sc_hd__xnor2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater84_A peripheralBus_data[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _12626_/Q vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09783_ _13499_/A _09787_/B vssd1 vssd1 vccd1 vccd1 _09783_/X sky130_fd_sc_hd__or2_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06995_ _06995_/A _06995_/B vssd1 vssd1 vccd1 vccd1 _06996_/A sky130_fd_sc_hd__or2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08734_ _13777_/A vssd1 vssd1 vccd1 vccd1 _08887_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_100_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _12456_/Q vssd1 vssd1 vccd1 vccd1 _10130_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _07616_/A _07626_/B _07621_/C vssd1 vssd1 vccd1 vccd1 _07617_/A sky130_fd_sc_hd__or3_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _08588_/X _08591_/X _08593_/X _08595_/X _08583_/X _08563_/X vssd1 vssd1 vccd1
+ vccd1 _08596_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13077__233 vssd1 vssd1 vccd1 vccd1 _13077__233/HI _13572_/A sky130_fd_sc_hd__conb_1
X_07547_ _07590_/A vssd1 vssd1 vccd1 vccd1 _07558_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07478_ _07478_/A _07484_/B vssd1 vssd1 vccd1 vccd1 _07479_/A sky130_fd_sc_hd__or2_1
XFILLER_10_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09217_ _09271_/C vssd1 vssd1 vccd1 vccd1 _09217_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13118__274 vssd1 vssd1 vccd1 vccd1 _13118__274/HI _13643_/A sky130_fd_sc_hd__conb_1
X_06429_ _06429_/A vssd1 vssd1 vccd1 vccd1 _06429_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09148_ _11490_/A vssd1 vssd1 vccd1 vccd1 _09148_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09079_ _10941_/B vssd1 vssd1 vccd1 vccd1 _11386_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11110_ _11110_/A vssd1 vssd1 vccd1 vccd1 _12704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12090_ _14073_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12090_/X sky130_fd_sc_hd__or2_1
X_11041_ _11055_/A vssd1 vssd1 vccd1 vccd1 _11041_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13554__A _13554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input13_A peripheralBus_address[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11943_ _11977_/S vssd1 vssd1 vccd1 vccd1 _11957_/S sky130_fd_sc_hd__buf_2
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11874_ _11874_/A vssd1 vssd1 vccd1 vccd1 _12894_/D sky130_fd_sc_hd__clkbuf_1
X_13613_ _13613_/A _07329_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
X_10825_ _10825_/A _10825_/B vssd1 vssd1 vccd1 vccd1 _12632_/D sky130_fd_sc_hd__nor2_1
XANTENNA__12065__C1 _11497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13544_ _13544_/A _07505_/X vssd1 vssd1 vccd1 vccd1 _13992_/Z sky130_fd_sc_hd__ebufn_8
X_10756_ _10773_/D vssd1 vssd1 vccd1 vccd1 _10863_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13475_ _13475_/A _07687_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
X_10687_ _10552_/X _10673_/A _10686_/X _10682_/X vssd1 vssd1 vccd1 vccd1 _12599_/D
+ sky130_fd_sc_hd__o211a_1
X_12426_ _12659_/CLK _12426_/D vssd1 vssd1 vccd1 vccd1 _12426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09784__A1 _09092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ _12367_/CLK _12357_/D vssd1 vssd1 vccd1 vccd1 _13568_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_154_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11308_ _13879_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11308_/X sky130_fd_sc_hd__or2_1
XFILLER_141_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12288_ _12290_/CLK _12288_/D vssd1 vssd1 vccd1 vccd1 _12288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14027_ _14027_/A _08061_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
X_11239_ _11239_/A _11239_/B vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__and2_1
XFILLER_68_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06780_ _06788_/A _06780_/B _06780_/C vssd1 vssd1 vccd1 vccd1 _06781_/A sky130_fd_sc_hd__or3_1
XFILLER_36_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11646__A2 _11649_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08450_ _08437_/X _08439_/X _08443_/X _08447_/X _08448_/X _08449_/X vssd1 vssd1 vccd1
+ vccd1 _08450_/X sky130_fd_sc_hd__mux4_1
X_07401_ _07822_/A _07404_/B _07401_/C vssd1 vssd1 vccd1 vccd1 _07402_/A sky130_fd_sc_hd__or3_1
X_08381_ _12240_/Q _12241_/Q _12242_/Q _12243_/Q _08379_/X _08380_/X vssd1 vssd1 vccd1
+ vccd1 _08381_/X sky130_fd_sc_hd__mux4_2
XFILLER_90_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07332_ _07332_/A vssd1 vssd1 vccd1 vccd1 _07332_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11712__A _11763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09389__A _09389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06806__A _07857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07263_ _07266_/A _07263_/B _07273_/C vssd1 vssd1 vccd1 vccd1 _07264_/A sky130_fd_sc_hd__or3_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ _11641_/C _12831_/Q _11640_/B _11641_/B _08967_/X _08968_/X vssd1 vssd1 vccd1
+ vccd1 _09002_/X sky130_fd_sc_hd__mux4_2
X_07194_ _07194_/A vssd1 vssd1 vccd1 vccd1 _07194_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09775__A1 _09773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07637__A _09484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09904_ _13529_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09904_/X sky130_fd_sc_hd__or2_1
XFILLER_59_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09835_ _09835_/A vssd1 vssd1 vccd1 vccd1 _12386_/D sky130_fd_sc_hd__clkbuf_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input5_A peripheralBus_address[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13374__A _13374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _09763_/X _09759_/X _09764_/X _09765_/X vssd1 vssd1 vccd1 vccd1 _12364_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06978_ _06978_/A vssd1 vssd1 vccd1 vccd1 _06978_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08717_ _08714_/X _08716_/X _09941_/A vssd1 vssd1 vccd1 vccd1 _09399_/B sky130_fd_sc_hd__mux2_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09697_ _09697_/A vssd1 vssd1 vccd1 vccd1 _12351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _08637_/X _08640_/X _08643_/X _08646_/X _08632_/X _08647_/X vssd1 vssd1 vccd1
+ vccd1 _08648_/X sky130_fd_sc_hd__mux4_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _13585_/A vssd1 vssd1 vccd1 vccd1 _08579_/X sky130_fd_sc_hd__buf_2
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10610_/A vssd1 vssd1 vccd1 vccd1 _12582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11590_ _11590_/A _11590_/B vssd1 vssd1 vccd1 vccd1 _12826_/D sky130_fd_sc_hd__nor2_1
X_10541_ _10408_/X _10538_/X _10540_/X _10536_/X vssd1 vssd1 vccd1 vccd1 _12561_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10472_ _10472_/A vssd1 vssd1 vccd1 vccd1 _12546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09766__A1 _09763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ _12968_/CLK _12211_/D vssd1 vssd1 vccd1 vccd1 _14108_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07547__A _07590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ _12964_/Q _14106_/A _12151_/S vssd1 vssd1 vccd1 vccd1 _12143_/B sky130_fd_sc_hd__mux2_1
XFILLER_135_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12172__B _13364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ _14067_/A _12073_/B vssd1 vssd1 vccd1 vccd1 _12073_/X sky130_fd_sc_hd__or2_1
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11024_ _11039_/A vssd1 vssd1 vccd1 vccd1 _11024_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12975_ _12980_/CLK _12975_/D vssd1 vssd1 vccd1 vccd1 _14100_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11926_ _14063_/Z _14031_/A _11940_/S vssd1 vssd1 vccd1 vccd1 _11927_/B sky130_fd_sc_hd__mux2_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _11857_/A vssd1 vssd1 vccd1 vccd1 _12889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10808_ _10864_/A _10864_/B _10865_/C _10865_/D vssd1 vssd1 vccd1 vccd1 _10809_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_60_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11788_ _13378_/A _11787_/Y _11711_/B _09404_/A _13404_/A vssd1 vssd1 vccd1 vccd1
+ _12870_/D sky130_fd_sc_hd__o2111a_1
XFILLER_41_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13527_ _13527_/A _07552_/X vssd1 vssd1 vccd1 vccd1 _13623_/Z sky130_fd_sc_hd__ebufn_8
X_10739_ _10820_/C vssd1 vssd1 vccd1 vccd1 _10895_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__09937__A _09937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ _13458_/A _07733_/X vssd1 vssd1 vccd1 vccd1 _14034_/Z sky130_fd_sc_hd__ebufn_8
X_12409_ _12470_/CLK _12409_/D vssd1 vssd1 vccd1 vccd1 _13585_/A sky130_fd_sc_hd__dfxtp_1
X_13389_ _13389_/A _08348_/X vssd1 vssd1 vccd1 vccd1 _14125_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07950_ _08004_/A vssd1 vssd1 vccd1 vccd1 _07962_/C sky130_fd_sc_hd__buf_2
XFILLER_141_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09672__A _09711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06901_ _07090_/A vssd1 vssd1 vccd1 vccd1 _07073_/C sky130_fd_sc_hd__clkbuf_2
X_07881_ _07881_/A _07890_/B _07890_/C vssd1 vssd1 vccd1 vccd1 _07882_/A sky130_fd_sc_hd__or3_1
XFILLER_110_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09620_ _09620_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09620_/X sky130_fd_sc_hd__or2_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06832_ _06832_/A vssd1 vssd1 vccd1 vccd1 _06843_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07192__A _07205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _09551_/A vssd1 vssd1 vccd1 vccd1 _12313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06763_ _06775_/A _06765_/B _06765_/C vssd1 vssd1 vccd1 vccd1 _06764_/A sky130_fd_sc_hd__or3_1
X_08502_ _09362_/B _12266_/Q _12267_/Q _12268_/Q _08368_/X _08370_/X vssd1 vssd1 vccd1
+ vccd1 _08502_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13922__A _13922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10827__B1 _10781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09482_ _11026_/B _09873_/B _10637_/B vssd1 vssd1 vccd1 vccd1 _09513_/A sky130_fd_sc_hd__nor3_4
X_06694_ _06694_/A vssd1 vssd1 vccd1 vccd1 _06753_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07920__A _07920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08433_ _08425_/X _08432_/X _08498_/S vssd1 vssd1 vccd1 vccd1 _11706_/C sky130_fd_sc_hd__mux2_2
XANTENNA__08591__S1 _08557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ _08364_/A _08364_/B _08364_/C vssd1 vssd1 vccd1 vccd1 _08365_/A sky130_fd_sc_hd__or3_1
XANTENNA__06536__A _06688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11788__D1 _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ _07315_/A vssd1 vssd1 vccd1 vccd1 _07315_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08295_ _08300_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08296_/A sky130_fd_sc_hd__or2_1
XFILLER_149_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07246_ _07253_/A _07250_/B _07246_/C vssd1 vssd1 vccd1 vccd1 _07247_/A sky130_fd_sc_hd__or3_1
XFILLER_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13369__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189__345 vssd1 vssd1 vccd1 vccd1 _13189__345/HI _13796_/A sky130_fd_sc_hd__conb_1
X_07177_ _07180_/A _07177_/B _07187_/C vssd1 vssd1 vccd1 vccd1 _07178_/A sky130_fd_sc_hd__or3_1
XFILLER_118_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10108__C_N _09987_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11307__A1 _10662_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09818_ _09818_/A vssd1 vssd1 vccd1 vccd1 _12381_/D sky130_fd_sc_hd__clkbuf_1
X_09749_ _09139_/X _09741_/X _09747_/X _09748_/X vssd1 vssd1 vccd1 vccd1 _12359_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10240__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12776_/CLK _12760_/D vssd1 vssd1 vccd1 vccd1 _12760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _13404_/A _11711_/B vssd1 vssd1 vccd1 vccd1 _11763_/S sky130_fd_sc_hd__nand2_4
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10294__A1 _09120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07830__A _09125_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08582__S1 _08557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12710_/CLK _12691_/D vssd1 vssd1 vccd1 vccd1 _13820_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11642_/A _11642_/B _11642_/C _11642_/D vssd1 vssd1 vccd1 vccd1 _11649_/D
+ sky130_fd_sc_hd__and4_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12167__B _13361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11573_ _11689_/A _11649_/C vssd1 vssd1 vccd1 vccd1 _11643_/B sky130_fd_sc_hd__and2_1
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 peripheralBus_address[3] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10524_ _09756_/X _10511_/X _10522_/X _10523_/X vssd1 vssd1 vccd1 vccd1 _12555_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09476__B _13562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ _10455_/A vssd1 vssd1 vccd1 vccd1 _12541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10386_ _13648_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10386_/X sky130_fd_sc_hd__or2_1
XFILLER_123_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12125_ _12959_/Q _14101_/A _12135_/S vssd1 vssd1 vccd1 vccd1 _12126_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater115_A _14112_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09492__A _09623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ _12056_/A _12056_/B _12056_/C vssd1 vssd1 vccd1 vccd1 _12057_/B sky130_fd_sc_hd__or3_1
XFILLER_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11007_ _12671_/Q _13945_/A vssd1 vssd1 vccd1 vccd1 _11011_/A sky130_fd_sc_hd__xor2_1
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output44_A _13375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12958_ _12962_/CLK _12958_/D vssd1 vssd1 vccd1 vccd1 _12958_/Q sky130_fd_sc_hd__dfxtp_1
X_13023__179 vssd1 vssd1 vccd1 vccd1 _13023__179/HI _13450_/A sky130_fd_sc_hd__conb_1
XFILLER_18_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08573__S1 _08551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909_ _12901_/Q _13373_/A vssd1 vssd1 vccd1 vccd1 _11910_/D sky130_fd_sc_hd__xor2_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _12895_/CLK _12889_/D vssd1 vssd1 vccd1 vccd1 _12889_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07100_ _07100_/A vssd1 vssd1 vccd1 vccd1 _07100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_158_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ _11026_/B vssd1 vssd1 vccd1 vccd1 _08113_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_146_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07031_ _07031_/A _07031_/B vssd1 vssd1 vccd1 vccd1 _07032_/A sky130_fd_sc_hd__or2_1
XFILLER_162_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10606__A _10952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08982_ _08973_/X _08981_/X _09043_/S vssd1 vssd1 vccd1 vccd1 _10939_/C sky130_fd_sc_hd__mux2_2
XFILLER_114_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07933_ _11154_/B vssd1 vssd1 vccd1 vccd1 _07945_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_96_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07864_ _07864_/A vssd1 vssd1 vccd1 vccd1 _07864_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09603_ _12308_/Q _13551_/A vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11156__B _11156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06815_ _06983_/B vssd1 vssd1 vccd1 vccd1 _10512_/B sky130_fd_sc_hd__clkbuf_2
X_07795_ _08064_/A vssd1 vssd1 vccd1 vccd1 _07806_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_37_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09534_ _09534_/A vssd1 vssd1 vccd1 vccd1 _12308_/D sky130_fd_sc_hd__clkbuf_1
X_06746_ _06746_/A _06751_/B _06751_/C vssd1 vssd1 vccd1 vccd1 _06747_/A sky130_fd_sc_hd__or3_1
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08746__A _13777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09465_ _12278_/Q _13554_/A vssd1 vssd1 vccd1 vccd1 _09467_/C sky130_fd_sc_hd__xnor2_1
X_06677_ _06677_/A vssd1 vssd1 vccd1 vccd1 _06677_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11172__A _11199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08416_ _12230_/Q vssd1 vssd1 vccd1 vccd1 _09210_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09396_ _09867_/B _09396_/B _09396_/C _09396_/D vssd1 vssd1 vccd1 vccd1 _09400_/A
+ sky130_fd_sc_hd__or4_1
XANTENNA__06266__A _06377_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08347_ _08347_/A _08349_/B vssd1 vssd1 vccd1 vccd1 _08348_/A sky130_fd_sc_hd__or2_1
X_08278_ _08314_/A vssd1 vssd1 vccd1 vccd1 _08288_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_153_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07229_ _07229_/A vssd1 vssd1 vccd1 vccd1 _07229_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10240_ _12473_/Q _13748_/A vssd1 vssd1 vccd1 vccd1 _10242_/C sky130_fd_sc_hd__xor2_1
XFILLER_154_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10235__B _13745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10171_ _10171_/A vssd1 vssd1 vccd1 vccd1 _12468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07825__A _09125_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09743__C _11156_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13930_ _13930_/A _06473_/X vssd1 vssd1 vccd1 vccd1 _13994_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10251__A _11028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13861_ _13861_/A _06665_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
XFILLER_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13562__A _13562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ _12813_/CLK _12812_/D vssd1 vssd1 vccd1 vccd1 _12812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13792_ _13792_/A _06858_/X vssd1 vssd1 vccd1 vccd1 _14112_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__07560__A _07590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10267__A1 _09160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_70_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ _12743_/CLK _12743_/D vssd1 vssd1 vccd1 vccd1 _13952_/A sky130_fd_sc_hd__dfxtp_4
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12710_/CLK _12674_/D vssd1 vssd1 vccd1 vccd1 _12674_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11625_ _11625_/A _11625_/B _11625_/C _11625_/D vssd1 vssd1 vccd1 vccd1 _11628_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11556_ _11703_/A _11556_/B _11556_/C vssd1 vssd1 vccd1 vccd1 _11557_/A sky130_fd_sc_hd__and3_1
XANTENNA__06904__A _06913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ _11151_/A _10507_/B _10507_/C vssd1 vssd1 vccd1 vccd1 _10508_/A sky130_fd_sc_hd__and3_1
XFILLER_7_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11487_ _11490_/A _11487_/B vssd1 vssd1 vccd1 vccd1 _11488_/A sky130_fd_sc_hd__or2_1
XFILLER_109_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ _10438_/A vssd1 vssd1 vccd1 vccd1 _12536_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12192__A1 _10652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _12505_/Q _13747_/A vssd1 vssd1 vccd1 vccd1 _10372_/B sky130_fd_sc_hd__xor2_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _12954_/Q _14096_/A _12118_/S vssd1 vssd1 vccd1 vccd1 _12109_/B sky130_fd_sc_hd__mux2_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_23_clk_A _12881_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__C1 _09263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ _12921_/Q _13360_/A vssd1 vssd1 vccd1 vccd1 _12040_/D sky130_fd_sc_hd__xor2_1
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_clk clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_06600_ _06610_/A _06602_/B _06602_/C vssd1 vssd1 vccd1 vccd1 _06601_/A sky130_fd_sc_hd__or3_1
XFILLER_92_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07580_ _07588_/A _07585_/B _07580_/C vssd1 vssd1 vccd1 vccd1 _07581_/A sky130_fd_sc_hd__or3_1
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_38_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06531_ _06531_/A vssd1 vssd1 vccd1 vccd1 _06531_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09250_ _09315_/B _09253_/C vssd1 vssd1 vccd1 vccd1 _09251_/B sky130_fd_sc_hd__and2_1
X_06462_ _06462_/A vssd1 vssd1 vccd1 vccd1 _06729_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11207__A0 _13872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08201_ _08228_/A vssd1 vssd1 vccd1 vccd1 _08212_/C sky130_fd_sc_hd__clkbuf_1
X_06393_ _07861_/A vssd1 vssd1 vccd1 vccd1 _06403_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09181_ _13625_/Z vssd1 vssd1 vccd1 vccd1 _11184_/A sky130_fd_sc_hd__buf_4
XANTENNA__11720__A _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ _08132_/A vssd1 vssd1 vccd1 vccd1 _08132_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08063_ _08063_/A vssd1 vssd1 vccd1 vccd1 _08063_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07014_ _07014_/A vssd1 vssd1 vccd1 vccd1 _07014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08482__S0 _08373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10733__A2 _10703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ _11388_/B vssd1 vssd1 vccd1 vccd1 _13936_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07916_ _07916_/A vssd1 vssd1 vccd1 vccd1 _07916_/X sky130_fd_sc_hd__clkbuf_1
X_08896_ _08892_/X _08895_/X _10710_/A vssd1 vssd1 vccd1 vccd1 _10165_/B sky130_fd_sc_hd__mux2_1
XFILLER_130_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07847_ _07964_/A vssd1 vssd1 vccd1 vccd1 _07962_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07778_ _07778_/A vssd1 vssd1 vccd1 vccd1 _07778_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09517_ _11189_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09517_/X sky130_fd_sc_hd__or2_1
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08537__S1 _09146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06729_ _06729_/A _07323_/B _06738_/C vssd1 vssd1 vccd1 vccd1 _06730_/A sky130_fd_sc_hd__or3_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13351__507 vssd1 vssd1 vccd1 vccd1 _13351__507/HI _14120_/A sky130_fd_sc_hd__conb_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09448_ _13436_/A _12288_/Q _09448_/S vssd1 vssd1 vccd1 vccd1 _09449_/B sky130_fd_sc_hd__mux2_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _09379_/A _09379_/B vssd1 vssd1 vccd1 vccd1 _09380_/C sky130_fd_sc_hd__nand2_1
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ _11410_/A _11412_/B _11410_/C vssd1 vssd1 vccd1 vccd1 _11438_/A sky130_fd_sc_hd__or3_2
XFILLER_165_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12390_ _12414_/CLK _12390_/D vssd1 vssd1 vccd1 vccd1 _13567_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_20_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11341_ _11341_/A vssd1 vssd1 vccd1 vccd1 _12763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14060_ _14060_/A _07942_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[29] sky130_fd_sc_hd__ebufn_8
X_11272_ _12729_/Q _13937_/A vssd1 vssd1 vccd1 vccd1 _11273_/D sky130_fd_sc_hd__xor2_1
XFILLER_141_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13557__A _13557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ _12481_/Q _13756_/A vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__xor2_1
XFILLER_106_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245__401 vssd1 vssd1 vccd1 vccd1 _13245__401/HI _13900_/A sky130_fd_sc_hd__conb_1
XFILLER_121_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10154_ _10155_/B _10155_/C _10153_/Y _09987_/X vssd1 vssd1 vccd1 vccd1 _12465_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10085_ _10085_/A vssd1 vssd1 vccd1 vccd1 _12449_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09770__A _10665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13913_ _13913_/A _06520_/X vssd1 vssd1 vccd1 vccd1 _14009_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_75_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13844_ _13844_/A _06713_/X vssd1 vssd1 vccd1 vccd1 _14068_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13775_ _13775_/A _07957_/X vssd1 vssd1 vccd1 vccd1 _13775_/Z sky130_fd_sc_hd__ebufn_8
X_10987_ _10987_/A vssd1 vssd1 vccd1 vccd1 _12673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12726_ _12726_/CLK _12726_/D vssd1 vssd1 vccd1 vccd1 _13854_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ _12659_/CLK _12657_/D vssd1 vssd1 vccd1 vccd1 _12657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11540__A _11582_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11608_ _11640_/C _11610_/C _11540_/X vssd1 vssd1 vccd1 vccd1 _11609_/B sky130_fd_sc_hd__o21ai_1
XFILLER_156_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12588_ _12589_/CLK _12588_/D vssd1 vssd1 vccd1 vccd1 _13715_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11539_ _11627_/D _11547_/D vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__and2_1
XFILLER_128_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09945__A _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08736_/X _08741_/X _08744_/X _08747_/X _08748_/X _08749_/X vssd1 vssd1 vccd1
+ vccd1 _08750_/X sky130_fd_sc_hd__mux4_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13029__185 vssd1 vssd1 vccd1 vccd1 _13029__185/HI _13472_/A sky130_fd_sc_hd__conb_1
X_07701_ _07729_/A vssd1 vssd1 vccd1 vccd1 _07714_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08681_ _08567_/X _08568_/X _08654_/X _08680_/X _08583_/X _08584_/X vssd1 vssd1 vccd1
+ vccd1 _08681_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08541__A0 _08447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ _07661_/A vssd1 vssd1 vccd1 vccd1 _07644_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__06809__A _06809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ _07563_/A vssd1 vssd1 vccd1 vccd1 _07563_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09302_ _09306_/C _09302_/B vssd1 vssd1 vccd1 vccd1 _12253_/D sky130_fd_sc_hd__nor2_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06514_ _06528_/A vssd1 vssd1 vccd1 vccd1 _06526_/B sky130_fd_sc_hd__clkbuf_1
X_07494_ _07504_/A _07504_/B _07496_/C vssd1 vssd1 vccd1 vccd1 _07495_/A sky130_fd_sc_hd__or3_1
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ _09317_/D _09235_/C _09217_/X vssd1 vssd1 vccd1 vccd1 _09234_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10651__A1 _10648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06445_ _06451_/A _06449_/B vssd1 vssd1 vccd1 vccd1 _06446_/A sky130_fd_sc_hd__or2_1
XFILLER_139_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09164_ peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 _09631_/A sky130_fd_sc_hd__buf_4
XFILLER_21_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06376_ input17/X vssd1 vssd1 vccd1 vccd1 _12059_/A sky130_fd_sc_hd__inv_2
XANTENNA__06544__A _07507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10403__A1 _09767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08115_ _11026_/B vssd1 vssd1 vccd1 vccd1 _08128_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_119_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11600__B1 _11505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ _10250_/A vssd1 vssd1 vccd1 vccd1 _12060_/A sky130_fd_sc_hd__buf_2
XFILLER_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08046_ _08072_/A vssd1 vssd1 vccd1 vccd1 _08057_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_135_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13377__A _13377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08455__S0 _08373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09997_ _09997_/A _09997_/B _09997_/C _09997_/D vssd1 vssd1 vccd1 vccd1 _10030_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08948_ _12812_/Q _12813_/Q _11626_/C _11571_/D _08946_/X _08947_/X vssd1 vssd1 vccd1
+ vccd1 _08948_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08879_ _10922_/A _10921_/C _12655_/Q _12656_/Q _08779_/X _08780_/X vssd1 vssd1 vccd1
+ vccd1 _08879_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10910_ _10872_/A _10909_/X _10820_/C vssd1 vssd1 vccd1 vccd1 _10910_/X sky130_fd_sc_hd__a21bo_1
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07822__B _07822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ _11927_/A _11890_/B vssd1 vssd1 vccd1 vccd1 _11891_/A sky130_fd_sc_hd__and2_1
XFILLER_84_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10841_ _10869_/B _10833_/A _10877_/A _10876_/C vssd1 vssd1 vccd1 vccd1 _10842_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13840__A _13840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13560_ _13560_/A _07467_/X vssd1 vssd1 vccd1 vccd1 _14104_/Z sky130_fd_sc_hd__ebufn_8
X_10772_ _12622_/Q vssd1 vssd1 vccd1 vccd1 _10865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12511_ _12517_/CLK _12511_/D vssd1 vssd1 vccd1 vccd1 _12511_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10642__A1 _10377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13491_ _13491_/A _07648_/X vssd1 vssd1 vccd1 vccd1 _14035_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12442_ _12443_/CLK _12442_/D vssd1 vssd1 vccd1 vccd1 _12442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12175__B _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12373_ _12555_/CLK _12373_/D vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfxtp_2
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14112_ _14112_/A _08243_/X vssd1 vssd1 vccd1 vccd1 _14112_/Z sky130_fd_sc_hd__ebufn_8
X_11324_ _10548_/X _11312_/X _11323_/X _11319_/X vssd1 vssd1 vccd1 vccd1 _12758_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14043_ _14043_/A _07895_/X vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__ebufn_8
X_11255_ _11255_/A _11255_/B vssd1 vssd1 vccd1 vccd1 _11256_/A sky130_fd_sc_hd__and2_1
XANTENNA__09484__B _09484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10206_ _10206_/A vssd1 vssd1 vccd1 vccd1 _12478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ _11199_/B vssd1 vssd1 vccd1 vccd1 _11197_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__10423__B _10423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10137_ _10148_/C _10137_/B _10137_/C _10137_/D vssd1 vssd1 vccd1 vccd1 _10142_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10068_ _10086_/B _10076_/D vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__or2_1
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11535__A _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13827_ _13827_/A _06759_/X vssd1 vssd1 vccd1 vccd1 _13987_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_51_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13750__A _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13758_ _13758_/A _06947_/X vssd1 vssd1 vccd1 vccd1 _14078_/Z sky130_fd_sc_hd__ebufn_8
X_12709_ _12724_/CLK _12709_/D vssd1 vssd1 vccd1 vccd1 _12709_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11830__A0 peripheralBus_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13689_ _13689_/A _07122_/X vssd1 vssd1 vccd1 vccd1 _14105_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__06364__A _11457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08685__S0 _08549_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ _09937_/A vssd1 vssd1 vccd1 vccd1 _09934_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__08437__S0 _08417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09851_ _12375_/Q _09851_/B vssd1 vssd1 vccd1 vccd1 _09851_/X sky130_fd_sc_hd__and2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _10864_/C _12622_/Q _12623_/Q _12624_/Q _08733_/X _08735_/X vssd1 vssd1 vccd1
+ vccd1 _08802_/X sky130_fd_sc_hd__mux4_2
XFILLER_86_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09186_/X _09776_/X _09780_/X _09781_/X vssd1 vssd1 vccd1 vccd1 _12369_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06994_ _06994_/A vssd1 vssd1 vccd1 vccd1 _06994_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _08886_/A vssd1 vssd1 vccd1 vccd1 _08733_/X sky130_fd_sc_hd__buf_4
XANTENNA__07923__A _07923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _08606_/X _08612_/X _08610_/X _08614_/X _08663_/X _08652_/X vssd1 vssd1 vccd1
+ vccd1 _08664_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07615_ _07615_/A vssd1 vssd1 vccd1 vccd1 _07626_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _12450_/Q _12451_/Q _10101_/A _12453_/Q _08556_/X _08557_/X vssd1 vssd1 vccd1
+ vccd1 _08595_/X sky130_fd_sc_hd__mux4_2
XFILLER_42_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07546_ _07546_/A vssd1 vssd1 vccd1 vccd1 _07546_/X sky130_fd_sc_hd__clkbuf_1
X_07477_ _07477_/A vssd1 vssd1 vccd1 vccd1 _07477_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11180__A _11195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09216_ _09269_/A _09315_/D _09318_/A vssd1 vssd1 vccd1 vccd1 _09224_/C sky130_fd_sc_hd__and3_1
X_06428_ _06428_/A _06437_/B vssd1 vssd1 vccd1 vccd1 _06429_/A sky130_fd_sc_hd__or2_1
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09147_ input27/X vssd1 vssd1 vccd1 vccd1 _11490_/A sky130_fd_sc_hd__buf_6
X_06359_ _06359_/A _06362_/B _06362_/C vssd1 vssd1 vccd1 vccd1 _06360_/A sky130_fd_sc_hd__or3_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09585__A _11443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09078_ _09073_/X _09077_/X _09089_/S vssd1 vssd1 vccd1 vccd1 _10941_/B sky130_fd_sc_hd__mux2_2
XFILLER_150_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08029_ _08029_/A vssd1 vssd1 vccd1 vccd1 _08029_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11040_ _10652_/X _11027_/X _11038_/X _11039_/X vssd1 vssd1 vccd1 vccd1 _12682_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11942_ _11942_/A vssd1 vssd1 vccd1 vccd1 _12908_/D sky130_fd_sc_hd__clkbuf_1
X_13357__513 vssd1 vssd1 vccd1 vccd1 _13357__513/HI _14126_/A sky130_fd_sc_hd__conb_1
XFILLER_33_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11873_ _11886_/A _11873_/B vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__and2_1
XFILLER_60_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13570__A _13570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13612_ _13612_/A _07332_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824_ _10869_/D _10833_/A _10781_/X vssd1 vssd1 vccd1 vccd1 _10825_/B sky130_fd_sc_hd__o21ai_1
XFILLER_32_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11812__A0 _09631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13543_ _13543_/A _07509_/X vssd1 vssd1 vccd1 vccd1 _14087_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_158_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ _10774_/B _10755_/B vssd1 vssd1 vccd1 vccd1 _12617_/D sky130_fd_sc_hd__nor2_1
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13474_ _13474_/A _07690_/X vssd1 vssd1 vccd1 vccd1 _13666_/Z sky130_fd_sc_hd__ebufn_8
X_10686_ _13726_/A _10686_/B vssd1 vssd1 vccd1 vccd1 _10686_/X sky130_fd_sc_hd__or2_1
X_12425_ _12659_/CLK _12425_/D vssd1 vssd1 vccd1 vccd1 _12425_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11040__A1 _10652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09495__A _12134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12356_ _12356_/CLK _12356_/D vssd1 vssd1 vccd1 vccd1 _12356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11307_ _10662_/X _11299_/X _11305_/X _11306_/X vssd1 vssd1 vccd1 vccd1 _12751_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08419__S0 _08417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ _12289_/CLK _12287_/D vssd1 vssd1 vccd1 vccd1 _12287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14026_ _14026_/A _08082_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
X_11238_ _13881_/A _12737_/Q _11248_/S vssd1 vssd1 vccd1 vccd1 _11239_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13745__A _13745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11169_ _10652_/X _11155_/X _11168_/X _11166_/X vssd1 vssd1 vccd1 vccd1 _12715_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11500__C1 _11497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07400_ _07400_/A vssd1 vssd1 vccd1 vccd1 _07400_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08380_ _13393_/A vssd1 vssd1 vccd1 vccd1 _08380_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07331_ _07342_/A _07336_/B _07739_/C vssd1 vssd1 vccd1 vccd1 _07332_/A sky130_fd_sc_hd__or3_1
XFILLER_149_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10609__A _10952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07262_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07273_/C sky130_fd_sc_hd__clkbuf_1
X_13150__306 vssd1 vssd1 vccd1 vccd1 _13150__306/HI _13707_/A sky130_fd_sc_hd__conb_1
X_09001_ _12832_/Q vssd1 vssd1 vccd1 vccd1 _11640_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07193_ _07193_/A _07203_/B _07200_/C vssd1 vssd1 vccd1 vccd1 _07194_/A sky130_fd_sc_hd__or3_1
XANTENNA__11031__A1 _10377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09527__A2 _09513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09903_ _09915_/B vssd1 vssd1 vccd1 vccd1 _09913_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_116_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09834_ _09834_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _09835_/A sky130_fd_sc_hd__and2_1
XANTENNA__09852__B _13564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044__200 vssd1 vssd1 vccd1 vccd1 _13044__200/HI _13503_/A sky130_fd_sc_hd__conb_1
XFILLER_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09765_ _09878_/A vssd1 vssd1 vccd1 vccd1 _09765_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06977_ _07417_/A _06977_/B vssd1 vssd1 vccd1 vccd1 _06978_/A sky130_fd_sc_hd__or2_1
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08716_ _08595_/X _08659_/X _08685_/X _08715_/X _08694_/X _08634_/X vssd1 vssd1 vccd1
+ vccd1 _08716_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09696_ _09705_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09697_/A sky130_fd_sc_hd__and2_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06269__A _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10510__C _11410_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08647_ _13587_/A vssd1 vssd1 vccd1 vccd1 _08647_/X sky130_fd_sc_hd__clkbuf_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _13584_/A vssd1 vssd1 vccd1 vccd1 _08578_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _07531_/A _07531_/B _07538_/C vssd1 vssd1 vccd1 vccd1 _07530_/A sky130_fd_sc_hd__or3_1
X_10540_ _13689_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10540_/X sky130_fd_sc_hd__or2_1
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10238__B _13751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ _10477_/A _10471_/B vssd1 vssd1 vccd1 vccd1 _10472_/A sky130_fd_sc_hd__and2_1
X_12210_ _12968_/CLK _12210_/D vssd1 vssd1 vccd1 vccd1 _14107_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08569__A3 _08568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12141_ _12141_/A vssd1 vssd1 vccd1 vccd1 _12963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06451__B _07845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12072_ _10648_/A _12061_/X _12070_/X _12071_/X vssd1 vssd1 vccd1 vccd1 _12940_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11023_ _10999_/X _11000_/Y _11006_/X _11022_/X vssd1 vssd1 vccd1 vccd1 _11023_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__13565__A _13565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12974_ _12974_/CLK _12974_/D vssd1 vssd1 vccd1 vccd1 _14099_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11925_ _11977_/S vssd1 vssd1 vccd1 vccd1 _11940_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11856_ _11869_/A _11856_/B vssd1 vssd1 vccd1 vccd1 _11857_/A sky130_fd_sc_hd__and2_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06907__A _08168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10807_ _10863_/A _10863_/B _10865_/A _10865_/B vssd1 vssd1 vccd1 vccd1 _10809_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_13_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11787_ _11787_/A _11787_/B vssd1 vssd1 vccd1 vccd1 _11787_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__10429__A _10480_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08888__S0 _10697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13526_ _13526_/A _07555_/X vssd1 vssd1 vccd1 vccd1 _14102_/Z sky130_fd_sc_hd__ebufn_8
X_10738_ _10768_/A vssd1 vssd1 vccd1 vccd1 _10820_/C sky130_fd_sc_hd__buf_2
XFILLER_158_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13457_ _13457_/A _07736_/X vssd1 vssd1 vccd1 vccd1 _14033_/Z sky130_fd_sc_hd__ebufn_8
X_10669_ _10665_/X _10655_/X _10666_/X _10668_/X vssd1 vssd1 vccd1 vccd1 _12592_/D
+ sky130_fd_sc_hd__o211a_1
X_12408_ _12418_/CLK _12408_/D vssd1 vssd1 vccd1 vccd1 _13584_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_127_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13388_ _13388_/A _08346_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[29] sky130_fd_sc_hd__ebufn_8
XFILLER_126_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06642__A _06729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12339_ _12340_/CLK _12339_/D vssd1 vssd1 vccd1 vccd1 _13469_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_142_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14009_ _14009_/A _08134_/X vssd1 vssd1 vccd1 vccd1 _14009_/Z sky130_fd_sc_hd__ebufn_8
X_06900_ _06900_/A vssd1 vssd1 vccd1 vccd1 _07336_/B sky130_fd_sc_hd__buf_2
X_07880_ _07920_/A vssd1 vssd1 vccd1 vccd1 _07890_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_95_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07473__A _07473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06831_ _06831_/A vssd1 vssd1 vccd1 vccd1 _06831_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10611__B _13752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09550_ _09563_/A _09550_/B vssd1 vssd1 vccd1 vccd1 _09551_/A sky130_fd_sc_hd__and2_1
X_06762_ _06803_/A vssd1 vssd1 vccd1 vccd1 _06775_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08501_ _12265_/Q vssd1 vssd1 vccd1 vccd1 _09362_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09481_ _10250_/A vssd1 vssd1 vccd1 vccd1 _10637_/B sky130_fd_sc_hd__clkbuf_4
X_06693_ _06693_/A vssd1 vssd1 vccd1 vccd1 _06693_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ _08427_/X _08428_/X _08430_/X _08431_/X _08382_/X _08424_/X vssd1 vssd1 vccd1
+ vccd1 _08432_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11723__A _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08363_ _08363_/A vssd1 vssd1 vccd1 vccd1 _08363_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11788__C1 _09404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07314_ _07490_/A _07317_/B _07314_/C vssd1 vssd1 vccd1 vccd1 _07315_/A sky130_fd_sc_hd__or3_1
X_08294_ _08294_/A vssd1 vssd1 vccd1 vccd1 _08294_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07245_ _07245_/A vssd1 vssd1 vccd1 vccd1 _07245_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09847__B _13560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07176_ _07230_/A vssd1 vssd1 vccd1 vccd1 _07187_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_117_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06552__A _06729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09817_ _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09818_/A sky130_fd_sc_hd__and2_1
XFILLER_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08198__B _08208_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09748_ _09878_/A vssd1 vssd1 vccd1 vccd1 _09748_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _13493_/A _12347_/Q _09685_/S vssd1 vssd1 vccd1 vccd1 _09680_/B sky130_fd_sc_hd__mux2_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11710_ _12103_/B vssd1 vssd1 vccd1 vccd1 _11711_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10294__A2 _10278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12710_/CLK _12690_/D vssd1 vssd1 vccd1 vccd1 _13819_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06727__A _11028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11641_/A _11641_/B _11641_/C _11641_/D vssd1 vssd1 vccd1 vccd1 _11642_/D
+ sky130_fd_sc_hd__and4_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10249__A _10278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11572_ _11628_/A _11572_/B _11572_/C _11572_/D vssd1 vssd1 vccd1 vccd1 _11649_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 peripheralBus_address[4] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_2
X_10523_ _10650_/A vssd1 vssd1 vccd1 vccd1 _10523_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10454_ _10461_/A _10454_/B vssd1 vssd1 vccd1 vccd1 _10455_/A sky130_fd_sc_hd__and2_1
XFILLER_108_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06462__A _06462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10385_ _11160_/A vssd1 vssd1 vccd1 vccd1 _10385_/X sky130_fd_sc_hd__buf_6
XANTENNA__10754__B1 _10749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09773__A _10670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ _12124_/A vssd1 vssd1 vccd1 vccd1 _12958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12055_ _12055_/A _12055_/B _12055_/C _12055_/D vssd1 vssd1 vccd1 vccd1 _12056_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater108_A _14096_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__B1 _13760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11006_ _11001_/X _11002_/Y _11003_/X _11004_/Y _11005_/X vssd1 vssd1 vccd1 vccd1
+ _11006_/X sky130_fd_sc_hd__a221o_1
XFILLER_77_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output37_A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12957_ _12962_/CLK _12957_/D vssd1 vssd1 vccd1 vccd1 _12957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11908_ _12897_/Q _13369_/A vssd1 vssd1 vccd1 vccd1 _11910_/C sky130_fd_sc_hd__xor2_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12904_/CLK _12888_/D vssd1 vssd1 vccd1 vccd1 _12888_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11262__B _13946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11839_ _11839_/A vssd1 vssd1 vccd1 vccd1 _12884_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09948__A _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13509_ _13509_/A _07597_/X vssd1 vssd1 vccd1 vccd1 _13765_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_9_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07030_ _07030_/A vssd1 vssd1 vccd1 vccd1 _07030_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07468__A _07468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08981_ _08975_/X _08976_/X _08978_/X _08980_/X _08924_/X _08925_/X vssd1 vssd1 vccd1
+ vccd1 _08981_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13262__418 vssd1 vssd1 vccd1 vccd1 _13262__418/HI _13933_/A sky130_fd_sc_hd__conb_1
XFILLER_130_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07932_ _07932_/A vssd1 vssd1 vccd1 vccd1 _07932_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07863_ _08180_/A _07863_/B _08349_/B vssd1 vssd1 vccd1 vccd1 _07864_/A sky130_fd_sc_hd__or3_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09602_ _09602_/A _09602_/B _09602_/C _09602_/D vssd1 vssd1 vccd1 vccd1 _09608_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06814_ _11789_/B _07824_/C _11789_/A vssd1 vssd1 vccd1 vccd1 _06983_/B sky130_fd_sc_hd__or3b_4
X_13303__459 vssd1 vssd1 vccd1 vccd1 _13303__459/HI _14024_/A sky130_fd_sc_hd__conb_1
XFILLER_110_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11156__C _11156_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07794_ _09484_/A vssd1 vssd1 vccd1 vccd1 _08064_/A sky130_fd_sc_hd__buf_4
X_09533_ _09546_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _09534_/A sky130_fd_sc_hd__and2_1
XFILLER_71_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06745_ _06745_/A vssd1 vssd1 vccd1 vccd1 _06745_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09464_ _12287_/Q _13563_/A vssd1 vssd1 vccd1 vccd1 _09467_/B sky130_fd_sc_hd__xnor2_1
X_06676_ _06686_/A _06678_/B _06678_/C vssd1 vssd1 vccd1 vccd1 _06677_/A sky130_fd_sc_hd__or3_1
XANTENNA__06547__A _06547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13156__312 vssd1 vssd1 vccd1 vccd1 _13156__312/HI _13729_/A sky130_fd_sc_hd__conb_1
X_08415_ _11706_/B vssd1 vssd1 vccd1 vccd1 _13360_/A sky130_fd_sc_hd__buf_4
X_09395_ _09846_/A vssd1 vssd1 vccd1 vccd1 _09404_/A sky130_fd_sc_hd__buf_2
XFILLER_52_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08346_ _08346_/A vssd1 vssd1 vccd1 vccd1 _08346_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08277_ _08277_/A vssd1 vssd1 vccd1 vccd1 _08277_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07228_ _07239_/A _07231_/B _07228_/C vssd1 vssd1 vccd1 vccd1 _07229_/A sky130_fd_sc_hd__or3_1
XFILLER_164_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06282__A _07603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07159_ _07159_/A vssd1 vssd1 vccd1 vccd1 _07159_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10170_ _10173_/A _10170_/B vssd1 vssd1 vccd1 vccd1 _10171_/A sky130_fd_sc_hd__and2_1
XFILLER_121_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09354__B1 _09248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10251__B _11412_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13860_ _13860_/A _06670_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[21] sky130_fd_sc_hd__ebufn_8
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12811_ _12811_/CLK _12811_/D vssd1 vssd1 vccd1 vccd1 _12811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13791_ _13791_/A _06862_/X vssd1 vssd1 vccd1 vccd1 _13983_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11363__A _11363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12758_/CLK _12742_/D vssd1 vssd1 vccd1 vccd1 _12742_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06457__A _08210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12673_ _12699_/CLK _12673_/D vssd1 vssd1 vccd1 vccd1 _12673_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11624_ _11624_/A vssd1 vssd1 vccd1 vccd1 _12835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09768__A _13494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11555_ _11627_/A _11558_/C vssd1 vssd1 vccd1 vccd1 _11556_/C sky130_fd_sc_hd__nand2_1
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10506_ _10483_/Y _10489_/X _10505_/Y _13760_/A vssd1 vssd1 vccd1 vccd1 _10507_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11486_ _14103_/Z _13975_/A _11489_/S vssd1 vssd1 vccd1 vccd1 _11487_/B sky130_fd_sc_hd__mux2_1
X_10437_ _10444_/A _10437_/B vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__and2_1
XFILLER_124_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _12509_/Q _13751_/A vssd1 vssd1 vccd1 vccd1 _10372_/A sky130_fd_sc_hd__xor2_1
XFILLER_124_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12107_/A vssd1 vssd1 vccd1 vccd1 _12953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10442__A _10480_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10299_ _10299_/A vssd1 vssd1 vccd1 vccd1 _12501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12038_ _12933_/Q _13372_/A vssd1 vssd1 vccd1 vccd1 _12040_/C sky130_fd_sc_hd__xor2_1
XANTENNA__11257__B _13944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13753__A _13753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13989_ _13989_/A _06317_/X vssd1 vssd1 vccd1 vccd1 _14117_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_19_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06530_ _06534_/A _06540_/B _06540_/C vssd1 vssd1 vccd1 vccd1 _06531_/A sky130_fd_sc_hd__or3_1
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06461_ _06461_/A vssd1 vssd1 vccd1 vccd1 _06461_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08200_ _08240_/A vssd1 vssd1 vccd1 vccd1 _08212_/A sky130_fd_sc_hd__clkbuf_1
X_09180_ _10670_/A _09145_/A _09179_/X _09939_/A vssd1 vssd1 vccd1 vccd1 _12223_/D
+ sky130_fd_sc_hd__a211o_1
X_06392_ _06392_/A vssd1 vssd1 vccd1 vccd1 _06392_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08131_ _08135_/A _08189_/B _08131_/C vssd1 vssd1 vccd1 vccd1 _08132_/A sky130_fd_sc_hd__or3_4
XFILLER_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08062_ _08065_/A _08062_/B _08070_/C vssd1 vssd1 vccd1 vccd1 _08063_/A sky130_fd_sc_hd__or3_1
X_07013_ _07019_/A _07019_/B vssd1 vssd1 vccd1 vccd1 _07014_/A sky130_fd_sc_hd__or2_1
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08482__S1 _08374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ _10939_/B vssd1 vssd1 vccd1 vccd1 _11388_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07915_ _07921_/A _07917_/B _07917_/C vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__or3_1
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08895_ _08774_/X _08840_/X _08866_/X _08894_/X _08810_/X _08812_/X vssd1 vssd1 vccd1
+ vccd1 _08895_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09887__A1 _09756_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09860__B _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _07846_/A vssd1 vssd1 vccd1 vccd1 _07846_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07777_ _07782_/A _07779_/B _07787_/C vssd1 vssd1 vccd1 vccd1 _07778_/A sky130_fd_sc_hd__or3_1
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09516_ _13433_/A _09513_/X _09515_/X _09509_/X vssd1 vssd1 vccd1 vccd1 _12302_/D
+ sky130_fd_sc_hd__o211a_1
X_06728_ _08195_/B vssd1 vssd1 vccd1 vccd1 _06738_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09447_ _09447_/A vssd1 vssd1 vccd1 vccd1 _12287_/D sky130_fd_sc_hd__clkbuf_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06659_ _06659_/A _06664_/B _06664_/C vssd1 vssd1 vccd1 vccd1 _06660_/A sky130_fd_sc_hd__or3_1
XFILLER_25_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09378_ _09382_/B _09382_/C vssd1 vssd1 vccd1 vccd1 _09379_/B sky130_fd_sc_hd__and2_1
XFILLER_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ _08336_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08330_/A sky130_fd_sc_hd__or2_1
XFILLER_149_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11340_ _11344_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11341_/A sky130_fd_sc_hd__and2_1
XFILLER_137_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11271_ _12739_/Q _13947_/A vssd1 vssd1 vccd1 vccd1 _11273_/C sky130_fd_sc_hd__xor2_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10222_ _10222_/A vssd1 vssd1 vccd1 vccd1 _12483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13284__440 vssd1 vssd1 vccd1 vccd1 _13284__440/HI _13989_/A sky130_fd_sc_hd__conb_1
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10153_ _10155_/B _10155_/C vssd1 vssd1 vccd1 vccd1 _10153_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10084_ _10146_/A _10084_/B _10084_/C vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__and3_1
X_13325__481 vssd1 vssd1 vccd1 vccd1 _13325__481/HI _14062_/A sky130_fd_sc_hd__conb_1
XFILLER_75_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13912_ _13912_/A _06522_/X vssd1 vssd1 vccd1 vccd1 _13976_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_63_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13843_ _13843_/A _06715_/X vssd1 vssd1 vccd1 vccd1 _14067_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11437__A1 _10670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10986_ _10986_/A _10986_/B vssd1 vssd1 vccd1 vccd1 _10987_/A sky130_fd_sc_hd__and2_1
X_13774_ _13774_/A _06908_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
X_12725_ _12743_/CLK _12725_/D vssd1 vssd1 vccd1 vccd1 _13853_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09498__A _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11821__A _11834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12656_ _12656_/CLK _12656_/D vssd1 vssd1 vccd1 vccd1 _12656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ _11640_/C _11610_/C vssd1 vssd1 vccd1 vccd1 _11609_/A sky130_fd_sc_hd__and2_1
XFILLER_128_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12587_ _12589_/CLK _12587_/D vssd1 vssd1 vccd1 vccd1 _13714_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11538_ _11571_/D vssd1 vssd1 vccd1 vccd1 _11627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13748__A _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11469_ _11481_/A _11469_/B vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__or2_1
XFILLER_99_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09961__A _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07700_ _07700_/A vssd1 vssd1 vccd1 vccd1 _07700_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08680_ _12457_/Q _12458_/Q _10130_/A _12460_/Q _08629_/X _08630_/X vssd1 vssd1 vccd1
+ vccd1 _08680_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08541__A1 _08452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07631_ _07631_/A vssd1 vssd1 vccd1 vccd1 _07631_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11428__A1 _11170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ _07575_/A _08103_/B _07564_/C vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__or3_1
XFILLER_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09301_ _09329_/B _09299_/A _09236_/X vssd1 vssd1 vccd1 vccd1 _09302_/B sky130_fd_sc_hd__o21ai_1
X_06513_ _06513_/A vssd1 vssd1 vccd1 vccd1 _06513_/X sky130_fd_sc_hd__clkbuf_1
X_07493_ _07507_/A vssd1 vssd1 vccd1 vccd1 _07504_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_110_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09232_ _09317_/D _09235_/C vssd1 vssd1 vccd1 vccd1 _09234_/A sky130_fd_sc_hd__and2_1
X_06444_ _06444_/A vssd1 vssd1 vccd1 vccd1 _06444_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09201__A _09269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ _09160_/X _09130_/X _09162_/X _09141_/X vssd1 vssd1 vccd1 vccd1 _12219_/D
+ sky130_fd_sc_hd__o211a_1
X_06375_ _07861_/A vssd1 vssd1 vccd1 vccd1 _06391_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08114_ _08114_/A vssd1 vssd1 vccd1 vccd1 _08114_/X sky130_fd_sc_hd__clkbuf_1
X_09094_ _11924_/B vssd1 vssd1 vccd1 vccd1 _10250_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13268__424 vssd1 vssd1 vccd1 vccd1 _13268__424/HI _13959_/A sky130_fd_sc_hd__conb_1
X_08045_ _08045_/A vssd1 vssd1 vccd1 vccd1 _08045_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09855__B _13557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08455__S1 _08374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13309__465 vssd1 vssd1 vccd1 vccd1 _13309__465/HI _14030_/A sky130_fd_sc_hd__conb_1
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09996_ _09996_/A _09996_/B vssd1 vssd1 vccd1 vccd1 _12427_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09871__A _11151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08947_ _09068_/A vssd1 vssd1 vccd1 vccd1 _08947_/X sky130_fd_sc_hd__buf_2
X_12982__138 vssd1 vssd1 vccd1 vccd1 _12982__138/HI _13379_/A sky130_fd_sc_hd__conb_1
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13393__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__B _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__A _10872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08878_ _12654_/Q vssd1 vssd1 vccd1 vccd1 _10921_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07829_ _07964_/A vssd1 vssd1 vccd1 vccd1 _07843_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07822__C _07822_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10840_ _10876_/C _10869_/B _10840_/C _10877_/A vssd1 vssd1 vccd1 vccd1 _10848_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_60_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_99_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ _10771_/A vssd1 vssd1 vccd1 vccd1 _12621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ _12517_/CLK _12510_/D vssd1 vssd1 vccd1 vccd1 _12510_/Q sky130_fd_sc_hd__dfxtp_1
X_13490_ _13490_/A _07650_/X vssd1 vssd1 vccd1 vccd1 _14034_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_13_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12441_ _12443_/CLK _12441_/D vssd1 vssd1 vccd1 vccd1 _12441_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09111__A _13628_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_22_clk_A _12881_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12372_ _12404_/CLK _12372_/D vssd1 vssd1 vccd1 vccd1 _13501_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11323_ _13885_/A _11323_/B vssd1 vssd1 vccd1 vccd1 _11323_/X sky130_fd_sc_hd__or2_1
X_14111_ _14111_/A _08239_/X vssd1 vssd1 vccd1 vccd1 _14111_/Z sky130_fd_sc_hd__ebufn_8
Xclkbuf_4_0_0_clk clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_clk/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13568__A _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07566__A _09484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ _13886_/A _12742_/Q _11254_/S vssd1 vssd1 vccd1 vccd1 _11255_/B sky130_fd_sc_hd__mux2_1
X_14042_ _14042_/A _07891_/X vssd1 vssd1 vccd1 vccd1 _14106_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__06470__A _06481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09484__C _12062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10205_ _10208_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__and2_1
XFILLER_134_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11185_ _11185_/A vssd1 vssd1 vccd1 vccd1 _11185_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10136_ _10136_/A vssd1 vssd1 vccd1 vccd1 _12460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061__217 vssd1 vssd1 vccd1 vccd1 _13061__217/HI _13536_/A sky130_fd_sc_hd__conb_1
X_10067_ _10098_/B vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08397__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13826_ _13826_/A _06761_/X vssd1 vssd1 vccd1 vccd1 _14082_/Z sky130_fd_sc_hd__ebufn_8
X_13102__258 vssd1 vssd1 vccd1 vccd1 _13102__258/HI _13611_/A sky130_fd_sc_hd__conb_1
XFILLER_90_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13757_ _13757_/A _06949_/X vssd1 vssd1 vccd1 vccd1 _14077_/Z sky130_fd_sc_hd__ebufn_8
X_10969_ _10969_/A _10969_/B vssd1 vssd1 vccd1 vccd1 _10970_/A sky130_fd_sc_hd__and2_1
X_12708_ _12743_/CLK _12708_/D vssd1 vssd1 vccd1 vccd1 _12708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13688_ _13688_/A _07125_/X vssd1 vssd1 vccd1 vccd1 _14072_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11270__B _13950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ _12820_/CLK _12639_/D vssd1 vssd1 vccd1 vccd1 _12639_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10167__A _13788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09956__A _13593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08685__S1 _08551_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06380__A _08338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08437__S1 _08418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10614__B _10614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09850_ _12375_/Q _13552_/A vssd1 vssd1 vccd1 vccd1 _09850_/Y sky130_fd_sc_hd__nor2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__A _09711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ _12621_/Q vssd1 vssd1 vccd1 vccd1 _10864_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _06995_/A _06995_/B vssd1 vssd1 vccd1 vccd1 _06994_/A sky130_fd_sc_hd__or2_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _09878_/A vssd1 vssd1 vccd1 vccd1 _09781_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _13776_/A vssd1 vssd1 vccd1 vccd1 _08886_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09711__A0 hold2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08663_ _13587_/A vssd1 vssd1 vccd1 vccd1 _08663_/X sky130_fd_sc_hd__buf_2
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13941__A _13941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07614_ _07614_/A vssd1 vssd1 vccd1 vccd1 _07614_/X sky130_fd_sc_hd__clkbuf_1
X_08594_ _12452_/Q vssd1 vssd1 vccd1 vccd1 _10101_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07545_ _07545_/A _07545_/B _07551_/C vssd1 vssd1 vccd1 vccd1 _07546_/A sky130_fd_sc_hd__or3_1
XANTENNA__12074__A1 _10652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ _07478_/A _07484_/B vssd1 vssd1 vccd1 vccd1 _07477_/A sky130_fd_sc_hd__or2_1
X_06427_ _06913_/A vssd1 vssd1 vccd1 vccd1 _06437_/B sky130_fd_sc_hd__clkbuf_1
X_09215_ _09215_/A vssd1 vssd1 vccd1 vccd1 _12231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06274__B _09097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ _09146_/A _09152_/B vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__and2_1
X_06358_ _06358_/A vssd1 vssd1 vccd1 vccd1 _06358_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09077_ _08960_/X _09020_/X _09046_/X _09076_/X _09056_/X _09057_/X vssd1 vssd1 vccd1
+ vccd1 _09077_/X sky130_fd_sc_hd__mux4_1
X_06289_ _06289_/A vssd1 vssd1 vccd1 vccd1 _06289_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08028_ _08039_/A _08033_/B _08030_/C vssd1 vssd1 vccd1 vccd1 _08029_/A sky130_fd_sc_hd__or3_1
XFILLER_135_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06290__A _08364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09950__A0 _13623_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09979_ _09981_/B _09972_/X _09978_/X vssd1 vssd1 vccd1 vccd1 _09979_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07833__B _07840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09106__A _11503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ _11945_/A _11941_/B vssd1 vssd1 vccd1 vccd1 _11942_/A sky130_fd_sc_hd__and2_1
XFILLER_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11872_ _12894_/Q _14038_/A _11878_/S vssd1 vssd1 vccd1 vccd1 _11873_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ _13611_/A _07334_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
X_10823_ _10869_/D _10833_/A vssd1 vssd1 vccd1 vccd1 _10825_/A sky130_fd_sc_hd__and2_1
XANTENNA__12065__A1 _11153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_118_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _12264_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13542_ _13542_/A _07511_/X vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_8
X_10754_ _10806_/A _10760_/D _10749_/X vssd1 vssd1 vccd1 vccd1 _10755_/B sky130_fd_sc_hd__o21ai_1
XFILLER_158_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13473_ _13473_/A _07692_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
X_10685_ _10548_/X _10673_/X _10684_/X _10682_/X vssd1 vssd1 vccd1 vccd1 _12598_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09776__A _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ _12659_/CLK _12424_/D vssd1 vssd1 vccd1 vccd1 _12424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12355_ _12377_/CLK _12355_/D vssd1 vssd1 vccd1 vccd1 _12355_/Q sky130_fd_sc_hd__dfxtp_1
X_11306_ _11430_/A vssd1 vssd1 vccd1 vccd1 _11306_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12286_ _12290_/CLK _12286_/D vssd1 vssd1 vccd1 vccd1 _12286_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08419__S1 _08418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11237_ _11237_/A vssd1 vssd1 vccd1 vccd1 _12736_/D sky130_fd_sc_hd__clkbuf_1
X_14025_ _14025_/A _08078_/X vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_141_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11168_ _13843_/A _11168_/B vssd1 vssd1 vccd1 vccd1 _11168_/X sky130_fd_sc_hd__or2_1
XANTENNA__10551__A1 _10548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ _10126_/C _10114_/X _10123_/A vssd1 vssd1 vccd1 vccd1 _10119_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_121_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11099_ _11112_/A _11099_/B vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__and2_1
XFILLER_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11265__B _13949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13761__A _13761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13809_ _13809_/A _06807_/X vssd1 vssd1 vccd1 vccd1 _14065_/Z sky130_fd_sc_hd__ebufn_8
Xclkbuf_leaf_109_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _12320_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11281__A _11408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07330_ _07371_/A vssd1 vssd1 vccd1 vccd1 _07342_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06375__A _07861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07261_ _07261_/A vssd1 vssd1 vccd1 vccd1 _07261_/X sky130_fd_sc_hd__clkbuf_1
X_09000_ _12830_/Q vssd1 vssd1 vccd1 vccd1 _11641_/C sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk/X sky130_fd_sc_hd__clkbuf_2
X_07192_ _07205_/A vssd1 vssd1 vccd1 vccd1 _07203_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08432__A0 _08427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13230__386 vssd1 vssd1 vccd1 vccd1 _13230__386/HI _13869_/A sky130_fd_sc_hd__conb_1
XFILLER_160_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09902_ _09902_/A vssd1 vssd1 vccd1 vccd1 _09902_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13936__A _13936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09833_ _13531_/A _12386_/Q _09837_/S vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__mux2_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11456__A _11634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09764_ _13493_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09764_/X sky130_fd_sc_hd__or2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06976_ _06976_/A vssd1 vssd1 vccd1 vccd1 _06976_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08715_ _10148_/B _12463_/Q _12464_/Q _12465_/Q _09929_/A _08709_/X vssd1 vssd1 vccd1
+ vccd1 _08715_/X sky130_fd_sc_hd__mux4_1
X_09695_ _13497_/A _12351_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09696_/B sky130_fd_sc_hd__mux2_1
XFILLER_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13124__280 vssd1 vssd1 vccd1 vccd1 _13124__280/HI _13665_/A sky130_fd_sc_hd__conb_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08646_ _10101_/A _10111_/C _10111_/B _10111_/A _08629_/X _08630_/X vssd1 vssd1 vccd1
+ vccd1 _08646_/X sky130_fd_sc_hd__mux4_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11903__B _13372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _12426_/Q _12427_/Q _09997_/A _12429_/Q _08575_/X _08576_/X vssd1 vssd1 vccd1
+ vccd1 _08577_/X sky130_fd_sc_hd__mux4_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10058__B1 _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09999__B1 _09994_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07528_ _07528_/A vssd1 vssd1 vccd1 vccd1 _07528_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06285__A _06547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07459_ _07466_/A _07459_/B vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__or2_1
XFILLER_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10470_ _13691_/A _12546_/Q _10473_/S vssd1 vssd1 vccd1 vccd1 _10471_/B sky130_fd_sc_hd__mux2_1
X_09129_ _09156_/A vssd1 vssd1 vccd1 vccd1 _09152_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14007__A _14007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ _12149_/A _12140_/B vssd1 vssd1 vccd1 vccd1 _12141_/A sky130_fd_sc_hd__and2_1
XFILLER_151_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12988__144 vssd1 vssd1 vccd1 vccd1 _12988__144/HI _13385_/A sky130_fd_sc_hd__conb_1
X_12071_ _12084_/A vssd1 vssd1 vccd1 vccd1 _12071_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ _11022_/A _11022_/B _11022_/C vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__or3_1
XFILLER_150_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12973_ _12980_/CLK _12973_/D vssd1 vssd1 vccd1 vccd1 _14098_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11924_ _11924_/A _11924_/B _11924_/C vssd1 vssd1 vccd1 vccd1 _11977_/S sky130_fd_sc_hd__or3_2
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _12889_/Q _14033_/A _11861_/S vssd1 vssd1 vccd1 vccd1 _11856_/B sky130_fd_sc_hd__mux2_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ _10806_/A _10806_/B _10806_/C _10806_/D vssd1 vssd1 vccd1 vccd1 _10866_/A
+ sky130_fd_sc_hd__and4_1
X_13173__329 vssd1 vssd1 vccd1 vccd1 _13173__329/HI _13766_/A sky130_fd_sc_hd__conb_1
XFILLER_158_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11786_ _11786_/A _11786_/B _11786_/C vssd1 vssd1 vccd1 vccd1 _11787_/B sky130_fd_sc_hd__or3_1
X_13525_ _13525_/A _07557_/X vssd1 vssd1 vccd1 vccd1 _14037_/Z sky130_fd_sc_hd__ebufn_8
X_10737_ _10915_/A _11503_/B _10737_/C vssd1 vssd1 vccd1 vccd1 _10768_/A sky130_fd_sc_hd__and3_1
XFILLER_158_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13456_ _13456_/A _07738_/X vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_8
X_10668_ _11039_/A vssd1 vssd1 vccd1 vccd1 _10668_/X sky130_fd_sc_hd__clkbuf_2
X_12407_ _12418_/CLK _12407_/D vssd1 vssd1 vccd1 vccd1 _13583_/A sky130_fd_sc_hd__dfxtp_4
X_10599_ _10602_/A _10599_/B vssd1 vssd1 vccd1 vccd1 _10600_/A sky130_fd_sc_hd__and2_1
X_13387_ _13387_/A _08344_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
XFILLER_127_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06642__B _07323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12338_ _12340_/CLK _12338_/D vssd1 vssd1 vccd1 vccd1 _13468_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13756__A _13756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13067__223 vssd1 vssd1 vccd1 vccd1 _13067__223/HI _13542_/A sky130_fd_sc_hd__conb_1
X_12269_ _12912_/CLK _12269_/D vssd1 vssd1 vccd1 vccd1 _12269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14008_ _14008_/A _08139_/X vssd1 vssd1 vccd1 vccd1 _14072_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10524__A1 _09756_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06830_ _06836_/A _06830_/B _07234_/C vssd1 vssd1 vccd1 vccd1 _06831_/A sky130_fd_sc_hd__or3_1
X_13108__264 vssd1 vssd1 vccd1 vccd1 _13108__264/HI _13633_/A sky130_fd_sc_hd__conb_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06761_ _06761_/A vssd1 vssd1 vccd1 vccd1 _06761_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09142__A1 _09139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ _08400_/X _08401_/X _08406_/X _08407_/X _08492_/X _08449_/X vssd1 vssd1 vccd1
+ vccd1 _08500_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09480_ _13570_/A _09479_/X _09414_/S _09192_/X vssd1 vssd1 vccd1 vccd1 _12291_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06692_ _06701_/A _06692_/B _06692_/C vssd1 vssd1 vccd1 vccd1 _06693_/A sky130_fd_sc_hd__or3_1
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08431_ _12258_/Q _12259_/Q _12260_/Q _12261_/Q _08404_/X _08405_/X vssd1 vssd1 vccd1
+ vccd1 _08431_/X sky130_fd_sc_hd__mux4_2
XANTENNA__06817__B _07323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ _08364_/A _08364_/B _08364_/C vssd1 vssd1 vccd1 vccd1 _08363_/A sky130_fd_sc_hd__or3_1
XFILLER_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07313_ _07313_/A vssd1 vssd1 vccd1 vccd1 _07313_/X sky130_fd_sc_hd__clkbuf_1
X_08293_ _08300_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08294_/A sky130_fd_sc_hd__or2_1
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07244_ _07253_/A _07250_/B _07246_/C vssd1 vssd1 vccd1 vccd1 _07245_/A sky130_fd_sc_hd__or3_1
XANTENNA__06833__A _06967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12881__CLK _12881_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12201__A1 _10662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07175_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07230_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06552__B _07323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10515__A1 _10377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11186__A _11199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09816_ _13526_/A _12381_/Q _09820_/S vssd1 vssd1 vccd1 vccd1 _09817_/B sky130_fd_sc_hd__mux2_1
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09747_ _13488_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09747_/X sky130_fd_sc_hd__or2_1
X_06959_ _06959_/A vssd1 vssd1 vccd1 vccd1 _06959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08567__S0 _08559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09678_ _09678_/A vssd1 vssd1 vccd1 vccd1 _12346_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08708_/A vssd1 vssd1 vccd1 vccd1 _08629_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A _11640_/B _11640_/C vssd1 vssd1 vccd1 vccd1 _11642_/C sky130_fd_sc_hd__and3_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ _11626_/A _11626_/B _11627_/C _11571_/D vssd1 vssd1 vccd1 vccd1 _11572_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_128_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07839__A _08335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10522_ _13683_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _10522_/X sky130_fd_sc_hd__or2_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10453_ _13686_/A _12541_/Q _10456_/S vssd1 vssd1 vccd1 vccd1 _10454_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10265__A _10293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10384_ _10377_/X _10379_/X _10382_/X _10383_/X vssd1 vssd1 vccd1 vccd1 _12518_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11951__A0 _09633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ _12132_/A _12123_/B vssd1 vssd1 vccd1 vccd1 _12124_/A sky130_fd_sc_hd__and2_1
XFILLER_151_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07574__A _07615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12054_ _12920_/Q _13359_/A vssd1 vssd1 vccd1 vccd1 _12055_/D sky130_fd_sc_hd__xor2_1
XFILLER_77_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11005_ _12672_/Q _13946_/A vssd1 vssd1 vccd1 vccd1 _11005_/X sky130_fd_sc_hd__xor2_1
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08558__S0 _08556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11824__A _11834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12956_ _12981_/CLK _12956_/D vssd1 vssd1 vccd1 vccd1 _12956_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06918__A _06955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11907_ _12893_/Q _13365_/A vssd1 vssd1 vccd1 vccd1 _11910_/B sky130_fd_sc_hd__xor2_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _12961_/CLK _12887_/D vssd1 vssd1 vccd1 vccd1 _12887_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06637__B _09096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11838_ _11852_/A _11838_/B vssd1 vssd1 vccd1 vccd1 _11839_/A sky130_fd_sc_hd__and2_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11769_ _12855_/Q _13360_/A vssd1 vssd1 vccd1 vccd1 _11770_/D sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_40_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _12938_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ _13508_/A _07599_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__06653__A _06680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13439_ _13439_/A _07780_/X vssd1 vssd1 vccd1 vccd1 _14111_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10175__A _10988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ _12837_/Q _11649_/A _12839_/Q _12840_/Q _08918_/X _08919_/X vssd1 vssd1 vccd1
+ vccd1 _08980_/X sky130_fd_sc_hd__mux4_2
XFILLER_102_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07484__A _08089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07931_ _07936_/A _07931_/B _07931_/C vssd1 vssd1 vccd1 vccd1 _07932_/A sky130_fd_sc_hd__or3_1
X_07862_ _07862_/A vssd1 vssd1 vccd1 vccd1 _07862_/X sky130_fd_sc_hd__clkbuf_1
X_09601_ _12315_/Q _13558_/A vssd1 vssd1 vccd1 vccd1 _09602_/D sky130_fd_sc_hd__xor2_1
X_13342__498 vssd1 vssd1 vccd1 vccd1 _13342__498/HI _14111_/A sky130_fd_sc_hd__conb_1
X_06813_ _09097_/A input6/X _09097_/B _09097_/C vssd1 vssd1 vccd1 vccd1 _07824_/C
+ sky130_fd_sc_hd__or4_1
X_07793_ _07793_/A vssd1 vssd1 vccd1 vccd1 _07793_/X sky130_fd_sc_hd__clkbuf_1
X_09532_ _13455_/A _12308_/Q _09610_/B vssd1 vssd1 vccd1 vccd1 _09533_/B sky130_fd_sc_hd__mux2_1
X_06744_ _06746_/A _06751_/B _06751_/C vssd1 vssd1 vccd1 vccd1 _06745_/A sky130_fd_sc_hd__or3_1
XFILLER_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09463_ _12281_/Q _13557_/A vssd1 vssd1 vccd1 vccd1 _09467_/A sky130_fd_sc_hd__xnor2_1
X_06675_ _06675_/A vssd1 vssd1 vccd1 vccd1 _06686_/A sky130_fd_sc_hd__buf_2
X_13195__351 vssd1 vssd1 vccd1 vccd1 _13195__351/HI _13802_/A sky130_fd_sc_hd__conb_1
X_08414_ _08402_/X _08413_/X _08498_/S vssd1 vssd1 vccd1 vccd1 _11706_/B sky130_fd_sc_hd__mux2_2
X_09394_ _09967_/B vssd1 vssd1 vccd1 vccd1 _09846_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08345_ _08347_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08346_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_31_clk _12759_/CLK vssd1 vssd1 vccd1 vccd1 _12786_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_165_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13236__392 vssd1 vssd1 vccd1 vccd1 _13236__392/HI _13891_/A sky130_fd_sc_hd__conb_1
X_08276_ _08276_/A _08276_/B _08276_/C vssd1 vssd1 vccd1 vccd1 _08277_/A sky130_fd_sc_hd__or3_1
XFILLER_138_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07227_ _07227_/A vssd1 vssd1 vccd1 vccd1 _07227_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09874__A _09902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07158_ _07166_/A _07163_/B _07160_/C vssd1 vssd1 vccd1 vccd1 _07159_/A sky130_fd_sc_hd__or3_1
XFILLER_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09593__B _13561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07089_ _07089_/A vssd1 vssd1 vccd1 vccd1 _07089_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_98_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _12367_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11697__C1 _11515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10251__C _10693_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12810_ _12811_/CLK _12810_/D vssd1 vssd1 vccd1 vccd1 _12810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13790_ _13790_/A _06864_/X vssd1 vssd1 vccd1 vccd1 _14078_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_15_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12758_/CLK _12741_/D vssd1 vssd1 vccd1 vccd1 _12741_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08865__A0 _08765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12687_/CLK _12672_/D vssd1 vssd1 vccd1 vccd1 _12672_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11703_/A _11623_/B _11623_/C vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__and3_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_clk _12881_/CLK vssd1 vssd1 vccd1 vccd1 _12873_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11554_ _11627_/A _11558_/C vssd1 vssd1 vccd1 vccd1 _11556_/B sky130_fd_sc_hd__or2_1
XANTENNA__09290__B1 _09392_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10505_ _10505_/A _10505_/B _10505_/C vssd1 vssd1 vccd1 vccd1 _10505_/Y sky130_fd_sc_hd__nor3_1
X_11485_ _11485_/A vssd1 vssd1 vccd1 vccd1 _12800_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10436_ _13681_/A _12536_/Q _10507_/B vssd1 vssd1 vccd1 vccd1 _10437_/B sky130_fd_sc_hd__mux2_1
XFILLER_164_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10727__A1 _10408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater120_A peripheralBus_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ _10367_/A _10367_/B _10367_/C _10367_/D vssd1 vssd1 vccd1 vccd1 _10373_/B
+ sky130_fd_sc_hd__or4_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _12115_/A _12106_/B vssd1 vssd1 vccd1 vccd1 _12107_/A sky130_fd_sc_hd__and2_1
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10298_/A _10298_/B vssd1 vssd1 vccd1 vccd1 _10299_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_89_clk _12438_/CLK vssd1 vssd1 vccd1 vccd1 _12461_/CLK sky130_fd_sc_hd__clkbuf_16
X_12037_ _12931_/Q _13370_/A vssd1 vssd1 vccd1 vccd1 _12040_/B sky130_fd_sc_hd__xor2_1
XFILLER_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13179__335 vssd1 vssd1 vccd1 vccd1 _13179__335/HI _13772_/A sky130_fd_sc_hd__conb_1
X_13988_ _13988_/A _06319_/X vssd1 vssd1 vccd1 vccd1 _13988_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_92_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12939_ _12946_/CLK _12939_/D vssd1 vssd1 vccd1 vccd1 _14065_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06367__B _07822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06460_ _07822_/B _07822_/C _06472_/C vssd1 vssd1 vccd1 vccd1 _06461_/A sky130_fd_sc_hd__or3_1
XFILLER_61_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06391_ _06391_/A _06400_/B vssd1 vssd1 vccd1 vccd1 _06392_/A sky130_fd_sc_hd__or2_1
XFILLER_159_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_clk _12217_/CLK vssd1 vssd1 vccd1 vccd1 _12968_/CLK sky130_fd_sc_hd__clkbuf_16
X_08130_ _11026_/B vssd1 vssd1 vccd1 vccd1 _08189_/B sky130_fd_sc_hd__clkbuf_2
X_08061_ _08061_/A vssd1 vssd1 vccd1 vccd1 _08061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ _07012_/A vssd1 vssd1 vccd1 vccd1 _07012_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11729__A _11763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08963_ _08954_/X _08961_/X _09071_/S vssd1 vssd1 vccd1 vccd1 _10939_/B sky130_fd_sc_hd__mux2_2
XANTENNA__08103__A _08110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__B _13754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13944__A _13944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07914_ _07914_/A vssd1 vssd1 vccd1 vccd1 _07914_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08894_ _10921_/B _10921_/A _12657_/Q _12658_/Q _10697_/A _08887_/X vssd1 vssd1 vccd1
+ vccd1 _08894_/X sky130_fd_sc_hd__mux4_2
XFILLER_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07845_ _07845_/A _07845_/B vssd1 vssd1 vccd1 vccd1 _07846_/A sky130_fd_sc_hd__or2_1
XFILLER_83_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11464__A _12084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07776_ _07817_/A vssd1 vssd1 vccd1 vccd1 _07787_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09515_ _11184_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09515_/X sky130_fd_sc_hd__or2_1
X_06727_ _11028_/B vssd1 vssd1 vccd1 vccd1 _08195_/B sky130_fd_sc_hd__clkbuf_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09455_/A _09446_/B vssd1 vssd1 vccd1 vccd1 _09447_/A sky130_fd_sc_hd__and2_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ _06658_/A vssd1 vssd1 vccd1 vccd1 _06658_/X sky130_fd_sc_hd__clkbuf_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11911__B _13361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09377_ _09377_/A _09377_/B _09377_/C vssd1 vssd1 vccd1 vccd1 _09382_/C sky130_fd_sc_hd__and3_1
XANTENNA__09588__B _13562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06589_ _06597_/A _06589_/B _06589_/C vssd1 vssd1 vccd1 vccd1 _06590_/A sky130_fd_sc_hd__or3_1
X_08328_ _08328_/A vssd1 vssd1 vccd1 vccd1 _08328_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06293__A _06442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08259_ _08264_/A _08261_/B _08264_/C vssd1 vssd1 vccd1 vccd1 _08260_/A sky130_fd_sc_hd__or3_1
XFILLER_4_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11270_ _12742_/Q _13950_/A vssd1 vssd1 vccd1 vccd1 _11273_/B sky130_fd_sc_hd__xor2_1
XFILLER_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13013__169 vssd1 vssd1 vccd1 vccd1 _13013__169/HI _13440_/A sky130_fd_sc_hd__conb_1
X_10221_ _10298_/A _10221_/B vssd1 vssd1 vccd1 vccd1 _10222_/A sky130_fd_sc_hd__and2_1
XFILLER_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10152_ _10152_/A vssd1 vssd1 vccd1 vccd1 _12464_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08013__A _08067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10083_ _10098_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10084_/C sky130_fd_sc_hd__nand2_1
XFILLER_59_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13911_ _13911_/A _06525_/X vssd1 vssd1 vccd1 vccd1 _14007_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13842_ _13842_/A _06718_/X vssd1 vssd1 vccd1 vccd1 _14066_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_28_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06468__A _06688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13773_ _13773_/A _06910_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
X_10985_ _13819_/A _12673_/Q _10990_/S vssd1 vssd1 vccd1 vccd1 _10986_/B sky130_fd_sc_hd__mux2_1
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12724_ _12724_/CLK _12724_/D vssd1 vssd1 vccd1 vccd1 _13852_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12655_ _12660_/CLK _12655_/D vssd1 vssd1 vccd1 vccd1 _12655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11606_ _12831_/Q vssd1 vssd1 vccd1 vccd1 _11640_/C sky130_fd_sc_hd__clkbuf_1
X_12586_ _12586_/CLK _12586_/D vssd1 vssd1 vccd1 vccd1 _13713_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06634__C _07995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11537_ _11547_/D _11537_/B vssd1 vssd1 vccd1 vccd1 _12814_/D sky130_fd_sc_hd__nor2_1
XFILLER_128_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06931__A _06955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ _14097_/Z _09068_/X _11499_/B vssd1 vssd1 vccd1 vccd1 _11469_/B sky130_fd_sc_hd__mux2_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ _13660_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__or2_1
XANTENNA__11373__A1 _12773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _12762_/Q _13937_/A vssd1 vssd1 vccd1 vccd1 _11400_/D sky130_fd_sc_hd__xor2_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09961__B _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11284__A _11312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__A2 _08455_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ _07630_/A _07641_/B _07635_/C vssd1 vssd1 vccd1 vccd1 _07631_/A sky130_fd_sc_hd__or3_1
XFILLER_81_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07561_ _08197_/A vssd1 vssd1 vccd1 vccd1 _08103_/B sky130_fd_sc_hd__clkbuf_1
X_09300_ _09329_/B _09329_/C _09300_/C vssd1 vssd1 vccd1 vccd1 _09306_/C sky130_fd_sc_hd__and3_1
X_06512_ _06521_/A _06512_/B _06512_/C vssd1 vssd1 vccd1 vccd1 _06513_/A sky130_fd_sc_hd__or3_1
XANTENNA__09689__A _10988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07492_ _07519_/A vssd1 vssd1 vccd1 vccd1 _07504_/A sky130_fd_sc_hd__clkbuf_1
X_09231_ _12236_/Q vssd1 vssd1 vccd1 vccd1 _09317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06443_ _06451_/A _06449_/B vssd1 vssd1 vccd1 vccd1 _06444_/A sky130_fd_sc_hd__or2_1
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09162_ _09162_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _09162_/X sky130_fd_sc_hd__or2_1
X_06374_ _11410_/A vssd1 vssd1 vccd1 vccd1 _07861_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_147_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08113_ _08122_/A _08113_/B _08122_/C vssd1 vssd1 vccd1 vccd1 _08114_/A sky130_fd_sc_hd__or3_1
XFILLER_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13939__A _13939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ input25/X input26/X vssd1 vssd1 vccd1 vccd1 _11924_/B sky130_fd_sc_hd__or2b_2
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08044_ _08052_/A _08047_/B _08044_/C vssd1 vssd1 vccd1 vccd1 _08045_/A sky130_fd_sc_hd__or3_1
XFILLER_116_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09995_ _09997_/B _09992_/A _09994_/X vssd1 vssd1 vccd1 vccd1 _09996_/B sky130_fd_sc_hd__o21ai_1
XFILLER_135_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08946_ _09067_/A vssd1 vssd1 vccd1 vccd1 _08946_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11906__B _13362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08877_ _08805_/X _08809_/X _08815_/X _08818_/X _08831_/X _08876_/X vssd1 vssd1 vccd1
+ vccd1 _08877_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07828_ _07828_/A vssd1 vssd1 vccd1 vccd1 _07828_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07759_ _07769_/A _07766_/B _07761_/C vssd1 vssd1 vccd1 vccd1 _07760_/A sky130_fd_sc_hd__or3_1
XFILLER_25_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10770_ _10785_/D _10936_/A _10770_/C vssd1 vssd1 vccd1 vccd1 _10771_/A sky130_fd_sc_hd__and3b_1
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09429_ _09439_/A _09429_/B vssd1 vssd1 vccd1 vccd1 _09430_/A sky130_fd_sc_hd__and2_1
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12440_ _12443_/CLK _12440_/D vssd1 vssd1 vccd1 vccd1 _12440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12371_ _12404_/CLK _12371_/D vssd1 vssd1 vccd1 vccd1 _13500_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ _14110_/A _08236_/X vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__ebufn_8
X_11322_ _11064_/X _11312_/X _11321_/X _11319_/X vssd1 vssd1 vccd1 vccd1 _12757_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07847__A _07964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14041_ _14041_/A _07889_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[10] sky130_fd_sc_hd__ebufn_8
X_11253_ _11253_/A vssd1 vssd1 vccd1 vccd1 _12741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10204_ _13625_/A _12478_/Q _10214_/S vssd1 vssd1 vccd1 vccd1 _10205_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11184_ _11184_/A vssd1 vssd1 vccd1 vccd1 _11184_/X sky130_fd_sc_hd__buf_6
XFILLER_121_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10135_ _10149_/B _10135_/B _10135_/C vssd1 vssd1 vccd1 vccd1 _10136_/A sky130_fd_sc_hd__and3b_1
XFILLER_121_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10066_ _10076_/D _10066_/B vssd1 vssd1 vccd1 vccd1 _12445_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13825_ _13825_/A _06764_/X vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13141__297 vssd1 vssd1 vccd1 vccd1 _13141__297/HI _13698_/A sky130_fd_sc_hd__conb_1
XFILLER_90_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13756_ _13756_/A _06952_/X vssd1 vssd1 vccd1 vccd1 _14108_/Z sky130_fd_sc_hd__ebufn_8
X_10968_ _13814_/A _12668_/Q _10972_/S vssd1 vssd1 vccd1 vccd1 _10969_/B sky130_fd_sc_hd__mux2_1
XFILLER_71_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12707_ _12743_/CLK _12707_/D vssd1 vssd1 vccd1 vccd1 _12707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13687_ _13687_/A _07127_/X vssd1 vssd1 vccd1 vccd1 _14103_/Z sky130_fd_sc_hd__ebufn_8
X_10899_ _10907_/C _10900_/B _10757_/X vssd1 vssd1 vccd1 vccd1 _10901_/A sky130_fd_sc_hd__o21ai_1
XFILLER_148_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12638_ _12820_/CLK _12638_/D vssd1 vssd1 vccd1 vccd1 _12638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13759__A _13759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ _12599_/CLK _12569_/D vssd1 vssd1 vccd1 vccd1 _12569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13035__191 vssd1 vssd1 vccd1 vccd1 _13035__191/HI _13478_/A sky130_fd_sc_hd__conb_1
XFILLER_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10183__A _10220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09972__A _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13494__A _13494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _12617_/Q _10773_/D _10863_/C _10773_/B _08779_/X _08780_/X vssd1 vssd1 vccd1
+ vccd1 _08800_/X sky130_fd_sc_hd__mux4_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _13498_/A _09787_/B vssd1 vssd1 vccd1 vccd1 _09780_/X sky130_fd_sc_hd__or2_1
X_06992_ _06992_/A vssd1 vssd1 vccd1 vccd1 _06992_/X sky130_fd_sc_hd__clkbuf_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _12616_/Q vssd1 vssd1 vccd1 vccd1 _10806_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10630__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08662_ _09396_/B vssd1 vssd1 vccd1 vccd1 _13556_/A sky130_fd_sc_hd__buf_6
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07613_ _07616_/A _07613_/B _07621_/C vssd1 vssd1 vccd1 vccd1 _07614_/A sky130_fd_sc_hd__or3_1
XFILLER_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08593_ _10098_/B _12447_/Q _12448_/Q _12449_/Q _08553_/X _08554_/X vssd1 vssd1 vccd1
+ vccd1 _08593_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07544_ _07544_/A vssd1 vssd1 vccd1 vccd1 _07544_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07475_ _07475_/A vssd1 vssd1 vccd1 vccd1 _07475_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09214_ _09211_/X _09214_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09215_/A sky130_fd_sc_hd__and3b_1
X_06426_ _06426_/A vssd1 vssd1 vccd1 vccd1 _06426_/X sky130_fd_sc_hd__clkbuf_1
X_09145_ _09145_/A vssd1 vssd1 vccd1 vccd1 _09145_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09866__B _13559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06357_ _06359_/A _06362_/B _06362_/C vssd1 vssd1 vccd1 vccd1 _06358_/A sky130_fd_sc_hd__or3_1
XFILLER_147_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09076_ _11687_/B _11687_/A _11695_/B _12851_/Q _09067_/X _09068_/X vssd1 vssd1 vccd1
+ vccd1 _09076_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06288_ _07827_/A _07845_/A _07979_/A vssd1 vssd1 vccd1 vccd1 _06289_/A sky130_fd_sc_hd__or3_1
XFILLER_30_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11189__A _11189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08027_ _08067_/A vssd1 vssd1 vccd1 vccd1 _08039_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_146_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09978_ _10049_/A vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_77_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11636__B _11682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08929_ _13969_/A vssd1 vssd1 vccd1 vccd1 _08929_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07833__C _08180_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11940_ _09625_/A _14035_/A _11940_/S vssd1 vssd1 vccd1 vccd1 _11941_/B sky130_fd_sc_hd__mux2_1
XFILLER_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11871_ _11888_/A vssd1 vssd1 vccd1 vccd1 _11886_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13610_ _13610_/A _07337_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10822_ _12632_/Q vssd1 vssd1 vccd1 vccd1 _10869_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ _13541_/A _07514_/X vssd1 vssd1 vccd1 vccd1 _13765_/Z sky130_fd_sc_hd__ebufn_8
X_10753_ _10806_/A _10760_/D vssd1 vssd1 vccd1 vccd1 _10774_/B sky130_fd_sc_hd__and2_1
XFILLER_111_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _13472_/A _07695_/X vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__ebufn_8
X_10684_ _13725_/A _10684_/B vssd1 vssd1 vccd1 vccd1 _10684_/X sky130_fd_sc_hd__or2_1
XFILLER_139_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09769__A1 _09767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _12470_/CLK _12423_/D vssd1 vssd1 vccd1 vccd1 _12423_/Q sky130_fd_sc_hd__dfxtp_1
X_13019__175 vssd1 vssd1 vccd1 vccd1 _13019__175/HI _13446_/A sky130_fd_sc_hd__conb_1
XFILLER_138_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07577__A _07590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12354_ _12356_/CLK _12354_/D vssd1 vssd1 vccd1 vccd1 _12354_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06481__A _06481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ _13878_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11305_/X sky130_fd_sc_hd__or2_1
XFILLER_114_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12285_ _12290_/CLK _12285_/D vssd1 vssd1 vccd1 vccd1 _12285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14024_ _14024_/A _08063_/X vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__ebufn_8
X_11236_ _11239_/A _11236_/B vssd1 vssd1 vccd1 vccd1 _11237_/A sky130_fd_sc_hd__and2_1
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11167_ _10648_/X _11155_/X _11165_/X _11166_/X vssd1 vssd1 vccd1 vccd1 _12714_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10118_ _10130_/D vssd1 vssd1 vccd1 vccd1 _10126_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11098_ _13846_/A _12701_/Q _11101_/S vssd1 vssd1 vccd1 vccd1 _11099_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08201__A _08228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10049_ _10049_/A vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__buf_2
XANTENNA__11500__A1 _13980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13808_ _13808_/A _06811_/X vssd1 vssd1 vccd1 vccd1 _14064_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13739_ _13739_/A _06994_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[28] sky130_fd_sc_hd__ebufn_8
XANTENNA__09967__A _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07260_ _07266_/A _07263_/B _07260_/C vssd1 vssd1 vccd1 vccd1 _07261_/A sky130_fd_sc_hd__or3_1
XFILLER_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07191_ _07191_/A vssd1 vssd1 vccd1 vccd1 _07191_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_83_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10625__B _13745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ _09773_/X _09888_/X _09900_/X _09892_/X vssd1 vssd1 vccd1 vccd1 _12400_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_98_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09832_ _09832_/A vssd1 vssd1 vccd1 vccd1 _12385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _10659_/A vssd1 vssd1 vccd1 vccd1 _09763_/X sky130_fd_sc_hd__buf_6
X_06975_ _07417_/A _06977_/B vssd1 vssd1 vccd1 vccd1 _06976_/A sky130_fd_sc_hd__or2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10360__B _13746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_21_clk_A _12881_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13952__A _13952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ _08582_/X _08591_/X _08588_/X _08593_/X _08663_/X _08670_/X vssd1 vssd1 vccd1
+ vccd1 _08714_/X sky130_fd_sc_hd__mux4_1
X_09694_ _09694_/A vssd1 vssd1 vccd1 vccd1 _12350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07950__A _08004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _12455_/Q vssd1 vssd1 vccd1 vccd1 _10111_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _08709_/A vssd1 vssd1 vccd1 vccd1 _08576_/X sky130_fd_sc_hd__buf_2
XFILLER_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_36_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07527_ _07531_/A _07531_/B _07538_/C vssd1 vssd1 vccd1 vccd1 _07528_/A sky130_fd_sc_hd__or3_1
XFILLER_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07458_ _07458_/A vssd1 vssd1 vccd1 vccd1 _07458_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06409_ _06409_/A vssd1 vssd1 vccd1 vccd1 _06409_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09596__B _13565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07389_ _07389_/A vssd1 vssd1 vccd1 vccd1 _07389_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09128_ _09134_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _09156_/A sky130_fd_sc_hd__nand2_1
XFILLER_136_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09059_ _12847_/Q vssd1 vssd1 vccd1 vccd1 _11687_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12070_ _14066_/A _12073_/B vssd1 vssd1 vccd1 vccd1 _12070_/X sky130_fd_sc_hd__or2_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11021_ _11021_/A _11021_/B _11021_/C _11021_/D vssd1 vssd1 vccd1 vccd1 _11022_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_104_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_109_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12972_ _12980_/CLK _12972_/D vssd1 vssd1 vccd1 vccd1 _14097_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input11_A peripheralBus_address[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _13377_/A _11922_/Y _11711_/B _09404_/A _13403_/A vssd1 vssd1 vccd1 vccd1
+ _12903_/D sky130_fd_sc_hd__o2111a_1
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11382__A _11723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _11888_/A vssd1 vssd1 vccd1 vccd1 _11869_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06476__A _08276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _10864_/B _10801_/B _10804_/Y vssd1 vssd1 vccd1 vccd1 _12628_/D sky130_fd_sc_hd__a21oi_1
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11785_ _11785_/A _11785_/B _11785_/C _11785_/D vssd1 vssd1 vccd1 vccd1 _11786_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_159_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09787__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13524_ _13524_/A _07559_/X vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_8
X_10736_ _13784_/A _13783_/A _10735_/X vssd1 vssd1 vccd1 vccd1 _10737_/C sky130_fd_sc_hd__or3b_2
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13455_ _13455_/A _08121_/X vssd1 vssd1 vccd1 vccd1 _13775_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_70_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10667_ _10667_/A vssd1 vssd1 vccd1 vccd1 _11039_/A sky130_fd_sc_hd__buf_2
XANTENNA__10726__A _13785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12406_ _12420_/CLK _12406_/D vssd1 vssd1 vccd1 vccd1 _13534_/A sky130_fd_sc_hd__dfxtp_1
X_13386_ _13386_/A _08342_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
X_10598_ _13723_/A _12579_/Q _10601_/S vssd1 vssd1 vccd1 vccd1 _10599_/B sky130_fd_sc_hd__mux2_1
XFILLER_142_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12337_ _12340_/CLK _12337_/D vssd1 vssd1 vccd1 vccd1 _13467_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12268_ _12274_/CLK _12268_/D vssd1 vssd1 vccd1 vccd1 _12268_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09914__A1 _09116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ _14007_/A _07948_/X vssd1 vssd1 vccd1 vccd1 _14007_/Z sky130_fd_sc_hd__ebufn_8
X_11219_ _11219_/A vssd1 vssd1 vccd1 vccd1 _12731_/D sky130_fd_sc_hd__clkbuf_1
X_12199_ _14102_/A _12206_/B vssd1 vssd1 vccd1 vccd1 _12199_/X sky130_fd_sc_hd__or2_1
XANTENNA__11276__B _13943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06760_ _06760_/A _06765_/B _06765_/C vssd1 vssd1 vccd1 vccd1 _06761_/A sky130_fd_sc_hd__or3_1
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06691_ _06691_/A vssd1 vssd1 vccd1 vccd1 _06691_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11292__A _11443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08430_ _09320_/D _12255_/Q _12256_/Q _09328_/A _08396_/X _08397_/X vssd1 vssd1 vccd1
+ vccd1 _08430_/X sky130_fd_sc_hd__mux4_2
XFILLER_91_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06817__C _07969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ _08361_/A vssd1 vssd1 vccd1 vccd1 _08361_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11788__A1 _13378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07312_ _07490_/A _07317_/B _07314_/C vssd1 vssd1 vccd1 vccd1 _07313_/A sky130_fd_sc_hd__or3_1
X_08292_ _08292_/A vssd1 vssd1 vccd1 vccd1 _08292_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07243_ _07243_/A vssd1 vssd1 vccd1 vccd1 _07243_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07174_ _07174_/A vssd1 vssd1 vccd1 vccd1 _07174_/X sky130_fd_sc_hd__clkbuf_1
X_13347__503 vssd1 vssd1 vccd1 vccd1 _13347__503/HI _14116_/A sky130_fd_sc_hd__conb_1
XANTENNA__10355__B _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07010__A _07979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13947__A _13947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09815_ _09815_/A vssd1 vssd1 vccd1 vccd1 _12380_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input3_A peripheralBus_address[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09746_ _09124_/X _09741_/X _09745_/X _09649_/X vssd1 vssd1 vccd1 vccd1 _12358_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06958_ _06960_/A _06965_/B vssd1 vssd1 vccd1 vccd1 _06959_/A sky130_fd_sc_hd__or2_1
XFILLER_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11914__B _13371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08567__S1 _08560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09677_ _09686_/A _09677_/B vssd1 vssd1 vccd1 vccd1 _09678_/A sky130_fd_sc_hd__and2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ _06889_/A vssd1 vssd1 vccd1 vccd1 _06889_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08628_ _10021_/C _10021_/B _10024_/B _10029_/B _08549_/X _08551_/X vssd1 vssd1 vccd1
+ vccd1 _08628_/X sky130_fd_sc_hd__mux4_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06296__A _07045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08559_ _13584_/A vssd1 vssd1 vccd1 vccd1 _08559_/X sky130_fd_sc_hd__buf_4
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11930__A _11998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ _11626_/A _11565_/X _11569_/X vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__o21ai_1
XFILLER_50_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10521_ _09753_/X _10511_/X _10520_/X _10425_/X vssd1 vssd1 vccd1 vccd1 _12554_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10452_ _10452_/A vssd1 vssd1 vccd1 vccd1 _12540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10383_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12122_ _12958_/Q _14100_/A _12135_/S vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12053_ _12924_/Q _13363_/A vssd1 vssd1 vccd1 vccd1 _12055_/C sky130_fd_sc_hd__xor2_1
XFILLER_111_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11004_ _12662_/Q _13936_/A vssd1 vssd1 vccd1 vccd1 _11004_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07590__A _07590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08558__S1 _08557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ _12962_/CLK _12955_/D vssd1 vssd1 vccd1 vccd1 _12955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11906_ _12890_/Q _13362_/A vssd1 vssd1 vccd1 vccd1 _11910_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10220__S _10220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _12886_/CLK _12886_/D vssd1 vssd1 vccd1 vccd1 _14014_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11837_ _14012_/Z _14012_/A _11840_/S vssd1 vssd1 vccd1 vccd1 _11838_/B sky130_fd_sc_hd__mux2_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _12867_/Q _13372_/A vssd1 vssd1 vccd1 vccd1 _11770_/C sky130_fd_sc_hd__xor2_1
XFILLER_14_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13507_ _13507_/A _07602_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
X_10719_ _14103_/Z _13783_/A _10723_/S vssd1 vssd1 vccd1 vccd1 _10720_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11699_ _12852_/Q _11699_/B vssd1 vssd1 vccd1 vccd1 _11702_/B sky130_fd_sc_hd__and2_1
X_13438_ _13438_/A _07783_/X vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_115_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ _13369_/A _08301_/X vssd1 vssd1 vccd1 vccd1 _13625_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07930_ _07930_/A vssd1 vssd1 vccd1 vccd1 _07930_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07861_ _07861_/A _07962_/B _07947_/B vssd1 vssd1 vccd1 vccd1 _07862_/A sky130_fd_sc_hd__or3_1
XFILLER_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09600_ _12323_/Q _13566_/A vssd1 vssd1 vccd1 vccd1 _09602_/C sky130_fd_sc_hd__xor2_1
XFILLER_96_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06812_ input4/X vssd1 vssd1 vccd1 vccd1 _09097_/A sky130_fd_sc_hd__inv_2
XFILLER_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07792_ _07796_/A _07792_/B _07801_/C vssd1 vssd1 vccd1 vccd1 _07793_/A sky130_fd_sc_hd__or3_1
XFILLER_95_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09531_ _09582_/S vssd1 vssd1 vccd1 vccd1 _09610_/B sky130_fd_sc_hd__clkbuf_2
X_06743_ _06743_/A vssd1 vssd1 vccd1 vccd1 _06743_/X sky130_fd_sc_hd__clkbuf_1
X_09462_ _09459_/Y _09460_/X _09461_/X vssd1 vssd1 vccd1 vccd1 _09468_/C sky130_fd_sc_hd__a21oi_1
X_06674_ _06674_/A vssd1 vssd1 vccd1 vccd1 _06674_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ _08406_/X _08407_/X _08409_/X _08411_/X _08479_/A _08383_/X vssd1 vssd1 vccd1
+ vccd1 _08413_/X sky130_fd_sc_hd__mux4_1
X_09393_ _09393_/A vssd1 vssd1 vccd1 vccd1 _12274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08344_ _08344_/A vssd1 vssd1 vccd1 vccd1 _08344_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08275_ _08275_/A vssd1 vssd1 vccd1 vccd1 _08275_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07226_ _07239_/A _07231_/B _07228_/C vssd1 vssd1 vccd1 vccd1 _07227_/A sky130_fd_sc_hd__or3_1
XFILLER_165_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07157_ _07157_/A vssd1 vssd1 vccd1 vccd1 _07157_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11909__B _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ _07094_/A _07091_/B _07088_/C vssd1 vssd1 vccd1 vccd1 _07089_/A sky130_fd_sc_hd__or3_1
XFILLER_78_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09729_ _12348_/Q _13558_/A vssd1 vssd1 vccd1 vccd1 _09730_/D sky130_fd_sc_hd__xor2_1
XFILLER_90_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12740_ _12758_/CLK _12740_/D vssd1 vssd1 vccd1 vccd1 _12740_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10672__A1 _10670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12671_ _12699_/CLK _12671_/D vssd1 vssd1 vccd1 vccd1 _12671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11622_ _11640_/A _11622_/B vssd1 vssd1 vccd1 vccd1 _11623_/C sky130_fd_sc_hd__nand2_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06754__A _11028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11553_ _11562_/C vssd1 vssd1 vccd1 vccd1 _11627_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10504_ _10504_/A _10504_/B _10504_/C _10504_/D vssd1 vssd1 vccd1 vccd1 _10505_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11484_ _11490_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _11485_/A sky130_fd_sc_hd__or2_1
XFILLER_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10435_ _10435_/A vssd1 vssd1 vccd1 vccd1 _12535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10366_ _12508_/Q _13750_/A vssd1 vssd1 vccd1 vccd1 _10367_/D sky130_fd_sc_hd__xor2_1
XFILLER_151_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12105_ _12953_/Q _14095_/A _12118_/S vssd1 vssd1 vccd1 vccd1 _12106_/B sky130_fd_sc_hd__mux2_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater113_A peripheralBus_data[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10297_ _13647_/A _12501_/Q _10375_/B vssd1 vssd1 vccd1 vccd1 _10298_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12036_ _12929_/Q _13368_/A vssd1 vssd1 vccd1 vccd1 _12040_/A sky130_fd_sc_hd__xor2_1
XFILLER_66_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output42_A _13785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13987_ _13987_/A _06321_/X vssd1 vssd1 vccd1 vccd1 _13987_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12938_ _12938_/CLK _12938_/D vssd1 vssd1 vccd1 vccd1 _14064_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06367__C _07822_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _12873_/CLK _12869_/D vssd1 vssd1 vccd1 vccd1 _12869_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06390_ _07845_/B vssd1 vssd1 vccd1 vccd1 _06400_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08060_ _08065_/A _08062_/B _08070_/C vssd1 vssd1 vccd1 vccd1 _08061_/A sky130_fd_sc_hd__or3_1
XFILLER_146_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07011_ _07019_/A _07019_/B vssd1 vssd1 vccd1 vccd1 _07012_/A sky130_fd_sc_hd__or2_1
XFILLER_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ _13972_/A vssd1 vssd1 vccd1 vccd1 _09071_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_142_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07913_ _07921_/A _07917_/B _07917_/C vssd1 vssd1 vccd1 vccd1 _07914_/A sky130_fd_sc_hd__or3_1
XFILLER_69_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08893_ _12655_/Q vssd1 vssd1 vccd1 vccd1 _10921_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07844_ _07844_/A vssd1 vssd1 vccd1 vccd1 _07844_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07775_ _07775_/A vssd1 vssd1 vccd1 vccd1 _07775_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09514_ _09526_/B vssd1 vssd1 vccd1 vccd1 _09524_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06726_ _11790_/A vssd1 vssd1 vccd1 vccd1 _11028_/B sky130_fd_sc_hd__buf_4
XFILLER_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09445_ _13435_/A _12287_/Q _09448_/S vssd1 vssd1 vccd1 vccd1 _09446_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10654__A1 _10652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06657_ _06659_/A _06664_/B _06664_/C vssd1 vssd1 vccd1 vccd1 _06658_/A sky130_fd_sc_hd__or3_1
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ _09377_/B _09370_/X _09377_/A vssd1 vssd1 vccd1 vccd1 _09380_/B sky130_fd_sc_hd__a21o_1
XFILLER_33_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06588_ _06588_/A vssd1 vssd1 vccd1 vccd1 _06588_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08327_ _08336_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08328_/A sky130_fd_sc_hd__or2_1
XFILLER_138_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08258_ _08258_/A vssd1 vssd1 vccd1 vccd1 _08258_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07209_ _07220_/A _07216_/B _07213_/C vssd1 vssd1 vccd1 vccd1 _07210_/A sky130_fd_sc_hd__or3_1
X_08189_ _08198_/A _08189_/B _08198_/C vssd1 vssd1 vccd1 vccd1 _08190_/A sky130_fd_sc_hd__or3_1
XFILLER_134_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10220_ _13630_/A _12483_/Q _10220_/S vssd1 vssd1 vccd1 vccd1 _10221_/B sky130_fd_sc_hd__mux2_1
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10151_ _10155_/C _10157_/B _10151_/C vssd1 vssd1 vccd1 vccd1 _10152_/A sky130_fd_sc_hd__and3b_1
XFILLER_133_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10082_ _10098_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10084_/B sky130_fd_sc_hd__or2_1
XFILLER_48_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13910_ _13910_/A _06527_/X vssd1 vssd1 vccd1 vccd1 _14070_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__07852__B _07854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__A _09125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ _13841_/A _06720_/X vssd1 vssd1 vccd1 vccd1 _14065_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13772_ _13772_/A _06912_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
X_10984_ _10984_/A vssd1 vssd1 vccd1 vccd1 _12672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08964__A _10939_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12723_ _12724_/CLK _12723_/D vssd1 vssd1 vccd1 vccd1 _13851_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252__408 vssd1 vssd1 vccd1 vccd1 _13252__408/HI _13923_/A sky130_fd_sc_hd__conb_1
X_12654_ _12660_/CLK _12654_/D vssd1 vssd1 vccd1 vccd1 _12654_/Q sky130_fd_sc_hd__dfxtp_1
X_11605_ _11605_/A vssd1 vssd1 vccd1 vccd1 _12830_/D sky130_fd_sc_hd__clkbuf_1
X_12585_ _12586_/CLK _12585_/D vssd1 vssd1 vccd1 vccd1 _13712_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11536_ _11626_/C _11533_/A _11521_/X vssd1 vssd1 vccd1 vccd1 _11537_/B sky130_fd_sc_hd__o21ai_1
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11467_ _09067_/X _11459_/X _11466_/X _11464_/X vssd1 vssd1 vccd1 vccd1 _12794_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10418_ _10285_/X _10409_/X _10417_/X _10412_/X vssd1 vssd1 vccd1 vccd1 _12530_/D
+ sky130_fd_sc_hd__o211a_1
X_11398_ _12772_/Q _13947_/A vssd1 vssd1 vccd1 vccd1 _11400_/C sky130_fd_sc_hd__xor2_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13146__302 vssd1 vssd1 vccd1 vccd1 _13146__302/HI _13703_/A sky130_fd_sc_hd__conb_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10349_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10350_/A sky130_fd_sc_hd__and2_1
XFILLER_140_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12019_ _12019_/A vssd1 vssd1 vccd1 vccd1 _12930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06378__B _07603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ _07590_/A vssd1 vssd1 vccd1 vccd1 _07575_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11833__A0 _13979_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06511_ _06511_/A vssd1 vssd1 vccd1 vccd1 _06511_/X sky130_fd_sc_hd__clkbuf_1
X_07491_ _07491_/A vssd1 vssd1 vccd1 vccd1 _07491_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09230_ _09235_/C _09230_/B vssd1 vssd1 vccd1 vccd1 _12235_/D sky130_fd_sc_hd__nor2_1
XFILLER_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06442_ _06442_/A vssd1 vssd1 vccd1 vccd1 _06451_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10628__B _13751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09161_ _09161_/A vssd1 vssd1 vccd1 vccd1 _09191_/B sky130_fd_sc_hd__clkbuf_1
X_06373_ _11457_/B vssd1 vssd1 vccd1 vccd1 _11410_/A sky130_fd_sc_hd__clkbuf_2
X_08112_ _08150_/A vssd1 vssd1 vccd1 vccd1 _08122_/A sky130_fd_sc_hd__buf_2
X_09092_ _11061_/A vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__buf_4
XFILLER_162_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08043_ _08043_/A vssd1 vssd1 vccd1 vccd1 _08043_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07656__C _07739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10363__B _13758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09962__C1 _09959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09994_ _10049_/A vssd1 vssd1 vccd1 vccd1 _09994_/X sky130_fd_sc_hd__buf_2
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07953__A _07999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ _12815_/Q vssd1 vssd1 vccd1 vccd1 _11571_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08876_ _08876_/A vssd1 vssd1 vccd1 vccd1 _08876_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07827_ _07827_/A _07827_/B _08349_/B vssd1 vssd1 vccd1 vccd1 _07828_/A sky130_fd_sc_hd__or3_1
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07758_ _07798_/A vssd1 vssd1 vccd1 vccd1 _07769_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_72_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06709_ _06722_/A vssd1 vssd1 vccd1 vccd1 _06719_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__09599__B _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ _07699_/A _07696_/B _07691_/C vssd1 vssd1 vccd1 vccd1 _07690_/A sky130_fd_sc_hd__or3_1
XFILLER_80_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09428_ _13430_/A _12282_/Q _09431_/S vssd1 vssd1 vccd1 vccd1 _09429_/B sky130_fd_sc_hd__mux2_1
XFILLER_80_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09359_ _09380_/A _09359_/B _09359_/C vssd1 vssd1 vccd1 vccd1 _09360_/A sky130_fd_sc_hd__and3_1
XFILLER_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12370_ _12404_/CLK _12370_/D vssd1 vssd1 vccd1 vccd1 _13499_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11321_ _13884_/A _11323_/B vssd1 vssd1 vccd1 vccd1 _11321_/X sky130_fd_sc_hd__or2_1
XFILLER_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ _14040_/A _07887_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[9] sky130_fd_sc_hd__ebufn_8
X_11252_ _11255_/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11253_/A sky130_fd_sc_hd__and2_1
XFILLER_134_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10203_ _10203_/A vssd1 vssd1 vccd1 vccd1 _12477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11183_ _10670_/X _11171_/X _11182_/X _11180_/X vssd1 vssd1 vccd1 vccd1 _12720_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10134_ _10133_/B _10133_/C _10137_/D _10137_/B vssd1 vssd1 vccd1 vccd1 _10135_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_95_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11385__A _12773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10065_ _10098_/C _10064_/B _09994_/X vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__06479__A _06481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13824_ _13824_/A _06766_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[17] sky130_fd_sc_hd__ebufn_8
XFILLER_16_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11815__A0 _09633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10967_ _10967_/A vssd1 vssd1 vccd1 vccd1 _12667_/D sky130_fd_sc_hd__clkbuf_1
X_13755_ _13755_/A _06954_/X vssd1 vssd1 vccd1 vccd1 _14075_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12706_ _12743_/CLK _12706_/D vssd1 vssd1 vccd1 vccd1 _12706_/Q sky130_fd_sc_hd__dfxtp_1
X_10898_ _10898_/A _10900_/B vssd1 vssd1 vccd1 vccd1 _12649_/D sky130_fd_sc_hd__nor2_1
X_13686_ _13686_/A _07129_/X vssd1 vssd1 vccd1 vccd1 _13974_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__07103__A _07248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12637_ _12820_/CLK _12637_/D vssd1 vssd1 vccd1 vccd1 _12637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12568_ _12586_/CLK _12568_/D vssd1 vssd1 vccd1 vccd1 _12568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11519_ _11658_/A _11628_/A vssd1 vssd1 vccd1 vccd1 _11523_/A sky130_fd_sc_hd__and2_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12499_ _12522_/CLK _12499_/D vssd1 vssd1 vccd1 vccd1 _13629_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13775__A _13775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06991_ _06995_/A _06995_/B vssd1 vssd1 vccd1 vccd1 _06992_/A sky130_fd_sc_hd__or2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11295__A _13874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _12615_/Q vssd1 vssd1 vccd1 vccd1 _10806_/C sky130_fd_sc_hd__clkbuf_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06389__A _08338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08661_ _08658_/X _08660_/X _08682_/S vssd1 vssd1 vccd1 vccd1 _09396_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07612_ _07612_/A vssd1 vssd1 vccd1 vccd1 _07612_/X sky130_fd_sc_hd__clkbuf_1
X_08592_ _12446_/Q vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07543_ _07545_/A _07545_/B _07551_/C vssd1 vssd1 vccd1 vccd1 _07544_/A sky130_fd_sc_hd__or3_1
X_13274__430 vssd1 vssd1 vccd1 vccd1 _13274__430/HI _13965_/A sky130_fd_sc_hd__conb_1
XFILLER_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07474_ _07478_/A _07484_/B vssd1 vssd1 vccd1 vccd1 _07475_/A sky130_fd_sc_hd__or2_1
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10358__B _13753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ _09281_/A vssd1 vssd1 vccd1 vccd1 _09271_/C sky130_fd_sc_hd__clkbuf_2
X_06425_ _06428_/A _06425_/B vssd1 vssd1 vccd1 vccd1 _06426_/A sky130_fd_sc_hd__or2_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13315__471 vssd1 vssd1 vccd1 vccd1 _13315__471/HI _14052_/A sky130_fd_sc_hd__conb_1
X_09144_ _09620_/A vssd1 vssd1 vccd1 vccd1 _10645_/A sky130_fd_sc_hd__buf_4
X_06356_ _06356_/A vssd1 vssd1 vccd1 vccd1 _06356_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09075_ _12850_/Q vssd1 vssd1 vccd1 vccd1 _11695_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06287_ _06287_/A vssd1 vssd1 vccd1 vccd1 _06287_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08026_ _08026_/A vssd1 vssd1 vccd1 vccd1 _08026_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11917__B _13367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09977_ _09977_/A vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08928_ _13968_/A vssd1 vssd1 vccd1 vccd1 _08928_/X sky130_fd_sc_hd__buf_2
X_08859_ _13779_/A vssd1 vssd1 vccd1 vccd1 _08859_/X sky130_fd_sc_hd__clkbuf_2
X_11870_ _11870_/A vssd1 vssd1 vccd1 vccd1 _12893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10821_ _10821_/A vssd1 vssd1 vccd1 vccd1 _12631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ _12617_/Q vssd1 vssd1 vccd1 vccd1 _10806_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13540_ _13540_/A _07516_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_111_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08019__A _08072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _13471_/A _07697_/X vssd1 vssd1 vccd1 vccd1 _14111_/Z sky130_fd_sc_hd__ebufn_8
X_10683_ _10288_/X _10673_/X _10681_/X _10682_/X vssd1 vssd1 vccd1 vccd1 _12597_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11025__A1 _13954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ _12470_/CLK _12422_/D vssd1 vssd1 vccd1 vccd1 _12422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ _12377_/CLK _12353_/D vssd1 vssd1 vccd1 vccd1 _12353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11304_ _10659_/X _11299_/X _11303_/X _11293_/X vssd1 vssd1 vccd1 vccd1 _12750_/D
+ sky130_fd_sc_hd__o211a_1
X_12284_ _12290_/CLK _12284_/D vssd1 vssd1 vccd1 vccd1 _12284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14023_ _14023_/A _08096_/X vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__ebufn_8
X_11235_ _13880_/A _12736_/Q _11248_/S vssd1 vssd1 vccd1 vccd1 _11236_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13595__A _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11166_ _11195_/A vssd1 vssd1 vccd1 vccd1 _11166_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10117_ _10117_/A vssd1 vssd1 vccd1 vccd1 _12455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11097_ _11206_/A vssd1 vssd1 vccd1 vccd1 _11112_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10048_ _10048_/A vssd1 vssd1 vccd1 vccd1 _12440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13258__414 vssd1 vssd1 vccd1 vccd1 _13258__414/HI _13929_/A sky130_fd_sc_hd__conb_1
XANTENNA__09313__A _09380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ _13807_/A _07862_/X vssd1 vssd1 vccd1 vccd1 _14063_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10459__A _10480_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11999_ _12033_/S vssd1 vssd1 vccd1 vccd1 _12012_/S sky130_fd_sc_hd__clkbuf_2
X_13738_ _13738_/A _06996_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[27] sky130_fd_sc_hd__ebufn_8
XANTENNA__09967__B _09967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13669_ _13669_/A _07174_/X vssd1 vssd1 vccd1 vccd1 _13765_/Z sky130_fd_sc_hd__ebufn_8
X_07190_ _07193_/A _07190_/B _07200_/C vssd1 vssd1 vccd1 vccd1 _07191_/A sky130_fd_sc_hd__or3_1
XFILLER_129_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _13528_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09900_/X sky130_fd_sc_hd__or2_1
XFILLER_160_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08815__S0 _08733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09831_ _09834_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _09832_/A sky130_fd_sc_hd__and2_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _09160_/X _09759_/X _09761_/X _09748_/X vssd1 vssd1 vccd1 vccd1 _12363_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ _06974_/A vssd1 vssd1 vccd1 vccd1 _07417_/A sky130_fd_sc_hd__buf_2
XFILLER_140_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _09399_/A vssd1 vssd1 vccd1 vccd1 _13563_/A sky130_fd_sc_hd__buf_4
XANTENNA_repeater75_A _14067_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09693_ _09705_/A _09693_/B vssd1 vssd1 vccd1 vccd1 _09694_/A sky130_fd_sc_hd__and2_1
XFILLER_67_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08644_ _12454_/Q vssd1 vssd1 vccd1 vccd1 _10111_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06847__A _06967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _08708_/A vssd1 vssd1 vccd1 vccd1 _08575_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07526_ _07553_/A vssd1 vssd1 vccd1 vccd1 _07538_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_07457_ _07466_/A _07459_/B vssd1 vssd1 vccd1 vccd1 _07458_/A sky130_fd_sc_hd__or2_1
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08671__A2 _08628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06408_ _06416_/A _06412_/B vssd1 vssd1 vccd1 vccd1 _06409_/A sky130_fd_sc_hd__or2_1
XFILLER_41_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07388_ _07396_/A _07391_/B _07388_/C vssd1 vssd1 vccd1 vccd1 _07389_/A sky130_fd_sc_hd__or3_1
X_13051__207 vssd1 vssd1 vccd1 vccd1 _13051__207/HI _13510_/A sky130_fd_sc_hd__conb_1
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09127_ _09919_/B vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06339_ _07045_/A vssd1 vssd1 vccd1 vccd1 _06349_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_108_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09058_ _08991_/X _08993_/X _08999_/X _09002_/X _09056_/X _09057_/X vssd1 vssd1 vccd1
+ vccd1 _09058_/X sky130_fd_sc_hd__mux4_1
X_08009_ _08009_/A vssd1 vssd1 vccd1 vccd1 _08009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11020_ _12665_/Q _13939_/A vssd1 vssd1 vccd1 vccd1 _11021_/D sky130_fd_sc_hd__xor2_1
XANTENNA__11647__B _11682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12971_ _12974_/CLK _12971_/D vssd1 vssd1 vccd1 vccd1 _14096_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11922_ _11922_/A _11922_/B vssd1 vssd1 vccd1 vccd1 _11922_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _11853_/A vssd1 vssd1 vccd1 vccd1 _12888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10279__A _10293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10804_ _10864_/B _10801_/B _10803_/X vssd1 vssd1 vccd1 vccd1 _10804_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ _12854_/Q _13359_/A vssd1 vssd1 vccd1 vccd1 _11785_/D sky130_fd_sc_hd__xor2_1
XFILLER_82_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _13523_/A _07563_/X vssd1 vssd1 vccd1 vccd1 _14035_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10735_ _10614_/B _10163_/C _10163_/D _10162_/A _13781_/A _13782_/A vssd1 vssd1 vccd1
+ vccd1 _10735_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13454_ _13454_/A _07740_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
X_10666_ _13719_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10666_/X sky130_fd_sc_hd__or2_1
XFILLER_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12405_ _12420_/CLK _12405_/D vssd1 vssd1 vccd1 vccd1 _13533_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13385_ _13385_/A _08340_/X vssd1 vssd1 vccd1 vccd1 _14121_/Z sky130_fd_sc_hd__ebufn_8
X_10597_ _10597_/A vssd1 vssd1 vccd1 vccd1 _12578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12336_ _12340_/CLK _12336_/D vssd1 vssd1 vccd1 vccd1 _13466_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_142_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11838__A _11852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10164__D _10613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ _12912_/CLK _12267_/D vssd1 vssd1 vccd1 vccd1 _12267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10742__A _10885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ _11221_/A _11218_/B vssd1 vssd1 vccd1 vccd1 _11219_/A sky130_fd_sc_hd__and2_1
X_14006_ _14006_/A _07961_/X vssd1 vssd1 vccd1 vccd1 _14070_/Z sky130_fd_sc_hd__ebufn_8
X_12198_ _10659_/A _12195_/X _12197_/X _12187_/X vssd1 vssd1 vccd1 vccd1 _12976_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11149_ _11149_/A _11149_/B _11149_/C vssd1 vssd1 vccd1 vccd1 _11149_/Y sky130_fd_sc_hd__nor3_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11573__A _11689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06690_ _06701_/A _06692_/B _06692_/C vssd1 vssd1 vccd1 vccd1 _06691_/A sky130_fd_sc_hd__or3_1
XANTENNA__06667__A _11156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08360_ _08364_/A _08364_/B _08360_/C vssd1 vssd1 vccd1 vccd1 _08361_/A sky130_fd_sc_hd__or3_1
XFILLER_51_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07311_ _07311_/A vssd1 vssd1 vccd1 vccd1 _07311_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11788__A2 _11787_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08291_ _08300_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08292_/A sky130_fd_sc_hd__or2_1
X_07242_ _07253_/A _07250_/B _07246_/C vssd1 vssd1 vccd1 vccd1 _07243_/A sky130_fd_sc_hd__or3_1
X_07173_ _07180_/A _07177_/B _07173_/C vssd1 vssd1 vccd1 vccd1 _07174_/A sky130_fd_sc_hd__or3_1
XFILLER_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10652__A _10652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14124__A _14124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10371__B _13743_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__A _08122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09814_ _09817_/A _09814_/B vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__and2_1
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09745_ _13487_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09745_/X sky130_fd_sc_hd__or2_1
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06957_ _06957_/A vssd1 vssd1 vccd1 vccd1 _06957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _13492_/A _12346_/Q _09685_/S vssd1 vssd1 vccd1 vccd1 _09677_/B sky130_fd_sc_hd__mux2_1
X_06888_ _06890_/A _06898_/B _06898_/C vssd1 vssd1 vccd1 vccd1 _06889_/A sky130_fd_sc_hd__or3_1
XFILLER_55_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _12432_/Q vssd1 vssd1 vccd1 vccd1 _10021_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09888__A _09902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _12429_/Q _12430_/Q _12431_/Q _12432_/Q _08556_/X _08557_/X vssd1 vssd1 vccd1
+ vccd1 _08558_/X sky130_fd_sc_hd__mux4_2
X_07509_ _07509_/A vssd1 vssd1 vccd1 vccd1 _07509_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08489_ _08455_/X _08461_/X _08458_/X _08488_/X _08470_/X _09152_/A vssd1 vssd1 vccd1
+ vccd1 _08489_/X sky130_fd_sc_hd__mux4_1
X_12994__150 vssd1 vssd1 vccd1 vccd1 _12994__150/HI _13405_/A sky130_fd_sc_hd__conb_1
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10520_ _13682_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _10520_/X sky130_fd_sc_hd__or2_1
XFILLER_156_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10451_ _10461_/A _10451_/B vssd1 vssd1 vccd1 vccd1 _10452_/A sky130_fd_sc_hd__and2_1
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10382_ _13647_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10382_/X sky130_fd_sc_hd__or2_1
X_12121_ _12154_/S vssd1 vssd1 vccd1 vccd1 _12135_/S sky130_fd_sc_hd__buf_2
XANTENNA__11658__A _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12052_ _12928_/Q _13367_/A vssd1 vssd1 vccd1 vccd1 _12055_/B sky130_fd_sc_hd__xor2_1
XFILLER_151_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08032__A _08072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ _12662_/Q _13936_/A vssd1 vssd1 vccd1 vccd1 _11003_/X sky130_fd_sc_hd__or2_1
XFILLER_93_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_82_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12954_ _12981_/CLK _12954_/D vssd1 vssd1 vccd1 vccd1 _12954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11905_ _11905_/A _11905_/B _11905_/C _11905_/D vssd1 vssd1 vccd1 vccd1 _11922_/A
+ sky130_fd_sc_hd__or4_1
X_13220__376 vssd1 vssd1 vccd1 vccd1 _13220__376/HI _13859_/A sky130_fd_sc_hd__conb_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ _12886_/CLK _12885_/D vssd1 vssd1 vccd1 vccd1 _14013_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _11888_/A vssd1 vssd1 vccd1 vccd1 _11852_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_97_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08635__A2 _08628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11767_ _12865_/Q _13370_/A vssd1 vssd1 vccd1 vccd1 _11770_/B sky130_fd_sc_hd__xor2_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13506_ _13506_/A _07607_/X vssd1 vssd1 vccd1 vccd1 _13666_/Z sky130_fd_sc_hd__ebufn_8
X_10718_ _10718_/A vssd1 vssd1 vccd1 vccd1 _12607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11698_ _12852_/Q _11699_/B _11576_/X vssd1 vssd1 vccd1 vccd1 _11700_/A sky130_fd_sc_hd__o21ai_1
XFILLER_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13437_ _13437_/A _07786_/X vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA_clkbuf_leaf_20_clk_A _12881_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10649_ _13714_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10649_/X sky130_fd_sc_hd__or2_1
XFILLER_161_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13114__270 vssd1 vssd1 vccd1 vccd1 _13114__270/HI _13639_/A sky130_fd_sc_hd__conb_1
X_13368_ _13368_/A _08298_/X vssd1 vssd1 vccd1 vccd1 _14104_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_115_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12319_ _12334_/CLK _12319_/D vssd1 vssd1 vccd1 vccd1 _12319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_35_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09899__A1 _09770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _07860_/A vssd1 vssd1 vccd1 vccd1 _07860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06811_ _06811_/A vssd1 vssd1 vccd1 vccd1 _06811_/X sky130_fd_sc_hd__clkbuf_1
X_07791_ _07791_/A vssd1 vssd1 vccd1 vccd1 _07791_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09530_ _13595_/A _09791_/B vssd1 vssd1 vccd1 vccd1 _09582_/S sky130_fd_sc_hd__and2_2
X_06742_ _06746_/A _06751_/B _06751_/C vssd1 vssd1 vccd1 vccd1 _06743_/A sky130_fd_sc_hd__or3_1
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09461_ _12280_/Q _13556_/A vssd1 vssd1 vccd1 vccd1 _09461_/X sky130_fd_sc_hd__xor2_1
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06673_ _06673_/A _06678_/B _06678_/C vssd1 vssd1 vccd1 vccd1 _06674_/A sky130_fd_sc_hd__or3_1
XANTENNA__09204__C _09372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08412_ _13394_/A vssd1 vssd1 vccd1 vccd1 _08479_/A sky130_fd_sc_hd__clkbuf_2
X_09392_ _09392_/A _09392_/B vssd1 vssd1 vccd1 vccd1 _09393_/A sky130_fd_sc_hd__and2_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08343_ _08347_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08344_/A sky130_fd_sc_hd__or2_1
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_108_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _08276_/A _08274_/B _08276_/C vssd1 vssd1 vccd1 vccd1 _08275_/A sky130_fd_sc_hd__or3_1
XFILLER_138_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10366__B _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07225_ _07225_/A vssd1 vssd1 vccd1 vccd1 _07225_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__07021__A _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07156_ _07166_/A _07163_/B _07160_/C vssd1 vssd1 vccd1 vccd1 _07157_/A sky130_fd_sc_hd__or3_1
XFILLER_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06860__A _06967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11478__A _14068_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07087_ _07087_/A vssd1 vssd1 vccd1 vccd1 _07087_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163__319 vssd1 vssd1 vccd1 vccd1 _13163__319/HI _13736_/A sky130_fd_sc_hd__conb_1
XFILLER_59_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07989_ _07997_/A _08005_/B _07993_/C vssd1 vssd1 vccd1 vccd1 _07990_/A sky130_fd_sc_hd__or3_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11449__A1 _11064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ _12356_/Q _13566_/A vssd1 vssd1 vccd1 vccd1 _09730_/C sky130_fd_sc_hd__xor2_1
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09659_ _13487_/A _12341_/Q _09738_/B vssd1 vssd1 vccd1 vccd1 _09660_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12687_/CLK _12670_/D vssd1 vssd1 vccd1 vccd1 _12670_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13057__213 vssd1 vssd1 vccd1 vccd1 _13057__213/HI _13516_/A sky130_fd_sc_hd__conb_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11640_/A _11622_/B vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__or2_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11552_ _11576_/A vssd1 vssd1 vccd1 vccd1 _11703_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__08027__A _08067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10503_ _12534_/Q _13743_/A vssd1 vssd1 vccd1 vccd1 _10504_/D sky130_fd_sc_hd__xor2_1
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11483_ _13974_/Z _13974_/A _11489_/S vssd1 vssd1 vccd1 vccd1 _11484_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09578__A0 _13469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ _10444_/A _10434_/B vssd1 vssd1 vccd1 vccd1 _10435_/A sky130_fd_sc_hd__and2_1
XANTENNA__06770__A _06809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10365_ _12503_/Q _13745_/A vssd1 vssd1 vccd1 vccd1 _10367_/C sky130_fd_sc_hd__xor2_1
XFILLER_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _12154_/S vssd1 vssd1 vccd1 vccd1 _12118_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_112_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10348_/S vssd1 vssd1 vccd1 vccd1 _10375_/B sky130_fd_sc_hd__buf_2
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12035_ _12035_/A vssd1 vssd1 vccd1 vccd1 _12935_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_repeater106_A _13987_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13986_ _13986_/A _06324_/X vssd1 vssd1 vccd1 vccd1 _14082_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_46_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output35_A _13402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12937_ _12946_/CLK _12937_/D vssd1 vssd1 vccd1 vccd1 _14063_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _12886_/CLK _12868_/D vssd1 vssd1 vccd1 vccd1 _12868_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11673__B1_N _11582_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11819_ _11888_/A vssd1 vssd1 vccd1 vccd1 _11834_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12799_/CLK _12799_/D vssd1 vssd1 vccd1 vccd1 _13973_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07010_ _07979_/B vssd1 vssd1 vccd1 vccd1 _07019_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06680__A _06680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08961_ _08955_/X _08957_/X _08959_/X _08960_/X _08952_/X _08953_/X vssd1 vssd1 vccd1
+ vccd1 _08961_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08103__C _08110_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07912_ _07912_/A vssd1 vssd1 vccd1 vccd1 _07912_/X sky130_fd_sc_hd__clkbuf_1
X_08892_ _08768_/X _08772_/X _08771_/X _08773_/X _08769_/X _08850_/X vssd1 vssd1 vccd1
+ vccd1 _08892_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07843_ _07843_/A _07854_/B _07852_/C vssd1 vssd1 vccd1 vccd1 _07844_/A sky130_fd_sc_hd__or3_1
XFILLER_69_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07774_ _07782_/A _07779_/B _07774_/C vssd1 vssd1 vccd1 vccd1 _07775_/A sky130_fd_sc_hd__or3_1
X_09513_ _09513_/A vssd1 vssd1 vccd1 vccd1 _09513_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06725_ _06725_/A _06725_/B vssd1 vssd1 vccd1 vccd1 _11790_/A sky130_fd_sc_hd__or2_4
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06656_ _06656_/A vssd1 vssd1 vccd1 vccd1 _06656_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11851__A1 _14032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _09444_/A vssd1 vssd1 vccd1 vccd1 _12286_/D sky130_fd_sc_hd__clkbuf_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ _09377_/B _09370_/X _09374_/Y vssd1 vssd1 vccd1 vccd1 _12269_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__10377__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06587_ _06597_/A _06589_/B _06589_/C vssd1 vssd1 vccd1 vccd1 _06588_/A sky130_fd_sc_hd__or3_1
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08326_ _08338_/A vssd1 vssd1 vccd1 vccd1 _08336_/A sky130_fd_sc_hd__clkbuf_1
X_08257_ _08264_/A _08261_/B _08264_/C vssd1 vssd1 vccd1 vccd1 _08258_/A sky130_fd_sc_hd__or3_1
XFILLER_138_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07208_ _07208_/A vssd1 vssd1 vccd1 vccd1 _07220_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08188_ _08228_/A vssd1 vssd1 vccd1 vccd1 _08198_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_07139_ _07139_/A vssd1 vssd1 vccd1 vccd1 _07139_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10150_ _10149_/B _10149_/C _10149_/A vssd1 vssd1 vccd1 vccd1 _10151_/C sky130_fd_sc_hd__a21o_1
XFILLER_121_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10081_ _12449_/Q vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09406__A _09846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09125__B _09125_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ _13840_/A _06724_/X vssd1 vssd1 vccd1 vccd1 _14064_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12095__A1 _11061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13771_ _13771_/A _06915_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
X_10983_ _10986_/A _10983_/B vssd1 vssd1 vccd1 vccd1 _10984_/A sky130_fd_sc_hd__and2_1
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ _12722_/CLK _12722_/D vssd1 vssd1 vccd1 vccd1 _13850_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13291__447 vssd1 vssd1 vccd1 vccd1 _13291__447/HI _13996_/A sky130_fd_sc_hd__conb_1
X_12653_ _12660_/CLK _12653_/D vssd1 vssd1 vccd1 vccd1 _12653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _11610_/C _11604_/B _11604_/C vssd1 vssd1 vccd1 vccd1 _11605_/A sky130_fd_sc_hd__and3b_1
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12584_ _12586_/CLK _12584_/D vssd1 vssd1 vccd1 vccd1 _13711_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11535_ _13967_/A _11628_/A _11572_/B vssd1 vssd1 vccd1 vccd1 _11547_/D sky130_fd_sc_hd__and3_1
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13332__488 vssd1 vssd1 vccd1 vccd1 _13332__488/HI _14085_/A sky130_fd_sc_hd__conb_1
XFILLER_128_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ _14064_/Z _11494_/B vssd1 vssd1 vccd1 vccd1 _11466_/X sky130_fd_sc_hd__or2_1
XFILLER_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10417_ _13659_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10417_/X sky130_fd_sc_hd__or2_1
X_11397_ _12775_/Q _13950_/A vssd1 vssd1 vccd1 vccd1 _11400_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08204__B _08208_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185__341 vssd1 vssd1 vccd1 vccd1 _13185__341/HI _13792_/A sky130_fd_sc_hd__conb_1
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _13662_/A _12516_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _10349_/B sky130_fd_sc_hd__mux2_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11846__A _13403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _10293_/B vssd1 vssd1 vccd1 vccd1 _10291_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12018_ _12030_/A _12018_/B vssd1 vssd1 vccd1 vccd1 _12019_/A sky130_fd_sc_hd__and2_1
X_13226__382 vssd1 vssd1 vccd1 vccd1 _13226__382/HI _13865_/A sky130_fd_sc_hd__conb_1
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09487__C1 _09192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13969_ _13969_/A _06370_/X vssd1 vssd1 vccd1 vccd1 _14097_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06510_ _06521_/A _06512_/B _06512_/C vssd1 vssd1 vccd1 vccd1 _06511_/A sky130_fd_sc_hd__or3_1
X_07490_ _07490_/A _08180_/B _07496_/C vssd1 vssd1 vccd1 vccd1 _07491_/A sky130_fd_sc_hd__or3_1
XFILLER_34_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06441_ _06441_/A vssd1 vssd1 vccd1 vccd1 _06441_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09160_ _11170_/A vssd1 vssd1 vccd1 vccd1 _09160_/X sky130_fd_sc_hd__buf_4
XANTENNA__09986__A _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06372_ _06372_/A vssd1 vssd1 vccd1 vccd1 _06372_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08111_ _08111_/A vssd1 vssd1 vccd1 vccd1 _08111_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08462__A0 _08452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09091_ _14107_/Z vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__buf_4
XFILLER_119_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08042_ _08052_/A _08047_/B _08044_/C vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__or3_1
XFILLER_147_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09993_ _09997_/B _09997_/C _09993_/C vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__and3_1
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ _12814_/Q vssd1 vssd1 vccd1 vccd1 _11626_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08130__A _11026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _10164_/C vssd1 vssd1 vccd1 vccd1 _13753_/A sky130_fd_sc_hd__buf_4
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09190__A1 _09092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07826_ _08351_/A vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__buf_2
XFILLER_72_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07757_ _07757_/A vssd1 vssd1 vccd1 vccd1 _07757_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06708_ _06753_/A vssd1 vssd1 vccd1 vccd1 _06719_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_44_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07688_ _07729_/A vssd1 vssd1 vccd1 vccd1 _07699_/A sky130_fd_sc_hd__clkbuf_1
X_09427_ _09427_/A vssd1 vssd1 vccd1 vccd1 _12281_/D sky130_fd_sc_hd__clkbuf_1
X_06639_ _11924_/A vssd1 vssd1 vccd1 vccd1 _11156_/B sky130_fd_sc_hd__buf_4
X_09358_ _09362_/B _09358_/B vssd1 vssd1 vccd1 vccd1 _09359_/C sky130_fd_sc_hd__nand2_1
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08309_ _08312_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08310_/A sky130_fd_sc_hd__or2_1
X_09289_ _09321_/B vssd1 vssd1 vccd1 vccd1 _09330_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11320_ _11061_/X _11312_/X _11318_/X _11319_/X vssd1 vssd1 vccd1 vccd1 _12756_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169__325 vssd1 vssd1 vccd1 vccd1 _13169__325/HI _13742_/A sky130_fd_sc_hd__conb_1
X_11251_ _13885_/A _12741_/Q _11254_/S vssd1 vssd1 vccd1 vccd1 _11252_/B sky130_fd_sc_hd__mux2_1
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09953__A0 _14104_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10202_ _10208_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _10203_/A sky130_fd_sc_hd__and2_1
XFILLER_109_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11182_ _13848_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11182_/X sky130_fd_sc_hd__or2_1
XFILLER_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10133_ _10137_/B _10133_/B _10133_/C _10137_/D vssd1 vssd1 vccd1 vccd1 _10149_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10570__A _10971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10064_ _10098_/C _10064_/B vssd1 vssd1 vccd1 vccd1 _10076_/D sky130_fd_sc_hd__and2_1
XANTENNA__09136__A _09379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13823_ _13823_/A _06772_/X vssd1 vssd1 vccd1 vccd1 _13983_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_63_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13754_ _13754_/A _06957_/X vssd1 vssd1 vccd1 vccd1 _14106_/Z sky130_fd_sc_hd__ebufn_8
X_10966_ _10969_/A _10966_/B vssd1 vssd1 vccd1 vccd1 _10967_/A sky130_fd_sc_hd__and2_1
XFILLER_71_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _12724_/CLK _12705_/D vssd1 vssd1 vccd1 vccd1 _12705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13685_ _13685_/A _07132_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[6] sky130_fd_sc_hd__ebufn_8
X_10897_ _10907_/D _10908_/A _10897_/C _10897_/D vssd1 vssd1 vccd1 vccd1 _10900_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12636_ _12820_/CLK _12636_/D vssd1 vssd1 vccd1 vccd1 _12636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12567_ _12589_/CLK _12567_/D vssd1 vssd1 vccd1 vccd1 _12567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11518_ _11518_/A _11518_/B _12808_/Q _12807_/Q vssd1 vssd1 vccd1 vccd1 _11628_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_157_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ _12522_/CLK _12498_/D vssd1 vssd1 vccd1 vccd1 _13628_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08215__A _08228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11449_ _11064_/X _11438_/X _11448_/X _11444_/X vssd1 vssd1 vccd1 vccd1 _12790_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09944__A0 _14037_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10003__B1 _09994_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10554__A1 _10552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06990_ _06990_/A vssd1 vssd1 vccd1 vccd1 _06990_/X sky130_fd_sc_hd__clkbuf_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _14099_/A _08207_/X vssd1 vssd1 vccd1 vccd1 _14099_/Z sky130_fd_sc_hd__ebufn_8
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08660_ _08591_/X _08595_/X _08593_/X _08659_/X _08695_/A _08652_/X vssd1 vssd1 vccd1
+ vccd1 _08660_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07611_ _07616_/A _07613_/B _07621_/C vssd1 vssd1 vccd1 vccd1 _07612_/A sky130_fd_sc_hd__or3_1
XFILLER_66_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08591_ _10052_/A _10099_/D _12444_/Q _12445_/Q _08556_/X _08557_/X vssd1 vssd1 vccd1
+ vccd1 _08591_/X sky130_fd_sc_hd__mux4_2
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ _07542_/A vssd1 vssd1 vccd1 vccd1 _07542_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__12200__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13003__159 vssd1 vssd1 vccd1 vccd1 _13003__159/HI _13414_/A sky130_fd_sc_hd__conb_1
X_07473_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07484_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_22_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09212_ _09210_/B _09201_/X _09210_/A vssd1 vssd1 vccd1 vccd1 _09214_/B sky130_fd_sc_hd__a21o_1
XFILLER_14_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06424_ _06424_/A vssd1 vssd1 vccd1 vccd1 _06424_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09143_ _14065_/Z vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__buf_4
X_06355_ _06359_/A _06362_/B _06362_/C vssd1 vssd1 vccd1 vccd1 _06356_/A sky130_fd_sc_hd__or3_1
XFILLER_147_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09074_ _12848_/Q vssd1 vssd1 vccd1 vccd1 _11687_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06286_ _07827_/A _07845_/A _07979_/A vssd1 vssd1 vccd1 vccd1 _06287_/A sky130_fd_sc_hd__or3_1
XFILLER_135_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08450__A3 _08447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08025_ _08025_/A _08033_/B _08030_/C vssd1 vssd1 vccd1 vccd1 _08026_/A sky130_fd_sc_hd__or3_1
XFILLER_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07964__A _07964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10545__A1 _10285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09976_ _09976_/A vssd1 vssd1 vccd1 vccd1 _12422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08927_ _12823_/Q vssd1 vssd1 vccd1 vccd1 _11639_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09163__A1 _09160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08858_ _10162_/D vssd1 vssd1 vccd1 vccd1 _13750_/A sky130_fd_sc_hd__buf_4
X_07809_ _07809_/A _07820_/B _07815_/C vssd1 vssd1 vccd1 vccd1 _07810_/A sky130_fd_sc_hd__or3_1
XFILLER_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08789_ _12635_/Q vssd1 vssd1 vccd1 vccd1 _10870_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10820_ _10833_/A _10820_/B _10820_/C vssd1 vssd1 vccd1 vccd1 _10821_/A sky130_fd_sc_hd__and3b_1
XFILLER_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10751_ _10760_/D _10751_/B vssd1 vssd1 vccd1 vccd1 _12616_/D sky130_fd_sc_hd__nor2_1
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _13470_/A _07700_/X vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10682_ _11039_/A vssd1 vssd1 vccd1 vccd1 _10682_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12421_ _12659_/CLK _12421_/D vssd1 vssd1 vccd1 vccd1 _12421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12352_ _12367_/CLK _12352_/D vssd1 vssd1 vccd1 vccd1 _12352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08035__A _08035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11303_ _13877_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11303_/X sky130_fd_sc_hd__or2_1
XFILLER_126_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12283_ _12301_/CLK _12283_/D vssd1 vssd1 vccd1 vccd1 _12283_/Q sky130_fd_sc_hd__dfxtp_1
X_14022_ _14022_/A _08066_/X vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__ebufn_8
X_11234_ _11254_/S vssd1 vssd1 vccd1 vccd1 _11248_/S sky130_fd_sc_hd__buf_2
XFILLER_141_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11165_ _13842_/A _11168_/B vssd1 vssd1 vccd1 vccd1 _11165_/X sky130_fd_sc_hd__or2_1
XFILLER_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10116_ _10114_/X _10135_/B _10116_/C vssd1 vssd1 vccd1 vccd1 _10117_/A sky130_fd_sc_hd__and3b_1
XFILLER_67_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11096_ _11096_/A vssd1 vssd1 vccd1 vccd1 _12700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10047_ _10045_/X _10062_/B _10047_/C vssd1 vssd1 vccd1 vccd1 _10048_/A sky130_fd_sc_hd__and3b_1
XFILLER_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13297__453 vssd1 vssd1 vccd1 vccd1 _13297__453/HI _14018_/A sky130_fd_sc_hd__conb_1
XFILLER_63_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13806_ _13806_/A _06818_/X vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_16_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11998_ _11998_/A vssd1 vssd1 vccd1 vccd1 _12013_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13737_ _13737_/A _07000_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[26] sky130_fd_sc_hd__ebufn_8
X_10949_ _10952_/A _10949_/B vssd1 vssd1 vccd1 vccd1 _10950_/A sky130_fd_sc_hd__and2_1
XFILLER_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13338__494 vssd1 vssd1 vccd1 vccd1 _13338__494/HI _14091_/A sky130_fd_sc_hd__conb_1
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _12583_/CLK sky130_fd_sc_hd__clkbuf_16
X_13668_ _13668_/A _07178_/X vssd1 vssd1 vccd1 vccd1 _14084_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12619_ _12660_/CLK _12619_/D vssd1 vssd1 vccd1 vccd1 _12619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13599_ _13599_/A _07368_/X vssd1 vssd1 vccd1 vccd1 _14111_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_117_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13786__A _13786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08815__S1 _08735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09830_ _13530_/A _12385_/Q _09837_/S vssd1 vssd1 vccd1 vccd1 _09831_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09761_ _13492_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09761_/X sky130_fd_sc_hd__or2_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06973_/X sky130_fd_sc_hd__clkbuf_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08704_/X _08711_/X _08712_/S vssd1 vssd1 vccd1 vccd1 _09399_/A sky130_fd_sc_hd__mux2_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09692_ _13496_/A _12350_/Q _09704_/S vssd1 vssd1 vccd1 vccd1 _09693_/B sky130_fd_sc_hd__mux2_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09504__A _09631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08643_ _10099_/A _12449_/Q _10097_/A _10101_/B _08629_/X _08630_/X vssd1 vssd1 vccd1
+ vccd1 _08643_/X sky130_fd_sc_hd__mux4_2
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _12428_/Q vssd1 vssd1 vccd1 vccd1 _09997_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10369__B _13747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ _07525_/A vssd1 vssd1 vccd1 vccd1 _07525_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_61_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _12823_/CLK sky130_fd_sc_hd__clkbuf_16
X_07456_ _07468_/A vssd1 vssd1 vccd1 vccd1 _07466_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06407_ _06407_/A vssd1 vssd1 vccd1 vccd1 _06407_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07387_ _07387_/A vssd1 vssd1 vccd1 vccd1 _07387_/X sky130_fd_sc_hd__clkbuf_1
X_13090__246 vssd1 vssd1 vccd1 vccd1 _13090__246/HI _13599_/A sky130_fd_sc_hd__conb_1
XANTENNA__10385__A _11160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09126_ input25/X input26/X vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__and2b_2
X_06338_ _06462_/A vssd1 vssd1 vccd1 vccd1 _06349_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06269_ _10693_/A vssd1 vssd1 vccd1 vccd1 _08364_/A sky130_fd_sc_hd__clkbuf_4
X_09057_ _09057_/A vssd1 vssd1 vccd1 vccd1 _09057_/X sky130_fd_sc_hd__clkbuf_2
X_13131__287 vssd1 vssd1 vccd1 vccd1 _13131__287/HI _13672_/A sky130_fd_sc_hd__conb_1
XFILLER_163_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08008_ _08010_/A _08020_/B _08016_/C vssd1 vssd1 vccd1 vccd1 _08009_/A sky130_fd_sc_hd__or3_1
XFILLER_104_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11191__A1 _11189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09959_ _10256_/A vssd1 vssd1 vccd1 vccd1 _09959_/X sky130_fd_sc_hd__buf_2
XFILLER_77_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12970_ _12981_/CLK _12970_/D vssd1 vssd1 vccd1 vccd1 _14095_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11921_ _11921_/A _11921_/B _11921_/C vssd1 vssd1 vccd1 vccd1 _11922_/B sky130_fd_sc_hd__or3_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025__181 vssd1 vssd1 vccd1 vccd1 _13025__181/HI _13452_/A sky130_fd_sc_hd__conb_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _11852_/A _11852_/B vssd1 vssd1 vccd1 vccd1 _11853_/A sky130_fd_sc_hd__and2_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _10803_/A vssd1 vssd1 vccd1 vccd1 _10803_/X sky130_fd_sc_hd__buf_2
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _12858_/Q _13363_/A vssd1 vssd1 vccd1 vccd1 _11785_/C sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_52_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _12687_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13522_ _13522_/A _07565_/X vssd1 vssd1 vccd1 vccd1 _14034_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_13_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10734_ _12614_/Q vssd1 vssd1 vccd1 vccd1 _10806_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13453_ _13453_/A _07743_/X vssd1 vssd1 vccd1 vccd1 _14029_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10295__A _13787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10665_ _10665_/A vssd1 vssd1 vccd1 vccd1 _10665_/X sky130_fd_sc_hd__buf_6
X_12404_ _12404_/CLK _12404_/D vssd1 vssd1 vccd1 vccd1 _13532_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13384_ _13384_/A _08337_/X vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11954__A0 _09636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10596_ _10602_/A _10596_/B vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__and2_1
X_12335_ _12340_/CLK _12335_/D vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater136_A peripheralBus_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12266_ _12912_/CLK _12266_/D vssd1 vssd1 vccd1 vccd1 _12266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14005_ _14005_/A _07959_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[6] sky130_fd_sc_hd__ebufn_8
X_11217_ _13875_/A _12731_/Q _11231_/S vssd1 vssd1 vccd1 vccd1 _11218_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09308__B _09372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12197_ _14101_/A _12206_/B vssd1 vssd1 vccd1 vccd1 _12197_/X sky130_fd_sc_hd__or2_1
XANTENNA__12015__A _12134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11148_ _11148_/A _11148_/B _11148_/C _11148_/D vssd1 vssd1 vccd1 vccd1 _11149_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_68_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11079_ _11079_/A vssd1 vssd1 vccd1 vccd1 _12695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09324__A _09347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__B _11649_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _12599_/CLK sky130_fd_sc_hd__clkbuf_16
X_07310_ _07490_/A _07317_/B _07314_/C vssd1 vssd1 vccd1 vccd1 _07311_/A sky130_fd_sc_hd__or3_1
X_08290_ _08314_/A vssd1 vssd1 vccd1 vccd1 _08300_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__10917__B _10917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_A _12917_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07241_ _07281_/A vssd1 vssd1 vccd1 vccd1 _07253_/A sky130_fd_sc_hd__clkbuf_1
X_07172_ _07172_/A vssd1 vssd1 vccd1 vccd1 _07172_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09813_ _13525_/A _12380_/Q _09820_/S vssd1 vssd1 vccd1 vccd1 _09814_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09118__A1 _09116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09744_ _09789_/B vssd1 vssd1 vccd1 vccd1 _09757_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_101_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06956_ _06960_/A _06965_/B vssd1 vssd1 vccd1 vccd1 _06957_/A sky130_fd_sc_hd__or2_1
X_13009__165 vssd1 vssd1 vccd1 vccd1 _13009__165/HI _13420_/A sky130_fd_sc_hd__conb_1
X_09675_ _09675_/A vssd1 vssd1 vccd1 vccd1 _12345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06887_ _07090_/A vssd1 vssd1 vccd1 vccd1 _06898_/C sky130_fd_sc_hd__clkbuf_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _09997_/A _12429_/Q _10029_/C _10021_/D _08549_/X _08551_/X vssd1 vssd1 vccd1
+ vccd1 _08626_/X sky130_fd_sc_hd__mux4_2
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _13585_/A vssd1 vssd1 vccd1 vccd1 _08557_/X sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_3_7_0_clk_A clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _12743_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07508_ _07517_/A _07517_/B _07510_/C vssd1 vssd1 vccd1 vccd1 _07509_/A sky130_fd_sc_hd__or3_1
X_08488_ _09362_/D _12264_/Q _12265_/Q _09362_/A _08368_/X _08370_/X vssd1 vssd1 vccd1
+ vccd1 _08488_/X sky130_fd_sc_hd__mux4_2
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07439_ _07439_/A vssd1 vssd1 vccd1 vccd1 _07439_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10450_ _13685_/A _12540_/Q _10456_/S vssd1 vssd1 vccd1 vccd1 _10451_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09109_ _12155_/A vssd1 vssd1 vccd1 vccd1 _09109_/X sky130_fd_sc_hd__clkbuf_2
X_10381_ _10423_/B vssd1 vssd1 vccd1 vccd1 _10392_/B sky130_fd_sc_hd__clkbuf_1
X_12120_ _12120_/A vssd1 vssd1 vccd1 vccd1 _12957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12051_ _12925_/Q _13364_/A vssd1 vssd1 vccd1 vccd1 _12055_/A sky130_fd_sc_hd__xor2_1
XFILLER_117_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09128__B _11460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11164__A1 _10645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11002_ _12674_/Q _13948_/A vssd1 vssd1 vccd1 vccd1 _11002_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06768__A _07406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11393__B _13941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09144__A _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12953_ _12981_/CLK _12953_/D vssd1 vssd1 vccd1 vccd1 _12953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11904_ _12888_/Q _13360_/A vssd1 vssd1 vccd1 vccd1 _11905_/D sky130_fd_sc_hd__xor2_1
XFILLER_73_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12886_/CLK _12884_/D vssd1 vssd1 vccd1 vccd1 _14012_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11835_ _11835_/A vssd1 vssd1 vccd1 vccd1 _12883_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08715__S0 _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _12863_/Q _13368_/A vssd1 vssd1 vccd1 vccd1 _11770_/A sky130_fd_sc_hd__xor2_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10737__B _11503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _13505_/A _07609_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
X_10717_ _10720_/A _10717_/B vssd1 vssd1 vccd1 vccd1 _10718_/A sky130_fd_sc_hd__or2_1
X_11697_ _12851_/Q _11694_/A _11696_/Y _11515_/X vssd1 vssd1 vccd1 vccd1 _12851_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13436_ _13436_/A _07788_/X vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10648_ _10648_/A vssd1 vssd1 vccd1 vccd1 _10648_/X sky130_fd_sc_hd__buf_4
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11849__A _11852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13367_ _13367_/A _08296_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[8] sky130_fd_sc_hd__ebufn_8
X_10579_ _10585_/A _10579_/B vssd1 vssd1 vccd1 vccd1 _10580_/A sky130_fd_sc_hd__and2_1
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12318_ _12334_/CLK _12318_/D vssd1 vssd1 vccd1 vccd1 _12318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12249_ _12251_/CLK _12249_/D vssd1 vssd1 vccd1 vccd1 _12249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06810_ _07857_/A _06830_/B _07947_/B vssd1 vssd1 vccd1 vccd1 _06811_/A sky130_fd_sc_hd__or3_1
XFILLER_56_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07790_ _07796_/A _07792_/B _07801_/C vssd1 vssd1 vccd1 vccd1 _07791_/A sky130_fd_sc_hd__or3_1
XANTENNA__06678__A _06686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06741_ _08195_/B vssd1 vssd1 vccd1 vccd1 _06751_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09460_ _12279_/Q _13555_/A vssd1 vssd1 vccd1 vccd1 _09460_/X sky130_fd_sc_hd__or2_1
XFILLER_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06672_ _06672_/A vssd1 vssd1 vccd1 vccd1 _06672_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08411_ _12257_/Q _12258_/Q _09343_/C _12260_/Q _08376_/X _08377_/X vssd1 vssd1 vccd1
+ vccd1 _08411_/X sky130_fd_sc_hd__mux4_2
XFILLER_52_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09391_ _12274_/Q _09391_/B vssd1 vssd1 vccd1 vccd1 _09392_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _12974_/CLK sky130_fd_sc_hd__clkbuf_16
X_08342_ _08342_/A vssd1 vssd1 vccd1 vccd1 _08342_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08273_ _08273_/A vssd1 vssd1 vccd1 vccd1 _08273_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07224_ _07239_/A _07231_/B _07228_/C vssd1 vssd1 vccd1 vccd1 _07225_/A sky130_fd_sc_hd__or3_1
XFILLER_164_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07956__B _07962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07155_ _07208_/A vssd1 vssd1 vccd1 vccd1 _07166_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_145_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07086_ _07094_/A _07091_/B _07088_/C vssd1 vssd1 vccd1 vccd1 _07087_/A sky130_fd_sc_hd__or3_1
XFILLER_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08133__A _08135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09339__A1 _09379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11494__A _13978_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07988_ _08022_/A vssd1 vssd1 vccd1 vccd1 _08005_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13243__399 vssd1 vssd1 vccd1 vccd1 _13243__399/HI _13898_/A sky130_fd_sc_hd__conb_1
X_09727_ _12353_/Q _13563_/A vssd1 vssd1 vccd1 vccd1 _09730_/B sky130_fd_sc_hd__xor2_1
XFILLER_101_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06939_ _06948_/A _06941_/B vssd1 vssd1 vccd1 vccd1 _06940_/A sky130_fd_sc_hd__or2_1
XFILLER_55_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09658_ _09711_/S vssd1 vssd1 vccd1 vccd1 _09738_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08609_ _12434_/Q vssd1 vssd1 vccd1 vccd1 _10024_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _12309_/Q _13552_/A vssd1 vssd1 vccd1 vccd1 _09589_/Y sky130_fd_sc_hd__nor2_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13096__252 vssd1 vssd1 vccd1 vccd1 _13096__252/HI _13605_/A sky130_fd_sc_hd__conb_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _12835_/Q vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11551_ _11551_/A vssd1 vssd1 vccd1 vccd1 _12817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10502_ _12539_/Q _13748_/A vssd1 vssd1 vccd1 vccd1 _10504_/C sky130_fd_sc_hd__xor2_1
X_13137__293 vssd1 vssd1 vccd1 vccd1 _13137__293/HI _13678_/A sky130_fd_sc_hd__conb_1
XFILLER_7_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11482_ _11482_/A vssd1 vssd1 vccd1 vccd1 _12799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10433_ _13680_/A _12535_/Q _10507_/B vssd1 vssd1 vccd1 vccd1 _10434_/B sky130_fd_sc_hd__mux2_1
XFILLER_136_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11388__B _11388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09139__A _11160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10364_ _12513_/Q _13755_/A vssd1 vssd1 vccd1 vccd1 _10367_/B sky130_fd_sc_hd__xor2_1
XFILLER_88_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ _13401_/A _12103_/B vssd1 vssd1 vccd1 vccd1 _12154_/S sky130_fd_sc_hd__nand2_2
XFILLER_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10295_ _13787_/A _10555_/B vssd1 vssd1 vccd1 vccd1 _10348_/S sky130_fd_sc_hd__and2_2
XFILLER_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12034_ _12115_/A _12034_/B vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__and2_1
XFILLER_2_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10896__B1 _10798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13985_ _13985_/A _06328_/X vssd1 vssd1 vccd1 vccd1 _14081_/Z sky130_fd_sc_hd__ebufn_8
X_12936_ _12969_/CLK _12936_/D vssd1 vssd1 vccd1 vccd1 _13376_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output28_A _13401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12867_ _12867_/CLK _12867_/D vssd1 vssd1 vccd1 vccd1 _12867_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _11929_/A vssd1 vssd1 vccd1 vccd1 _11888_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09266__B1 _09206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12798_ _12806_/CLK _12798_/D vssd1 vssd1 vccd1 vccd1 _13972_/A sky130_fd_sc_hd__dfxtp_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11749_ _11749_/A vssd1 vssd1 vccd1 vccd1 _12864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09975__C _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13419_ _13419_/A _07828_/X vssd1 vssd1 vccd1 vccd1 _13995_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11579__A _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09049__A _11384_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08960_ _12836_/Q _12837_/Q _12838_/Q _12839_/Q _08921_/X _08922_/X vssd1 vssd1 vccd1
+ vccd1 _08960_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_leaf_5_clk _12917_/CLK vssd1 vssd1 vccd1 vccd1 _12918_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07911_ _07921_/A _07917_/B _07917_/C vssd1 vssd1 vccd1 vccd1 _07912_/A sky130_fd_sc_hd__or3_1
XFILLER_130_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08891_ _10165_/A vssd1 vssd1 vccd1 vccd1 _13755_/A sky130_fd_sc_hd__buf_4
XFILLER_68_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10887__B1 _10798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ _08084_/A vssd1 vssd1 vccd1 vccd1 _07854_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07773_ _07773_/A vssd1 vssd1 vccd1 vccd1 _07773_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09512_ _13432_/A _09500_/X _09511_/X _09509_/X vssd1 vssd1 vccd1 vccd1 _12301_/D
+ sky130_fd_sc_hd__o211a_1
X_06724_ _06724_/A vssd1 vssd1 vccd1 vccd1 _06724_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _09455_/A _09443_/B vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__and2_1
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06655_ _06659_/A _06664_/B _06664_/C vssd1 vssd1 vccd1 vccd1 _06656_/A sky130_fd_sc_hd__or3_1
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09374_ _09377_/B _09370_/X _09392_/A vssd1 vssd1 vccd1 vccd1 _09374_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06586_ _06599_/A vssd1 vssd1 vccd1 vccd1 _06597_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__08128__A _08135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08325_ _08325_/A vssd1 vssd1 vccd1 vccd1 _08325_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08256_ _08256_/A vssd1 vssd1 vccd1 vccd1 _08256_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08480__A1 _08423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07207_ _07207_/A vssd1 vssd1 vccd1 vccd1 _07207_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08187_ _08240_/A vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_81_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07138_ _07152_/A _07145_/B _07142_/C vssd1 vssd1 vccd1 vccd1 _07139_/A sky130_fd_sc_hd__or3_1
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11001__B _13948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07069_ _07079_/A _07076_/B _07073_/C vssd1 vssd1 vccd1 vccd1 _07070_/A sky130_fd_sc_hd__or3_1
XFILLER_133_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_96_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ _10080_/A vssd1 vssd1 vccd1 vccd1 _12448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09193__C1 _09192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13770_ _13770_/A _06917_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
X_10982_ _13818_/A _12672_/Q _10990_/S vssd1 vssd1 vccd1 vccd1 _10983_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12721_ _12724_/CLK _12721_/D vssd1 vssd1 vccd1 vccd1 _13849_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12652_ _12652_/CLK _12652_/D vssd1 vssd1 vccd1 vccd1 _12652_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_34_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ _11631_/B _11595_/A _11642_/A _11641_/C vssd1 vssd1 vccd1 vccd1 _11604_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12583_ _12583_/CLK _12583_/D vssd1 vssd1 vccd1 vccd1 _13759_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_156_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11534_ _11626_/C _11626_/D _11625_/C _11625_/D vssd1 vssd1 vccd1 vccd1 _11572_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_11_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_49_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ _11689_/A _11459_/X _11463_/X _11464_/X vssd1 vssd1 vccd1 vccd1 _12793_/D
+ sky130_fd_sc_hd__o211a_1
X_10416_ _10414_/X _10409_/X _10415_/X _10412_/X vssd1 vssd1 vccd1 vccd1 _12529_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11396_ _12767_/Q _13942_/A vssd1 vssd1 vccd1 vccd1 _11400_/A sky130_fd_sc_hd__xor2_1
XFILLER_99_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10347_ _10347_/A vssd1 vssd1 vccd1 vccd1 _12515_/D sky130_fd_sc_hd__clkbuf_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10278_ _10278_/A vssd1 vssd1 vccd1 vccd1 _10278_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12017_ _12930_/Q _14073_/A _12029_/S vssd1 vssd1 vccd1 vccd1 _12018_/B sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_107_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13968_ _13968_/A _06372_/X vssd1 vssd1 vccd1 vccd1 _14064_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_19_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12919_ _12919_/CLK _12919_/D vssd1 vssd1 vccd1 vccd1 _14046_/A sky130_fd_sc_hd__dfxtp_1
X_13899_ _13899_/A _06560_/X vssd1 vssd1 vccd1 vccd1 _13995_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06440_ _06440_/A _06449_/B vssd1 vssd1 vccd1 vccd1 _06441_/A sky130_fd_sc_hd__or2_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06371_ _06822_/A _07822_/B _07822_/C vssd1 vssd1 vccd1 vccd1 _06372_/A sky130_fd_sc_hd__or3_1
XFILLER_159_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08110_ _08110_/A _08110_/B _08110_/C vssd1 vssd1 vccd1 vccd1 _08111_/A sky130_fd_sc_hd__or3_1
X_09090_ _10941_/D vssd1 vssd1 vccd1 vccd1 _13950_/A sky130_fd_sc_hd__buf_6
XANTENNA__08462__A1 _08455_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08041_ _08067_/A vssd1 vssd1 vccd1 vccd1 _08052_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_115_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09962__A1 _09092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ _09992_/A _09992_/B vssd1 vssd1 vccd1 vccd1 _12426_/D sky130_fd_sc_hd__nor2_1
XANTENNA_repeater98_A _14119_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08943_ _12808_/Q _11518_/B _11518_/A _11625_/D _08941_/X _08942_/X vssd1 vssd1 vccd1
+ vccd1 _08943_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_15_0_clk/X
+ sky130_fd_sc_hd__clkbuf_2
X_08874_ _08870_/X _08873_/X _08890_/S vssd1 vssd1 vccd1 vccd1 _10164_/C sky130_fd_sc_hd__mux2_1
XFILLER_57_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07825_ _09125_/B vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07756_ _07756_/A _07766_/B _07761_/C vssd1 vssd1 vccd1 vccd1 _07757_/A sky130_fd_sc_hd__or3_1
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06707_ _06707_/A vssd1 vssd1 vccd1 vccd1 _06707_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07687_ _07687_/A vssd1 vssd1 vccd1 vccd1 _07687_/X sky130_fd_sc_hd__clkbuf_1
X_09426_ _09439_/A _09426_/B vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__and2_1
X_06638_ input18/X _09102_/A _09096_/C _06725_/B vssd1 vssd1 vccd1 vccd1 _11924_/A
+ sky130_fd_sc_hd__or4_4
X_09357_ _09362_/B _09358_/B vssd1 vssd1 vccd1 vccd1 _09359_/B sky130_fd_sc_hd__or2_1
X_06569_ _06569_/A _06574_/B _06574_/C vssd1 vssd1 vccd1 vccd1 _06570_/A sky130_fd_sc_hd__or3_1
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08308_ _08308_/A vssd1 vssd1 vccd1 vccd1 _08308_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09288_ _09288_/A vssd1 vssd1 vccd1 vccd1 _12249_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10835__B _10917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08239_ _08239_/A vssd1 vssd1 vccd1 vccd1 _08239_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11250_ _11250_/A vssd1 vssd1 vccd1 vccd1 _12740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10201_ _13624_/A _12477_/Q _10214_/S vssd1 vssd1 vccd1 vccd1 _10202_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11947__A _11998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11181_ _10665_/X _11171_/X _11179_/X _11180_/X vssd1 vssd1 vccd1 vccd1 _12719_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10132_ _10129_/Y _10127_/C _10131_/X vssd1 vssd1 vccd1 vccd1 _12459_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__09417__A _09454_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08321__A _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07863__C _08349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10063_ _10063_/A vssd1 vssd1 vccd1 vccd1 _12444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input27_A rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13822_ _13822_/A _06774_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13753_ _13753_/A _06959_/X vssd1 vssd1 vccd1 vccd1 _14105_/Z sky130_fd_sc_hd__ebufn_8
X_10965_ _13813_/A _12667_/Q _10972_/S vssd1 vssd1 vccd1 vccd1 _10966_/B sky130_fd_sc_hd__mux2_1
XFILLER_141_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12704_ _12704_/CLK _12704_/D vssd1 vssd1 vccd1 vccd1 _12704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13684_ _13684_/A _07136_/X vssd1 vssd1 vccd1 vccd1 _14100_/Z sky130_fd_sc_hd__ebufn_8
X_10896_ _10907_/D _10895_/C _10798_/X vssd1 vssd1 vccd1 vccd1 _10898_/A sky130_fd_sc_hd__o21ai_1
XFILLER_93_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12635_ _12820_/CLK _12635_/D vssd1 vssd1 vccd1 vccd1 _12635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13402__A _13402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12566_ _12586_/CLK _12566_/D vssd1 vssd1 vccd1 vccd1 _13694_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11517_ _11517_/A _11517_/B vssd1 vssd1 vccd1 vccd1 _12809_/D sky130_fd_sc_hd__nor2_1
XFILLER_144_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _12522_/CLK _12497_/D vssd1 vssd1 vccd1 vccd1 _13627_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11448_ _13916_/A _11450_/B vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__or2_1
XFILLER_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11379_ _11929_/A vssd1 vssd1 vccd1 vccd1 _11801_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14098_ _14098_/A _08205_/X vssd1 vssd1 vccd1 vccd1 _14098_/Z sky130_fd_sc_hd__ebufn_8
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07610_ _07623_/A vssd1 vssd1 vccd1 vccd1 _07621_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_94_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08590_ _12443_/Q vssd1 vssd1 vccd1 vccd1 _10099_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__06686__A _06686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07541_ _07545_/A _07545_/B _07551_/C vssd1 vssd1 vccd1 vccd1 _07542_/A sky130_fd_sc_hd__or3_1
X_13042__198 vssd1 vssd1 vccd1 vccd1 _13042__198/HI _13485_/A sky130_fd_sc_hd__conb_1
XFILLER_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07472_ _07472_/A vssd1 vssd1 vccd1 vccd1 _07472_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09211_ _09347_/A _09318_/A vssd1 vssd1 vccd1 vccd1 _09211_/X sky130_fd_sc_hd__and2_1
X_06423_ _06428_/A _06425_/B vssd1 vssd1 vccd1 vccd1 _06424_/A sky130_fd_sc_hd__or2_1
XANTENNA__10936__A _10936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09142_ _09139_/X _09130_/X _09140_/X _09141_/X vssd1 vssd1 vccd1 vccd1 _12215_/D
+ sky130_fd_sc_hd__o211a_1
X_06354_ _06354_/A vssd1 vssd1 vccd1 vccd1 _06354_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09073_ _08951_/X _08957_/X _08955_/X _08959_/X _09024_/X _09030_/X vssd1 vssd1 vccd1
+ vccd1 _09073_/X sky130_fd_sc_hd__mux4_1
X_06285_ _06547_/A vssd1 vssd1 vccd1 vccd1 _07979_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08024_ _08024_/A vssd1 vssd1 vccd1 vccd1 _08024_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09975_ _09972_/X _09975_/B _10157_/B vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__and3b_1
XFILLER_115_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08926_ _08914_/X _08917_/X _08920_/X _08923_/X _08924_/X _08925_/X vssd1 vssd1 vccd1
+ vccd1 _08926_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08857_ _08851_/X _08856_/X _08890_/S vssd1 vssd1 vccd1 vccd1 _10162_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07808_ _08064_/A vssd1 vssd1 vccd1 vccd1 _07820_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08788_ _08781_/X _08782_/X _08783_/X _08787_/X _08748_/X _08749_/X vssd1 vssd1 vccd1
+ vccd1 _08788_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07739_ _07739_/A _07947_/B _07739_/C vssd1 vssd1 vccd1 vccd1 _07740_/A sky130_fd_sc_hd__or3_1
XFILLER_41_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10750_ _10806_/B _10742_/X _10749_/X vssd1 vssd1 vccd1 vccd1 _10751_/B sky130_fd_sc_hd__o21ai_1
XFILLER_158_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09409_ _09422_/A _09409_/B vssd1 vssd1 vccd1 vccd1 _09410_/A sky130_fd_sc_hd__and2_1
X_10681_ _13724_/A _10684_/B vssd1 vssd1 vccd1 vccd1 _10681_/X sky130_fd_sc_hd__or2_1
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12420_ _12420_/CLK _12420_/D vssd1 vssd1 vccd1 vccd1 _13596_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12351_ _12356_/CLK _12351_/D vssd1 vssd1 vccd1 vccd1 _12351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ _11170_/X _11299_/X _11301_/X _11293_/X vssd1 vssd1 vccd1 vccd1 _12749_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12282_ _12289_/CLK _12282_/D vssd1 vssd1 vccd1 vccd1 _12282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14021_ _14021_/A _08109_/X vssd1 vssd1 vccd1 vccd1 _14117_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_107_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ _11233_/A vssd1 vssd1 vccd1 vccd1 _12735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09147__A input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__B _13942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ _10645_/X _11155_/X _11163_/X _11068_/X vssd1 vssd1 vccd1 vccd1 _12713_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10115_ _10111_/B _10108_/B _10111_/A vssd1 vssd1 vccd1 vccd1 _10116_/C sky130_fd_sc_hd__a21o_1
XFILLER_96_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11095_ _11095_/A _11095_/B vssd1 vssd1 vccd1 vccd1 _11096_/A sky130_fd_sc_hd__and2_1
X_10046_ _10052_/D _10045_/C _10052_/C vssd1 vssd1 vccd1 vccd1 _10047_/C sky130_fd_sc_hd__a21o_1
XFILLER_48_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08901__A2 _08872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13805_ _13805_/A _06823_/X vssd1 vssd1 vccd1 vccd1 _14125_/Z sky130_fd_sc_hd__ebufn_8
X_11997_ _11997_/A vssd1 vssd1 vccd1 vccd1 _12924_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10948_ _13808_/A _12662_/Q _10955_/S vssd1 vssd1 vccd1 vccd1 _10949_/B sky130_fd_sc_hd__mux2_1
X_13736_ _13736_/A _07002_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[25] sky130_fd_sc_hd__ebufn_8
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ _13667_/A _07181_/X vssd1 vssd1 vccd1 vccd1 _14083_/Z sky130_fd_sc_hd__ebufn_8
X_10879_ _10881_/A _10872_/X _10878_/Y _10749_/X vssd1 vssd1 vccd1 vccd1 _12644_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12618_ _12660_/CLK _12618_/D vssd1 vssd1 vccd1 vccd1 _12618_/Q sky130_fd_sc_hd__dfxtp_1
X_13598_ _13598_/A _07370_/X vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__ebufn_8
X_12549_ _12599_/CLK _12549_/D vssd1 vssd1 vccd1 vccd1 _12549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09917__A1 _09120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _09789_/B vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__clkbuf_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06972_ _06972_/A _06977_/B vssd1 vssd1 vccd1 vccd1 _06973_/A sky130_fd_sc_hd__or2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _08568_/X _08654_/X _08680_/X _08710_/X _08632_/X _08634_/X vssd1 vssd1 vccd1
+ vccd1 _08711_/X sky130_fd_sc_hd__mux4_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09691_ _09711_/S vssd1 vssd1 vccd1 vccd1 _09704_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08642_ _12451_/Q vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _12422_/Q _12423_/Q _09981_/A _09997_/D _08549_/X _08551_/X vssd1 vssd1 vccd1
+ vccd1 _08573_/X sky130_fd_sc_hd__mux4_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07524_ _07531_/A _07531_/B _07524_/C vssd1 vssd1 vccd1 vccd1 _07525_/A sky130_fd_sc_hd__or3_1
XFILLER_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11660__B1 _11576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07455_ _07455_/A vssd1 vssd1 vccd1 vccd1 _07455_/X sky130_fd_sc_hd__clkbuf_1
X_06406_ _06416_/A _06412_/B vssd1 vssd1 vccd1 vccd1 _06407_/A sky130_fd_sc_hd__or2_1
XFILLER_10_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07386_ _07396_/A _07391_/B _07388_/C vssd1 vssd1 vccd1 vccd1 _07387_/A sky130_fd_sc_hd__or3_1
X_09125_ _09125_/A _09125_/B vssd1 vssd1 vccd1 vccd1 _09134_/A sky130_fd_sc_hd__nor2_1
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06337_ _06337_/A vssd1 vssd1 vccd1 vccd1 _06337_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__13977__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09056_ _13970_/A vssd1 vssd1 vccd1 vccd1 _09056_/X sky130_fd_sc_hd__buf_2
X_06268_ _11457_/A vssd1 vssd1 vccd1 vccd1 _10693_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11497__A _12084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09908__A1 _09186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ _08022_/A vssd1 vssd1 vccd1 vccd1 _08020_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_150_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_3_0_clk_A clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09958_ _13594_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _09958_/X sky130_fd_sc_hd__or2_1
XFILLER_106_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08909_ _12810_/Q vssd1 vssd1 vccd1 vccd1 _11518_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09889_ _09915_/B vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11920_ _11920_/A _11920_/B _11920_/C _11920_/D vssd1 vssd1 vccd1 vccd1 _11921_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_58_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _12888_/Q _14032_/A _11861_/S vssd1 vssd1 vccd1 vccd1 _11852_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _12628_/Q vssd1 vssd1 vccd1 vccd1 _10864_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11782_ _12862_/Q _13367_/A vssd1 vssd1 vccd1 vccd1 _11785_/B sky130_fd_sc_hd__xor2_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13521_ _13521_/A _07569_/X vssd1 vssd1 vccd1 vccd1 _14033_/Z sky130_fd_sc_hd__ebufn_8
X_10733_ _10288_/X _10703_/S _10732_/X _10711_/X vssd1 vssd1 vccd1 vccd1 _12613_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13452_ _13452_/A _07747_/X vssd1 vssd1 vccd1 vccd1 _13996_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10664_ _10662_/X _10655_/X _10663_/X _10650_/X vssd1 vssd1 vccd1 vccd1 _12591_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08046__A _08072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12403_ _12404_/CLK _12403_/D vssd1 vssd1 vccd1 vccd1 _13531_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13383_ _13383_/A _08334_/X vssd1 vssd1 vccd1 vccd1 _14119_/Z sky130_fd_sc_hd__ebufn_8
X_10595_ _13722_/A _12578_/Q _10601_/S vssd1 vssd1 vccd1 vccd1 _10596_/B sky130_fd_sc_hd__mux2_1
XFILLER_126_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12334_ _12334_/CLK _12334_/D vssd1 vssd1 vccd1 vccd1 _13464_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12265_ _12912_/CLK _12265_/D vssd1 vssd1 vccd1 vccd1 _12265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14004_ _14004_/A _07952_/X vssd1 vssd1 vccd1 vccd1 _14100_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_107_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11216_ _11254_/S vssd1 vssd1 vccd1 vccd1 _11231_/S sky130_fd_sc_hd__clkbuf_2
X_13264__420 vssd1 vssd1 vccd1 vccd1 _13264__420/HI _13955_/A sky130_fd_sc_hd__conb_1
X_12196_ _12208_/B vssd1 vssd1 vccd1 vccd1 _12206_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_122_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11147_ _12698_/Q _13939_/A vssd1 vssd1 vccd1 vccd1 _11148_/D sky130_fd_sc_hd__xor2_1
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output58_A _13759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11078_ _11078_/A _11078_/B vssd1 vssd1 vccd1 vccd1 _11079_/A sky130_fd_sc_hd__and2_1
X_13305__461 vssd1 vssd1 vccd1 vccd1 _13305__461/HI _14026_/A sky130_fd_sc_hd__conb_1
XFILLER_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10029_ _10029_/A _10029_/B _10029_/C _10029_/D vssd1 vssd1 vccd1 vccd1 _10030_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_48_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13719_ _13719_/A _07042_/X vssd1 vssd1 vccd1 vccd1 _14103_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_32_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07240_ _07240_/A vssd1 vssd1 vccd1 vccd1 _07240_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12198__A1 _10659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07171_ _07180_/A _07177_/B _07173_/C vssd1 vssd1 vccd1 vccd1 _07172_/A sky130_fd_sc_hd__or3_1
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07795__A _08064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09812_ _09812_/A vssd1 vssd1 vccd1 vccd1 _12379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater80_A peripheralBus_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09515__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ _11285_/B _09875_/B _11156_/C vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__nor3_4
X_06955_ _06955_/A vssd1 vssd1 vccd1 vccd1 _06965_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_100_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09674_ _09686_/A _09674_/B vssd1 vssd1 vccd1 vccd1 _09675_/A sky130_fd_sc_hd__and2_1
XFILLER_54_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08421__S0 _08373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06886_ _06900_/A vssd1 vssd1 vccd1 vccd1 _06898_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _12430_/Q vssd1 vssd1 vccd1 vccd1 _10029_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _13584_/A vssd1 vssd1 vccd1 vccd1 _08556_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06874__A _07090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ _07507_/A vssd1 vssd1 vccd1 vccd1 _07517_/B sky130_fd_sc_hd__clkbuf_1
X_08487_ _12266_/Q vssd1 vssd1 vccd1 vccd1 _09362_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10396__A _10423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07438_ _07442_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07439_/A sky130_fd_sc_hd__or2_1
XFILLER_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11004__B _13936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07369_ _07369_/A _07377_/B _07374_/C vssd1 vssd1 vccd1 vccd1 _07370_/A sky130_fd_sc_hd__or3_1
XANTENNA__08488__S0 _08368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09108_ _11443_/A vssd1 vssd1 vccd1 vccd1 _12155_/A sky130_fd_sc_hd__clkbuf_2
X_10380_ _11156_/B _11412_/C _10693_/C vssd1 vssd1 vccd1 vccd1 _10423_/B sky130_fd_sc_hd__nor3_4
X_13248__404 vssd1 vssd1 vccd1 vccd1 _13248__404/HI _13919_/A sky130_fd_sc_hd__conb_1
XFILLER_124_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _10938_/D vssd1 vssd1 vccd1 vccd1 _13942_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_136_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12050_ _12050_/A _12050_/B _12050_/C _12050_/D vssd1 vssd1 vccd1 vccd1 _12056_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_151_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11001_ _12674_/Q _13948_/A vssd1 vssd1 vccd1 vccd1 _11001_/X sky130_fd_sc_hd__or2_1
XFILLER_89_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12952_ _12952_/CLK _12952_/D vssd1 vssd1 vccd1 vccd1 _14078_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11903_ _12900_/Q _13372_/A vssd1 vssd1 vccd1 vccd1 _11905_/C sky130_fd_sc_hd__xor2_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12883_ _12886_/CLK _12883_/D vssd1 vssd1 vccd1 vccd1 _14011_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11690__A _11703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _11834_/A _11834_/B vssd1 vssd1 vccd1 vccd1 _11835_/A sky130_fd_sc_hd__and2_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09160__A _11170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _11765_/A vssd1 vssd1 vccd1 vccd1 _12869_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10737__C _10737_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _13504_/A _07612_/X vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__ebufn_8
X_10716_ _13974_/Z _13782_/A _10723_/S vssd1 vssd1 vccd1 vccd1 _10717_/B sky130_fd_sc_hd__mux2_1
XFILLER_147_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11696_ _11699_/B vssd1 vssd1 vccd1 vccd1 _11696_/Y sky130_fd_sc_hd__inv_2
X_13435_ _13435_/A _07791_/X vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__ebufn_8
X_10647_ _10645_/X _10638_/X _10646_/X _10550_/X vssd1 vssd1 vccd1 vccd1 _12586_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13366_ _13366_/A _08294_/X vssd1 vssd1 vccd1 vccd1 _14102_/Z sky130_fd_sc_hd__ebufn_8
X_10578_ _13717_/A _12573_/Q _10584_/S vssd1 vssd1 vccd1 vccd1 _10579_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12317_ _12320_/CLK _12317_/D vssd1 vssd1 vccd1 vccd1 _12317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12248_ _12251_/CLK _12248_/D vssd1 vssd1 vccd1 vccd1 _12248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12179_ _13375_/A _12178_/Y _11711_/B _09404_/A _13401_/A vssd1 vssd1 vccd1 vccd1
+ _12969_/D sky130_fd_sc_hd__o2111a_1
XFILLER_68_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06740_ _06753_/A vssd1 vssd1 vccd1 vccd1 _06751_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_83_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06671_ _06673_/A _06678_/B _06678_/C vssd1 vssd1 vccd1 vccd1 _06672_/A sky130_fd_sc_hd__or3_1
XFILLER_36_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08410_ _12259_/Q vssd1 vssd1 vccd1 vccd1 _09343_/C sky130_fd_sc_hd__clkbuf_2
X_09390_ _09390_/A vssd1 vssd1 vccd1 vccd1 _12273_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__06694__A _06694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10418__A1 _10285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08341_ _08347_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08342_/A sky130_fd_sc_hd__or2_1
X_08272_ _08276_/A _08274_/B _08276_/C vssd1 vssd1 vccd1 vccd1 _08273_/A sky130_fd_sc_hd__or3_1
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07223_ _07281_/A vssd1 vssd1 vccd1 vccd1 _07239_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater90 _13995_/Z vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__buf_12
XFILLER_118_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07154_ _07533_/A vssd1 vssd1 vccd1 vccd1 _07208_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__07956__C _07993_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07085_ _07085_/A vssd1 vssd1 vccd1 vccd1 _07085_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08133__B _08189_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input1_A peripheralBus_address[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07987_ _07987_/A vssd1 vssd1 vccd1 vccd1 _07987_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09726_ _12343_/Q _13553_/A vssd1 vssd1 vccd1 vccd1 _09730_/A sky130_fd_sc_hd__xor2_1
X_06938_ _06974_/A vssd1 vssd1 vccd1 vccd1 _06948_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09657_ _13594_/A _09791_/B vssd1 vssd1 vccd1 vccd1 _09711_/S sky130_fd_sc_hd__and2_2
X_06869_ _06869_/A vssd1 vssd1 vccd1 vccd1 _06869_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _12433_/Q vssd1 vssd1 vccd1 vccd1 _10021_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _12319_/Q _13562_/A vssd1 vssd1 vccd1 vccd1 _09588_/Y sky130_fd_sc_hd__nor2_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08536_/X _08538_/X _09162_/A vssd1 vssd1 vccd1 vccd1 _11708_/C sky130_fd_sc_hd__mux2_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11550_ _11558_/C _11604_/B _11550_/C vssd1 vssd1 vccd1 vccd1 _11551_/A sky130_fd_sc_hd__and3b_1
XFILLER_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ _12538_/Q _13747_/A vssd1 vssd1 vccd1 vccd1 _10504_/B sky130_fd_sc_hd__xor2_1
X_11481_ _11481_/A _11481_/B vssd1 vssd1 vccd1 vccd1 _11482_/A sky130_fd_sc_hd__or2_1
X_10432_ _10432_/A vssd1 vssd1 vccd1 vccd1 _12534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08324__A _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ _12516_/Q _13758_/A vssd1 vssd1 vccd1 vccd1 _10367_/A sky130_fd_sc_hd__xor2_1
XFILLER_136_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12102_ _10552_/A _12088_/A _12101_/X _12097_/X vssd1 vssd1 vccd1 vccd1 _12952_/D
+ sky130_fd_sc_hd__o211a_1
X_10294_ _09120_/X _10278_/A _10293_/X _10283_/X vssd1 vssd1 vccd1 vccd1 _12500_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _12935_/Q _14078_/A _12033_/S vssd1 vssd1 vccd1 vccd1 _12034_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_0_0_clk_A clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09155__A _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A _12917_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13984_ _13984_/A _06330_/X vssd1 vssd1 vccd1 vccd1 _14112_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12935_ _12935_/CLK _12935_/D vssd1 vssd1 vccd1 vccd1 _12935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12866_ _12886_/CLK _12866_/D vssd1 vssd1 vccd1 vccd1 _12866_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07403__A _07403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _11817_/A vssd1 vssd1 vccd1 vccd1 _12878_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12811_/CLK _12797_/D vssd1 vssd1 vccd1 vccd1 _13971_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _11757_/A _11748_/B vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__and2_1
X_11679_ _11679_/A _11680_/C vssd1 vssd1 vccd1 vccd1 _12846_/D sky130_fd_sc_hd__nor2_1
X_13418_ _13418_/A _07844_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__10483__B _13752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07910_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07921_/A sky130_fd_sc_hd__clkbuf_1
X_08890_ _08884_/X _08889_/X _08890_/S vssd1 vssd1 vccd1 vccd1 _10165_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10703__S _10703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08624__S0 _08602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07841_ _07841_/A vssd1 vssd1 vccd1 vccd1 _07841_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12984__140 vssd1 vssd1 vccd1 vccd1 _12984__140/HI _13381_/A sky130_fd_sc_hd__conb_1
XFILLER_96_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07772_ _07782_/A _07779_/B _07774_/C vssd1 vssd1 vccd1 vccd1 _07773_/A sky130_fd_sc_hd__or3_1
XFILLER_17_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09511_ _09638_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09511_/X sky130_fd_sc_hd__or2_1
X_06723_ _06733_/A _06738_/B _07863_/B vssd1 vssd1 vccd1 vccd1 _06724_/A sky130_fd_sc_hd__or3_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09442_ _13434_/A _12286_/Q _09448_/S vssd1 vssd1 vccd1 vccd1 _09443_/B sky130_fd_sc_hd__mux2_1
X_06654_ _08184_/B vssd1 vssd1 vccd1 vccd1 _06664_/C sky130_fd_sc_hd__clkbuf_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _09373_/A vssd1 vssd1 vccd1 vccd1 _12268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06585_ _06585_/A vssd1 vssd1 vccd1 vccd1 _06585_/X sky130_fd_sc_hd__clkbuf_1
X_08324_ _08324_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08325_/A sky130_fd_sc_hd__or2_1
XFILLER_32_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08255_ _08264_/A _08261_/B _08264_/C vssd1 vssd1 vccd1 vccd1 _08256_/A sky130_fd_sc_hd__or3_1
XFILLER_138_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10674__A _10686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07206_ _07206_/A _07216_/B _07213_/C vssd1 vssd1 vccd1 vccd1 _07207_/A sky130_fd_sc_hd__or3_1
X_08186_ _08186_/A vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__buf_4
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07137_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07152_/A sky130_fd_sc_hd__clkbuf_1
X_13210__366 vssd1 vssd1 vccd1 vccd1 _13210__366/HI _13833_/A sky130_fd_sc_hd__conb_1
XFILLER_106_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07068_ _08177_/A vssd1 vssd1 vccd1 vccd1 _07079_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_160_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11827__A0 _14009_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _09800_/A _09709_/B vssd1 vssd1 vccd1 vccd1 _09710_/A sky130_fd_sc_hd__and2_1
X_10981_ _10981_/A vssd1 vssd1 vccd1 vccd1 _12671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13104__260 vssd1 vssd1 vccd1 vccd1 _13104__260/HI _13613_/A sky130_fd_sc_hd__conb_1
XFILLER_71_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12720_ _12724_/CLK _12720_/D vssd1 vssd1 vccd1 vccd1 _13848_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08319__A _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12651_ _12652_/CLK _12651_/D vssd1 vssd1 vccd1 vccd1 _12651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11602_ _11641_/C _11631_/B _11602_/C _11642_/A vssd1 vssd1 vccd1 vccd1 _11610_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_30_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12582_ _12597_/CLK _12582_/D vssd1 vssd1 vccd1 vccd1 _12582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11533_ _11533_/A _11533_/B vssd1 vssd1 vccd1 vccd1 _12813_/D sky130_fd_sc_hd__nor2_1
XFILLER_156_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11399__B _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11464_ _12084_/A vssd1 vssd1 vccd1 vccd1 _11464_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__08054__A _08067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13895__A _13895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10415_ _13658_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10415_/X sky130_fd_sc_hd__or2_1
X_11395_ _11395_/A _11395_/B _11395_/C _11395_/D vssd1 vssd1 vccd1 vccd1 _11406_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_152_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07893__A _07920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ _10349_/A _10346_/B vssd1 vssd1 vccd1 vccd1 _10347_/A sky130_fd_sc_hd__and2_1
XFILLER_152_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10277_ _09773_/X _10264_/X _10276_/X _10270_/X vssd1 vssd1 vccd1 vccd1 _12494_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_repeater111_A _14082_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08606__S0 _08575_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12016_ _12033_/S vssd1 vssd1 vccd1 vccd1 _12029_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output40_A _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09613__A _09640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13967_ _13967_/A _07823_/X vssd1 vssd1 vccd1 vccd1 _14063_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11294__A1 _10645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12918_ _12918_/CLK _12918_/D vssd1 vssd1 vccd1 vccd1 _14045_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13898_ _13898_/A _06562_/X vssd1 vssd1 vccd1 vccd1 _13994_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_34_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07133__A _08035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _12850_/CLK _12849_/D vssd1 vssd1 vccd1 vccd1 _12849_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11046__A1 _10659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13153__309 vssd1 vssd1 vccd1 vccd1 _13153__309/HI _13710_/A sky130_fd_sc_hd__conb_1
X_06370_ _06370_/A vssd1 vssd1 vccd1 vccd1 _06370_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10254__C1 _09959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ _08040_/A vssd1 vssd1 vccd1 vccd1 _08040_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09991_ _09997_/C _09993_/C _09987_/X vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10941__B _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13047__203 vssd1 vssd1 vccd1 vccd1 _13047__203/HI _13506_/A sky130_fd_sc_hd__conb_1
XFILLER_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08942_ _09068_/A vssd1 vssd1 vccd1 vccd1 _08942_/X sky130_fd_sc_hd__buf_2
XFILLER_97_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08873_ _08793_/X _08795_/X _08846_/X _08872_/X _08826_/X _08859_/X vssd1 vssd1 vccd1
+ vccd1 _08873_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07824_ _11789_/A _11789_/B _07824_/C vssd1 vssd1 vccd1 vccd1 _09125_/B sky130_fd_sc_hd__or3_4
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11809__A0 _14068_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__B _13365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07755_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07766_/B sky130_fd_sc_hd__clkbuf_1
X_06706_ _06714_/A _06706_/B _06706_/C vssd1 vssd1 vccd1 vccd1 _06707_/A sky130_fd_sc_hd__or3_1
X_07686_ _07686_/A _07696_/B _07691_/C vssd1 vssd1 vccd1 vccd1 _07687_/A sky130_fd_sc_hd__or3_1
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ _13429_/A _12281_/Q _09431_/S vssd1 vssd1 vccd1 vccd1 _09426_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06637_ _06637_/A _09096_/B vssd1 vssd1 vccd1 vccd1 _06725_/B sky130_fd_sc_hd__or2_1
XANTENNA__11037__A1 _10648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _09356_/A _09358_/B vssd1 vssd1 vccd1 vccd1 _12264_/D sky130_fd_sc_hd__nor2_1
XFILLER_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06568_ _06568_/A vssd1 vssd1 vccd1 vccd1 _06568_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10245__C1 _09959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08307_ _08312_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08308_/A sky130_fd_sc_hd__or2_1
XFILLER_138_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09287_ _09292_/C _09389_/A _09287_/C vssd1 vssd1 vccd1 vccd1 _09288_/A sky130_fd_sc_hd__and3b_1
X_06499_ _06507_/A _06499_/B _06499_/C vssd1 vssd1 vccd1 vccd1 _06500_/A sky130_fd_sc_hd__or3_1
X_08238_ _08238_/A _08248_/B _08238_/C vssd1 vssd1 vccd1 vccd1 _08239_/A sky130_fd_sc_hd__or3_1
XFILLER_138_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11012__B _13942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08169_ _08169_/A vssd1 vssd1 vccd1 vccd1 _08169_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10200_ _10220_/S vssd1 vssd1 vccd1 vccd1 _10214_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11180_ _11195_/A vssd1 vssd1 vccd1 vccd1 _11180_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10131_ _10114_/X _10137_/D _10049_/A vssd1 vssd1 vccd1 vccd1 _10131_/X sky130_fd_sc_hd__a21bo_1
XFILLER_161_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10062_ _10064_/B _10062_/B _10062_/C vssd1 vssd1 vccd1 vccd1 _10063_/A sky130_fd_sc_hd__and3b_1
XFILLER_125_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11682__B _11682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ _13821_/A _06776_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[14] sky130_fd_sc_hd__ebufn_8
XFILLER_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13752_ _13752_/A _06961_/X vssd1 vssd1 vccd1 vccd1 _14072_/Z sky130_fd_sc_hd__ebufn_8
X_10964_ _10964_/A vssd1 vssd1 vccd1 vccd1 _12666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08049__A _11283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ _12704_/CLK _12703_/D vssd1 vssd1 vccd1 vccd1 _12703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13683_ _13683_/A _07139_/X vssd1 vssd1 vccd1 vccd1 _14099_/Z sky130_fd_sc_hd__ebufn_8
X_10895_ _10895_/A _10895_/B _10895_/C vssd1 vssd1 vccd1 vccd1 _12648_/D sky130_fd_sc_hd__nor3_1
XFILLER_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12634_ _12634_/CLK _12634_/D vssd1 vssd1 vccd1 vccd1 _12634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12565_ _12565_/CLK _12565_/D vssd1 vssd1 vccd1 vccd1 _13693_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10745__C _10917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ _11518_/B _11514_/B _11515_/X vssd1 vssd1 vccd1 vccd1 _11517_/B sky130_fd_sc_hd__o21ai_1
XFILLER_156_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ _12522_/CLK _12496_/D vssd1 vssd1 vccd1 vccd1 _13626_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11447_ _11061_/X _11438_/X _11446_/X _11444_/X vssd1 vssd1 vccd1 vccd1 _12789_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11200__A1 _10552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11378_ _11378_/A vssd1 vssd1 vccd1 vccd1 _12774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _10332_/A _10329_/B vssd1 vssd1 vccd1 vccd1 _10330_/A sky130_fd_sc_hd__and2_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _14097_/A _08203_/X vssd1 vssd1 vccd1 vccd1 _14097_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06967__A _06967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__A _13391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09004__S0 _08946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07540_ _07553_/A vssd1 vssd1 vccd1 vccd1 _07551_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_80_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07471_ _07478_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07472_/A sky130_fd_sc_hd__or2_1
XFILLER_34_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09210_ _09210_/A _09210_/B _12229_/Q _12228_/Q vssd1 vssd1 vccd1 vccd1 _09318_/A
+ sky130_fd_sc_hd__and4_1
X_06422_ _06422_/A vssd1 vssd1 vccd1 vccd1 _06422_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_95_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ _12155_/A vssd1 vssd1 vccd1 vccd1 _09141_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06353_ _06359_/A _06362_/B _06362_/C vssd1 vssd1 vccd1 vccd1 _06354_/A sky130_fd_sc_hd__or3_1
X_09072_ _10941_/A vssd1 vssd1 vccd1 vccd1 _13947_/A sky130_fd_sc_hd__buf_6
XANTENNA__07310__B _07317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06284_ _06694_/A vssd1 vssd1 vccd1 vccd1 _06547_/A sky130_fd_sc_hd__buf_2
XFILLER_107_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08023_ _08025_/A _08033_/B _08030_/C vssd1 vssd1 vccd1 vccd1 _08024_/A sky130_fd_sc_hd__or3_1
XANTENNA__10952__A _10952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__S0 _08807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11767__B _13370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _09977_/A vssd1 vssd1 vccd1 vccd1 _10157_/B sky130_fd_sc_hd__buf_2
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13281__437 vssd1 vssd1 vccd1 vccd1 _13281__437/HI _13986_/A sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_33_clk_A _12759_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08925_ _13971_/A vssd1 vssd1 vccd1 vccd1 _08925_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08856_ _08818_/X _08822_/X _08825_/X _08855_/X _08810_/X _08812_/X vssd1 vssd1 vccd1
+ vccd1 _08856_/X sky130_fd_sc_hd__mux4_1
X_13322__478 vssd1 vssd1 vccd1 vccd1 _13322__478/HI _14059_/A sky130_fd_sc_hd__conb_1
XFILLER_84_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07807_ _07807_/A vssd1 vssd1 vccd1 vccd1 _07807_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08787_ _12628_/Q _10864_/A _10874_/C _12631_/Q _08785_/X _08786_/X vssd1 vssd1 vccd1
+ vccd1 _08787_/X sky130_fd_sc_hd__mux4_2
XFILLER_72_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_48_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ _07738_/A vssd1 vssd1 vccd1 vccd1 _07738_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11007__B _13945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07669_ _07672_/A _07669_/B _07678_/C vssd1 vssd1 vccd1 vccd1 _07670_/A sky130_fd_sc_hd__or3_1
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13175__331 vssd1 vssd1 vccd1 vccd1 _13175__331/HI _13768_/A sky130_fd_sc_hd__conb_1
X_09408_ _13424_/A _12276_/Q _09414_/S vssd1 vssd1 vccd1 vccd1 _09409_/B sky130_fd_sc_hd__mux2_1
XFILLER_111_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ _10285_/X _10673_/X _10679_/X _10668_/X vssd1 vssd1 vccd1 vccd1 _12596_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09339_ _09379_/A _09363_/A _09346_/C vssd1 vssd1 vccd1 vccd1 _09341_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_106_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13216__372 vssd1 vssd1 vccd1 vccd1 _13216__372/HI _13855_/A sky130_fd_sc_hd__conb_1
XANTENNA__07220__B _07231_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ _12367_/CLK _12350_/D vssd1 vssd1 vccd1 vccd1 _12350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11301_ _13876_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11301_/X sky130_fd_sc_hd__or2_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12281_ _12289_/CLK _12281_/D vssd1 vssd1 vccd1 vccd1 _12281_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08809__S0 _08807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11232_ _11239_/A _11232_/B vssd1 vssd1 vccd1 vccd1 _11233_/A sky130_fd_sc_hd__and2_1
X_14020_ _14020_/A _08106_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[21] sky130_fd_sc_hd__ebufn_8
XFILLER_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ _13841_/A _11168_/B vssd1 vssd1 vccd1 vccd1 _11163_/X sky130_fd_sc_hd__or2_1
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10114_ _10126_/D vssd1 vssd1 vccd1 vccd1 _10114_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11094_ _13845_/A _12700_/Q _11101_/S vssd1 vssd1 vccd1 vccd1 _11095_/B sky130_fd_sc_hd__mux2_1
XFILLER_95_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10045_ _10052_/C _10052_/D _10045_/C vssd1 vssd1 vccd1 vccd1 _10045_/X sky130_fd_sc_hd__and3_1
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_10_0_clk_A clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13804_ _13804_/A _06827_/X vssd1 vssd1 vccd1 vccd1 _14028_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11996_ _11996_/A _11996_/B vssd1 vssd1 vccd1 vccd1 _11997_/A sky130_fd_sc_hd__and2_1
XFILLER_90_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13735_ _13735_/A _07004_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[24] sky130_fd_sc_hd__ebufn_8
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10947_ _10947_/A vssd1 vssd1 vccd1 vccd1 _12661_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13666_ _13666_/A _07184_/X vssd1 vssd1 vccd1 vccd1 _13666_/Z sky130_fd_sc_hd__ebufn_8
X_10878_ _10881_/A _10878_/B _10880_/D vssd1 vssd1 vccd1 vccd1 _10878_/Y sky130_fd_sc_hd__nand3_1
X_12617_ _12617_/CLK _12617_/D vssd1 vssd1 vccd1 vccd1 _12617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_clk/X
+ sky130_fd_sc_hd__clkbuf_2
X_13597_ _13597_/A _07373_/X vssd1 vssd1 vccd1 vccd1 _14109_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_157_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12548_ _12599_/CLK _12548_/D vssd1 vssd1 vccd1 vccd1 _12548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12479_ _12522_/CLK _12479_/D vssd1 vssd1 vccd1 vccd1 _12479_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09917__A2 _09902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10491__B _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _06971_/A vssd1 vssd1 vccd1 vccd1 _06971_/X sky130_fd_sc_hd__clkbuf_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _10148_/C _10148_/B _10148_/A _10149_/A _09929_/A _08709_/X vssd1 vssd1 vccd1
+ vccd1 _08710_/X sky130_fd_sc_hd__mux4_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _09836_/A vssd1 vssd1 vccd1 vccd1 _09705_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08641_ _12448_/Q vssd1 vssd1 vccd1 vccd1 _10099_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08572_ _12425_/Q vssd1 vssd1 vccd1 vccd1 _09997_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_13159__315 vssd1 vssd1 vccd1 vccd1 _13159__315/HI _13732_/A sky130_fd_sc_hd__conb_1
XFILLER_35_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07523_ _07523_/A vssd1 vssd1 vccd1 vccd1 _07523_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07454_ _07454_/A _07459_/B vssd1 vssd1 vccd1 vccd1 _07455_/A sky130_fd_sc_hd__or2_1
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07321__A _09484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06405_ _07861_/A vssd1 vssd1 vccd1 vccd1 _06416_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07385_ _07964_/A vssd1 vssd1 vccd1 vccd1 _07396_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09124_ _11153_/A vssd1 vssd1 vccd1 vccd1 _09124_/X sky130_fd_sc_hd__buf_4
X_06336_ _06346_/A _06336_/B _06336_/C vssd1 vssd1 vccd1 vccd1 _06337_/A sky130_fd_sc_hd__or3_1
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _10940_/C vssd1 vssd1 vccd1 vccd1 _13945_/A sky130_fd_sc_hd__buf_6
XFILLER_135_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06267_ input18/X _09102_/A _06548_/C _09096_/C vssd1 vssd1 vccd1 vccd1 _11457_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA__10682__A _11039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08006_ _08006_/A vssd1 vssd1 vccd1 vccd1 _08006_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07991__A _07997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09957_ _09182_/X _09921_/X _09956_/X _09916_/X vssd1 vssd1 vccd1 vccd1 _12417_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08908_ _10165_/D vssd1 vssd1 vccd1 vccd1 _13758_/A sky130_fd_sc_hd__buf_4
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09902_/A vssd1 vssd1 vccd1 vccd1 _09888_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08839_ _08764_/X _08768_/X _08765_/X _08771_/X _08837_/X _08838_/X vssd1 vssd1 vccd1
+ vccd1 _08839_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08895__A2 _08866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _11850_/A vssd1 vssd1 vccd1 vccd1 _12887_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _10801_/A _10801_/B vssd1 vssd1 vccd1 vccd1 _12627_/D sky130_fd_sc_hd__nor2_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11781_ _12859_/Q _13364_/A vssd1 vssd1 vccd1 vccd1 _11785_/A sky130_fd_sc_hd__xor2_1
X_13520_ _13520_/A _07571_/X vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10732_ _13788_/A _10732_/B vssd1 vssd1 vccd1 vccd1 _10732_/X sky130_fd_sc_hd__or2_1
XFILLER_41_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13451_ _13451_/A _07749_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
X_10663_ _13718_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10663_/X sky130_fd_sc_hd__or2_1
XFILLER_139_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12402_ _12404_/CLK _12402_/D vssd1 vssd1 vccd1 vccd1 _13530_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10594_ _10594_/A vssd1 vssd1 vccd1 vccd1 _12577_/D sky130_fd_sc_hd__clkbuf_1
X_13382_ _13382_/A _08332_/X vssd1 vssd1 vccd1 vccd1 _14086_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12333_ _12334_/CLK _12333_/D vssd1 vssd1 vccd1 vccd1 _13463_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12264_ _12264_/CLK _12264_/D vssd1 vssd1 vccd1 vccd1 _12264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14003_ _14003_/A _07972_/X vssd1 vssd1 vccd1 vccd1 _14067_/Z sky130_fd_sc_hd__ebufn_8
X_11215_ _11215_/A vssd1 vssd1 vccd1 vccd1 _12730_/D sky130_fd_sc_hd__clkbuf_1
X_12195_ _12195_/A vssd1 vssd1 vccd1 vccd1 _12195_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput50 _13954_/A vssd1 vssd1 vccd1 vccd1 pwm_out[15] sky130_fd_sc_hd__buf_2
X_11146_ _12702_/Q _13943_/A vssd1 vssd1 vccd1 vccd1 _11148_/C sky130_fd_sc_hd__xor2_1
XFILLER_150_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11077_ _13840_/A _12695_/Q _11151_/B vssd1 vssd1 vccd1 vccd1 _11078_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09605__B _13559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09532__A0 _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10028_ _10029_/A _10024_/X _09978_/X vssd1 vssd1 vccd1 vccd1 _10033_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__07406__A _07406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06310__A _11457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09621__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11979_ _11979_/A vssd1 vssd1 vccd1 vccd1 _12919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13718_ _13718_/A _07044_/X vssd1 vssd1 vccd1 vccd1 _13974_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__08237__A _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10486__B _10614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13649_ _13649_/A _07229_/X vssd1 vssd1 vccd1 vccd1 _14097_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07170_ _07170_/A vssd1 vssd1 vccd1 vccd1 _07170_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09811_ _09817_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__and2_1
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09742_ _10250_/A vssd1 vssd1 vccd1 vccd1 _11156_/C sky130_fd_sc_hd__buf_6
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06954_ _06954_/A vssd1 vssd1 vccd1 vccd1 _06954_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater73_A peripheralBus_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _13491_/A _12345_/Q _09685_/S vssd1 vssd1 vccd1 vccd1 _09674_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06885_ _06885_/A vssd1 vssd1 vccd1 vccd1 _06885_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08421__S1 _08374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _09981_/A _09997_/D _09997_/C _09997_/B _08602_/X _08603_/X vssd1 vssd1 vccd1
+ vccd1 _08624_/X sky130_fd_sc_hd__mux4_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09531__A _09582_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _12425_/Q _12426_/Q _12427_/Q _12428_/Q _08553_/X _08554_/X vssd1 vssd1 vccd1
+ vccd1 _08555_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07506_ _07519_/A vssd1 vssd1 vccd1 vccd1 _07517_/A sky130_fd_sc_hd__clkbuf_1
X_08486_ _08439_/X _08447_/X _08443_/X _08452_/X _08470_/X _09152_/A vssd1 vssd1 vccd1
+ vccd1 _08486_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07437_ _08131_/C vssd1 vssd1 vccd1 vccd1 _07447_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07986__A _07997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07368_ _07368_/A vssd1 vssd1 vccd1 vccd1 _07368_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08488__S1 _08370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09107_ _09967_/B vssd1 vssd1 vccd1 vccd1 _11443_/A sky130_fd_sc_hd__buf_4
X_06319_ _06319_/A vssd1 vssd1 vccd1 vccd1 _06319_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_111_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _12290_/CLK sky130_fd_sc_hd__clkbuf_16
X_07299_ _07299_/A vssd1 vssd1 vccd1 vccd1 _07299_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13287__443 vssd1 vssd1 vccd1 vccd1 _13287__443/HI _13992_/A sky130_fd_sc_hd__conb_1
X_09038_ _09031_/X _09037_/X _09071_/S vssd1 vssd1 vccd1 vccd1 _10938_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11020__B _13939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11000_ _12670_/Q _13944_/A vssd1 vssd1 vccd1 vccd1 _11000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13328__484 vssd1 vssd1 vccd1 vccd1 _13328__484/HI _14081_/A sky130_fd_sc_hd__conb_1
XFILLER_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ _12952_/CLK _12951_/D vssd1 vssd1 vccd1 vccd1 _14077_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11902_ _12898_/Q _13370_/A vssd1 vssd1 vccd1 vccd1 _11905_/B sky130_fd_sc_hd__xor2_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12882_ _12886_/CLK _12882_/D vssd1 vssd1 vccd1 vccd1 _14010_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09441__A _11408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11833_ _13979_/Z _14011_/A _11840_/S vssd1 vssd1 vccd1 vccd1 _11834_/B sky130_fd_sc_hd__mux2_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10587__A _10971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11799_/A _11764_/B vssd1 vssd1 vccd1 vccd1 _11765_/A sky130_fd_sc_hd__and2_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13503_ _13503_/A _07614_/X vssd1 vssd1 vccd1 vccd1 _14111_/Z sky130_fd_sc_hd__ebufn_8
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10715_/A vssd1 vssd1 vccd1 vccd1 _12606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11695_ _12851_/Q _11695_/B _11695_/C vssd1 vssd1 vccd1 vccd1 _11699_/B sky130_fd_sc_hd__and3_1
XFILLER_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13434_ _13434_/A _07793_/X vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__07896__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10646_ _13713_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10646_/X sky130_fd_sc_hd__or2_1
XFILLER_155_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13365_ _13365_/A _08292_/X vssd1 vssd1 vccd1 vccd1 _14037_/Z sky130_fd_sc_hd__ebufn_8
X_10577_ _10577_/A vssd1 vssd1 vccd1 vccd1 _12572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12316_ _12320_/CLK _12316_/D vssd1 vssd1 vccd1 vccd1 _12316_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06305__A _11457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12247_ _12251_/CLK _12247_/D vssd1 vssd1 vccd1 vccd1 _12247_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09616__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12178_ _12178_/A _12178_/B vssd1 vssd1 vccd1 vccd1 _12178_/Y sky130_fd_sc_hd__nor2_1
X_11129_ _12707_/Q _11386_/B vssd1 vssd1 vccd1 vccd1 _11129_/X sky130_fd_sc_hd__and2_1
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13080__236 vssd1 vssd1 vccd1 vccd1 _13080__236/HI _13575_/A sky130_fd_sc_hd__conb_1
XFILLER_83_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11881__A _11898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06670_ _06670_/A vssd1 vssd1 vccd1 vccd1 _06670_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06975__A _07417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13121__277 vssd1 vssd1 vccd1 vccd1 _13121__277/HI _13646_/A sky130_fd_sc_hd__conb_1
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08340_ _08340_/A vssd1 vssd1 vccd1 vccd1 _08340_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08271_ _08271_/A vssd1 vssd1 vccd1 vccd1 _08271_/X sky130_fd_sc_hd__clkbuf_1
X_07222_ _07533_/A vssd1 vssd1 vccd1 vccd1 _07281_/A sky130_fd_sc_hd__clkbuf_2
Xrepeater80 peripheralBus_data[3] vssd1 vssd1 vccd1 vccd1 _14034_/Z sky130_fd_sc_hd__buf_12
Xrepeater91 peripheralBus_data[28] vssd1 vssd1 vccd1 vccd1 _13995_/Z sky130_fd_sc_hd__buf_12
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07153_ _07153_/A vssd1 vssd1 vccd1 vccd1 _07153_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13015__171 vssd1 vssd1 vccd1 vccd1 _13015__171/HI _13442_/A sky130_fd_sc_hd__conb_1
X_07084_ _07094_/A _07091_/B _07088_/C vssd1 vssd1 vccd1 vccd1 _07085_/A sky130_fd_sc_hd__or3_1
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09526__A _10552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09245__B _09389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07986_ _07997_/A _08062_/B _08002_/C vssd1 vssd1 vccd1 vccd1 _07987_/A sky130_fd_sc_hd__or3_1
XFILLER_86_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07046__A _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09725_ _09725_/A _09725_/B _09725_/C _09725_/D vssd1 vssd1 vccd1 vccd1 _09736_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10106__A1 _09982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06937_ _06937_/A vssd1 vssd1 vccd1 vccd1 _06937_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09656_ _13470_/A _09640_/A _09655_/X _09649_/X vssd1 vssd1 vccd1 vccd1 _12340_/D
+ sky130_fd_sc_hd__o211a_1
X_06868_ _06877_/A _06870_/B _06870_/C vssd1 vssd1 vccd1 vccd1 _06869_/A sky130_fd_sc_hd__or3_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08607_ _12431_/Q vssd1 vssd1 vccd1 vccd1 _10021_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _12319_/Q _09848_/B vssd1 vssd1 vccd1 vccd1 _09587_/X sky130_fd_sc_hd__and2_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ _06801_/A _06806_/B _06806_/C vssd1 vssd1 vccd1 vccd1 _06800_/A sky130_fd_sc_hd__or3_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08431_/X _08482_/X _08507_/X _08537_/X _08511_/X _09157_/A vssd1 vssd1 vccd1
+ vccd1 _08538_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10200__A _10220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11015__B _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08469_ _12260_/Q _12261_/Q _12262_/Q _12263_/Q _08404_/X _08405_/X vssd1 vssd1 vccd1
+ vccd1 _08469_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10500_ _12542_/Q _13751_/A vssd1 vssd1 vccd1 vccd1 _10504_/A sky130_fd_sc_hd__xor2_1
XFILLER_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11480_ _13973_/Z _13973_/A _11489_/S vssd1 vssd1 vccd1 vccd1 _11481_/B sky130_fd_sc_hd__mux2_1
X_10431_ _10444_/A _10431_/B vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__and2_1
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10362_ _10362_/A _10362_/B _10362_/C _10362_/D vssd1 vssd1 vccd1 vccd1 _10373_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_109_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12101_ _14078_/A _12101_/B vssd1 vssd1 vccd1 vccd1 _12101_/X sky130_fd_sc_hd__or2_1
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10293_ _13630_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10293_/X sky130_fd_sc_hd__or2_1
X_12032_ _12134_/A vssd1 vssd1 vccd1 vccd1 _12115_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12098__A1 _11064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13983_ _13983_/A _06332_/X vssd1 vssd1 vccd1 vccd1 _13983_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_58_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12934_ _12952_/CLK _12934_/D vssd1 vssd1 vccd1 vccd1 _12934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12865_ _12886_/CLK _12865_/D vssd1 vssd1 vccd1 vccd1 _12865_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11206__A _11206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _11816_/A _11816_/B vssd1 vssd1 vccd1 vccd1 _11817_/A sky130_fd_sc_hd__and2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12799_/CLK _12796_/D vssd1 vssd1 vccd1 vccd1 _13970_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _12864_/Q _14009_/A _11760_/S vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__mux2_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _11688_/A _11688_/B _11688_/C vssd1 vssd1 vccd1 vccd1 _11680_/C sky130_fd_sc_hd__and3_1
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ _13417_/A _07968_/X vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_8
X_10629_ _12571_/Q _13747_/A vssd1 vssd1 vccd1 vccd1 _10632_/B sky130_fd_sc_hd__xor2_1
XFILLER_127_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08250__A _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08624__S1 _08603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _07843_/A _07840_/B _07852_/C vssd1 vssd1 vccd1 vccd1 _07841_/A sky130_fd_sc_hd__or3_1
XFILLER_69_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07771_ _07798_/A vssd1 vssd1 vccd1 vccd1 _07782_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09510_ _13431_/A _09500_/X _09508_/X _09509_/X vssd1 vssd1 vccd1 vccd1 _12300_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06722_ _06722_/A vssd1 vssd1 vccd1 vccd1 _07863_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10939__B _10939_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _11408_/A vssd1 vssd1 vccd1 vccd1 _09455_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06653_ _06680_/A vssd1 vssd1 vccd1 vccd1 _06664_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_80_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09372_ _09370_/X _09372_/B _09372_/C vssd1 vssd1 vccd1 vccd1 _09373_/A sky130_fd_sc_hd__and3b_1
XFILLER_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06584_ _06584_/A _06589_/B _06589_/C vssd1 vssd1 vccd1 vccd1 _06585_/A sky130_fd_sc_hd__or3_1
X_08323_ _08335_/A vssd1 vssd1 vccd1 vccd1 _08333_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_138_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08254_ _08351_/A vssd1 vssd1 vccd1 vccd1 _08264_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07967__C _07977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08480__A3 _08427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07205_ _07205_/A vssd1 vssd1 vccd1 vccd1 _07216_/B sky130_fd_sc_hd__clkbuf_1
X_08185_ _08185_/A vssd1 vssd1 vccd1 vccd1 _08185_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09965__A0 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07136_ _07136_/A vssd1 vssd1 vccd1 vccd1 _07136_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07983__B _08062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ _07067_/A vssd1 vssd1 vccd1 vccd1 _07067_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10690__A _10703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09193__A1 _09112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07969_ _08089_/A _07969_/B vssd1 vssd1 vccd1 vccd1 _07970_/A sky130_fd_sc_hd__or2_1
XFILLER_74_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09708_ _13501_/A _12355_/Q _09711_/S vssd1 vssd1 vccd1 vccd1 _09709_/B sky130_fd_sc_hd__mux2_1
X_10980_ _10986_/A _10980_/B vssd1 vssd1 vccd1 vccd1 _10981_/A sky130_fd_sc_hd__and2_1
XFILLER_55_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _13464_/A _09627_/X _09638_/X _09634_/X vssd1 vssd1 vccd1 vccd1 _12334_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12650_ _12652_/CLK _12650_/D vssd1 vssd1 vccd1 vccd1 _12650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11601_ _11631_/B _11595_/X _11600_/Y vssd1 vssd1 vccd1 vccd1 _12829_/D sky130_fd_sc_hd__a21oi_1
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12581_ _12598_/CLK _12581_/D vssd1 vssd1 vccd1 vccd1 _12581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ _11626_/D _11530_/A _11521_/X vssd1 vssd1 vccd1 vccd1 _11533_/B sky130_fd_sc_hd__o21ai_1
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08335__A _08335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ _14063_/Z _11494_/B vssd1 vssd1 vccd1 vccd1 _11463_/X sky130_fd_sc_hd__or2_1
XFILLER_125_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10414_ _11189_/A vssd1 vssd1 vccd1 vccd1 _10414_/X sky130_fd_sc_hd__buf_4
XFILLER_136_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11394_ _12763_/Q _13938_/A vssd1 vssd1 vccd1 vccd1 _11395_/D sky130_fd_sc_hd__xor2_1
XFILLER_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10345_ _13661_/A _12515_/Q _10348_/S vssd1 vssd1 vccd1 vccd1 _10346_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09708__A0 _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ _13624_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10276_/X sky130_fd_sc_hd__or2_1
XANTENNA__08606__S1 _08576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09184__A1 _09182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ _12134_/A vssd1 vssd1 vccd1 vccd1 _12030_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_repeater104_A peripheralBus_data[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13966_ _13966_/A _06382_/X vssd1 vssd1 vccd1 vccd1 _14126_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_81_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output33_A _13979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12917_ _12917_/CLK _12917_/D vssd1 vssd1 vccd1 vccd1 _14044_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13897_ _13897_/A _06566_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[26] sky130_fd_sc_hd__ebufn_8
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12848_ _12850_/CLK _12848_/D vssd1 vssd1 vccd1 vccd1 _12848_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13192__348 vssd1 vssd1 vccd1 vccd1 _13192__348/HI _13799_/A sky130_fd_sc_hd__conb_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _12782_/CLK _12779_/D vssd1 vssd1 vccd1 vccd1 _13905_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13233__389 vssd1 vssd1 vccd1 vccd1 _13233__389/HI _13888_/A sky130_fd_sc_hd__conb_1
XANTENNA__09947__A0 _14102_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10006__B1 _09994_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09990_ _09997_/C _09993_/C vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__and2_1
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13086__242 vssd1 vssd1 vccd1 vccd1 _13086__242/HI _13581_/A sky130_fd_sc_hd__conb_1
X_08941_ _09067_/A vssd1 vssd1 vccd1 vccd1 _08941_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ _10907_/A _10922_/A _12654_/Q _12655_/Q _08779_/X _08780_/X vssd1 vssd1 vccd1
+ vccd1 _08872_/X sky130_fd_sc_hd__mux4_2
XFILLER_69_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07823_ _07823_/A vssd1 vssd1 vccd1 vccd1 _07823_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13127__283 vssd1 vssd1 vccd1 vccd1 _13127__283/HI _13668_/A sky130_fd_sc_hd__conb_1
XFILLER_38_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07754_ _07754_/A vssd1 vssd1 vccd1 vccd1 _07754_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06705_ _06705_/A vssd1 vssd1 vccd1 vccd1 _06705_/X sky130_fd_sc_hd__clkbuf_1
X_07685_ _07698_/A vssd1 vssd1 vccd1 vccd1 _07696_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_25_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_91_clk _12438_/CLK vssd1 vssd1 vccd1 vccd1 _12414_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09424_ _11408_/A vssd1 vssd1 vccd1 vccd1 _09439_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06636_ input19/X vssd1 vssd1 vccd1 vccd1 _06637_/A sky130_fd_sc_hd__clkinv_2
XFILLER_12_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09355_ _09362_/C _09355_/B vssd1 vssd1 vccd1 vccd1 _09358_/B sky130_fd_sc_hd__and2_1
XFILLER_40_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06567_ _06569_/A _06574_/B _06574_/C vssd1 vssd1 vccd1 vccd1 _06568_/A sky130_fd_sc_hd__or3_1
X_08306_ _08306_/A vssd1 vssd1 vccd1 vccd1 _08306_/X sky130_fd_sc_hd__clkbuf_1
X_09286_ _09322_/B _09276_/X _09322_/A vssd1 vssd1 vccd1 vccd1 _09287_/C sky130_fd_sc_hd__a21o_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06498_ _06498_/A vssd1 vssd1 vccd1 vccd1 _06498_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08237_ _08263_/A vssd1 vssd1 vccd1 vccd1 _08248_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__13996__A _13996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09938__A0 _14035_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08168_ _08168_/A _08285_/B vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__or2_1
XFILLER_119_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07119_ _07119_/A vssd1 vssd1 vccd1 vccd1 _07119_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08099_ _08101_/A _08101_/B _08105_/C vssd1 vssd1 vccd1 vccd1 _08100_/A sky130_fd_sc_hd__or3_1
XFILLER_106_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10130_ _10130_/A _10130_/B _10130_/C _10130_/D vssd1 vssd1 vccd1 vccd1 _10137_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10061_ _10088_/C _10060_/C _10099_/C vssd1 vssd1 vccd1 vccd1 _10062_/C sky130_fd_sc_hd__a21o_1
XFILLER_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13820_ _13820_/A _06779_/X vssd1 vssd1 vccd1 vccd1 _14012_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13751_ _13751_/A _06964_/X vssd1 vssd1 vccd1 vccd1 _14103_/Z sky130_fd_sc_hd__ebufn_8
X_10963_ _10969_/A _10963_/B vssd1 vssd1 vccd1 vccd1 _10964_/A sky130_fd_sc_hd__and2_1
XFILLER_44_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_82_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _12617_/CLK sky130_fd_sc_hd__clkbuf_16
X_12702_ _12704_/CLK _12702_/D vssd1 vssd1 vccd1 vccd1 _12702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13682_ _13682_/A _07141_/X vssd1 vssd1 vccd1 vccd1 _14098_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10894_ _10908_/A _10897_/C _10908_/C _10894_/D vssd1 vssd1 vccd1 vccd1 _10895_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12633_ _12634_/CLK _12633_/D vssd1 vssd1 vccd1 vccd1 _12633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ _12565_/CLK _12564_/D vssd1 vssd1 vccd1 vccd1 _13692_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11515_ _11576_/A vssd1 vssd1 vccd1 vccd1 _11515_/X sky130_fd_sc_hd__clkbuf_4
X_12495_ _12522_/CLK _12495_/D vssd1 vssd1 vccd1 vccd1 _13625_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11446_ _13915_/A _11450_/B vssd1 vssd1 vccd1 vccd1 _11446_/X sky130_fd_sc_hd__or2_1
XFILLER_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11200__A2 _11185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11377_ _11377_/A _11377_/B vssd1 vssd1 vccd1 vccd1 _11378_/A sky130_fd_sc_hd__and2_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _13656_/A _12510_/Q _10342_/S vssd1 vssd1 vccd1 vccd1 _10329_/B sky130_fd_sc_hd__mux2_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _14096_/A _08199_/X vssd1 vssd1 vccd1 vccd1 _14096_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__06313__A _07045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _09750_/X _10249_/X _10258_/X _10256_/X vssd1 vssd1 vccd1 vccd1 _12487_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09004__S1 _08947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13949_ _13949_/A _06424_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[14] sky130_fd_sc_hd__ebufn_8
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _12554_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07470_ _07470_/A vssd1 vssd1 vccd1 vccd1 _07470_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06983__A _08210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06421_ _06428_/A _06425_/B vssd1 vssd1 vccd1 vccd1 _06422_/A sky130_fd_sc_hd__or2_1
XFILLER_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09140_ _09140_/A _09145_/A vssd1 vssd1 vccd1 vccd1 _09140_/X sky130_fd_sc_hd__or2_1
X_06352_ _06547_/A vssd1 vssd1 vccd1 vccd1 _06362_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09071_ _09066_/X _09070_/X _09071_/S vssd1 vssd1 vccd1 vccd1 _10941_/A sky130_fd_sc_hd__mux2_1
X_06283_ _08186_/A vssd1 vssd1 vccd1 vccd1 _06694_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ _08022_/A vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__08703__A _09848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__S1 _08808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09973_ _09982_/A _12421_/Q _12422_/Q vssd1 vssd1 vccd1 vccd1 _09975_/B sky130_fd_sc_hd__a21o_1
XFILLER_115_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08924_ _13970_/A vssd1 vssd1 vccd1 vccd1 _08924_/X sky130_fd_sc_hd__buf_2
XFILLER_85_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11783__B _13363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _10907_/D _10907_/C _10907_/B _10907_/A _08779_/X _08780_/X vssd1 vssd1 vccd1
+ vccd1 _08855_/X sky130_fd_sc_hd__mux4_2
XFILLER_57_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07806_ _07809_/A _07806_/B _07815_/C vssd1 vssd1 vccd1 vccd1 _07807_/A sky130_fd_sc_hd__or3_1
X_08786_ _13777_/A vssd1 vssd1 vccd1 vccd1 _08786_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07737_ _07742_/A _07737_/B _07748_/C vssd1 vssd1 vccd1 vccd1 _07738_/A sky130_fd_sc_hd__or3_1
XFILLER_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_64_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _12820_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__07989__A _07997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ _07668_/A vssd1 vssd1 vccd1 vccd1 _07668_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06893__A _07371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09407_ _11408_/A vssd1 vssd1 vccd1 vccd1 _09422_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12207__A1 _11184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06619_ _06680_/A vssd1 vssd1 vccd1 vccd1 _06630_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07599_ _07599_/A vssd1 vssd1 vccd1 vccd1 _07599_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11415__C1 _11319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09338_ _09363_/A _09338_/B vssd1 vssd1 vccd1 vccd1 _12259_/D sky130_fd_sc_hd__nor2_1
XFILLER_138_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ _09269_/A _09334_/C _09285_/C vssd1 vssd1 vccd1 vccd1 _09276_/C sky130_fd_sc_hd__and3_1
X_11300_ _11325_/B vssd1 vssd1 vccd1 vccd1 _11310_/B sky130_fd_sc_hd__clkbuf_1
X_12280_ _12289_/CLK _12280_/D vssd1 vssd1 vccd1 vccd1 _12280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08809__S1 _08808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ _13879_/A _12735_/Q _11231_/S vssd1 vssd1 vccd1 vccd1 _11232_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11162_ _11160_/X _11155_/X _11161_/X _11068_/X vssd1 vssd1 vccd1 vccd1 _12712_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _10137_/C vssd1 vssd1 vccd1 vccd1 _10126_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11093_ _11093_/A vssd1 vssd1 vccd1 vccd1 _12699_/D sky130_fd_sc_hd__clkbuf_1
X_10044_ _10052_/D _10045_/C _10043_/Y vssd1 vssd1 vccd1 vccd1 _12439_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__10154__C1 _09987_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08993__S0 _08946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13803_ _13803_/A _06829_/X vssd1 vssd1 vccd1 vccd1 _13995_/Z sky130_fd_sc_hd__ebufn_8
X_11995_ _12924_/Q _14067_/A _11995_/S vssd1 vssd1 vccd1 vccd1 _11996_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_55_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _12799_/CLK sky130_fd_sc_hd__clkbuf_16
X_13734_ _13734_/A _07006_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[23] sky130_fd_sc_hd__ebufn_8
X_10946_ _10952_/A _10946_/B vssd1 vssd1 vccd1 vccd1 _10947_/A sky130_fd_sc_hd__and2_1
XFILLER_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13665_ _13665_/A _07186_/X vssd1 vssd1 vccd1 vccd1 _14113_/Z sky130_fd_sc_hd__ebufn_8
X_10877_ _10877_/A _10877_/B _10877_/C _10877_/D vssd1 vssd1 vccd1 vccd1 _10880_/D
+ sky130_fd_sc_hd__and4_1
X_12616_ _12617_/CLK _12616_/D vssd1 vssd1 vccd1 vccd1 _12616_/Q sky130_fd_sc_hd__dfxtp_1
X_13596_ _13596_/A _07375_/X vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__11957__A0 _09638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12547_ _12599_/CLK _12547_/D vssd1 vssd1 vccd1 vccd1 _12547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12478_ _12656_/CLK _12478_/D vssd1 vssd1 vccd1 vccd1 _12478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11429_ _13909_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11429_/X sky130_fd_sc_hd__or2_1
XFILLER_6_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08242__B _08248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14079_ _14079_/A _08038_/X vssd1 vssd1 vccd1 vccd1 _14079_/Z sky130_fd_sc_hd__ebufn_8
X_06970_ _06972_/A _06977_/B vssd1 vssd1 vccd1 vccd1 _06971_/A sky130_fd_sc_hd__or2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08640_ _10099_/C _10098_/C _10098_/B _12447_/Q _08575_/X _08576_/X vssd1 vssd1 vccd1
+ vccd1 _08640_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08571_ _09397_/A vssd1 vssd1 vccd1 vccd1 _13551_/A sky130_fd_sc_hd__buf_4
X_13198__354 vssd1 vssd1 vccd1 vccd1 _13198__354/HI _13805_/A sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_46_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _12597_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07522_ _07531_/A _07531_/B _07524_/C vssd1 vssd1 vccd1 vccd1 _07523_/A sky130_fd_sc_hd__or3_1
XANTENNA__08736__S0 _08733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07453_ _07453_/A vssd1 vssd1 vccd1 vccd1 _07453_/X sky130_fd_sc_hd__clkbuf_1
X_13239__395 vssd1 vssd1 vccd1 vccd1 _13239__395/HI _13894_/A sky130_fd_sc_hd__conb_1
XFILLER_50_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06404_ _06404_/A vssd1 vssd1 vccd1 vccd1 _06404_/X sky130_fd_sc_hd__clkbuf_1
X_07384_ _09125_/A vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11948__A0 _09631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09123_ _13775_/Z vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__clkbuf_4
X_06335_ _06361_/A vssd1 vssd1 vccd1 vccd1 _06346_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09054_ _09050_/X _09053_/X _09071_/S vssd1 vssd1 vccd1 vccd1 _10940_/C sky130_fd_sc_hd__mux2_1
X_06266_ _06377_/C vssd1 vssd1 vccd1 vccd1 _09096_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__11778__B _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07975__C _07977_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08005_ _08010_/A _08005_/B _08016_/C vssd1 vssd1 vccd1 vccd1 _08006_/A sky130_fd_sc_hd__or3_1
XANTENNA__11176__A1 _10659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09956_ _13593_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _09956_/X sky130_fd_sc_hd__or2_1
XANTENNA__07991__B _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08907_ _08904_/X _08906_/X _10710_/A vssd1 vssd1 vccd1 vccd1 _10165_/D sky130_fd_sc_hd__mux2_1
XFILLER_131_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09756_/X _09874_/X _09886_/X _09878_/X vssd1 vssd1 vccd1 vccd1 _12395_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08838_ _08850_/A vssd1 vssd1 vccd1 vccd1 _08838_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11018__B _13935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _13779_/A vssd1 vssd1 vccd1 vccd1 _08769_/X sky130_fd_sc_hd__buf_2
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _12722_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _10863_/A _10800_/B vssd1 vssd1 vccd1 vccd1 _10801_/B sky130_fd_sc_hd__and2_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11780_/A _11780_/B _11780_/C _11780_/D vssd1 vssd1 vccd1 vccd1 _11786_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07512__A _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ _10285_/X _10703_/S _10730_/X _10711_/X vssd1 vssd1 vccd1 vccd1 _12612_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13450_ _13450_/A _07752_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__07231__B _07231_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10662_ _10662_/A vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__buf_6
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ _12404_/CLK _12401_/D vssd1 vssd1 vccd1 vccd1 _13529_/A sky130_fd_sc_hd__dfxtp_1
X_13381_ _13381_/A _08330_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
X_10593_ _10602_/A _10593_/B vssd1 vssd1 vccd1 vccd1 _10594_/A sky130_fd_sc_hd__and2_1
X_12332_ _12334_/CLK _12332_/D vssd1 vssd1 vccd1 vccd1 _13462_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ _12264_/CLK _12263_/D vssd1 vssd1 vccd1 vccd1 _12263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11167__A1 _10648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08062__B _08062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032__188 vssd1 vssd1 vccd1 vccd1 _13032__188/HI _13475_/A sky130_fd_sc_hd__conb_1
X_14002_ _14002_/A _07955_/X vssd1 vssd1 vccd1 vccd1 _14066_/Z sky130_fd_sc_hd__ebufn_8
X_11214_ _11221_/A _11214_/B vssd1 vssd1 vccd1 vccd1 _11215_/A sky130_fd_sc_hd__and2_1
X_12194_ _11170_/X _12182_/X _12193_/X _12187_/X vssd1 vssd1 vccd1 vccd1 _12975_/D
+ sky130_fd_sc_hd__o211a_1
Xoutput40 _13595_/A vssd1 vssd1 vccd1 vccd1 pwm_en[6] sky130_fd_sc_hd__buf_2
Xoutput51 _13376_/A vssd1 vssd1 vccd1 vccd1 pwm_out[1] sky130_fd_sc_hd__buf_2
XFILLER_122_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11145_ _12694_/Q _13935_/A vssd1 vssd1 vccd1 vccd1 _11148_/B sky130_fd_sc_hd__xor2_1
XFILLER_96_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11076_ _11076_/A vssd1 vssd1 vccd1 vccd1 _12694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_94_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10027_ _10027_/A vssd1 vssd1 vccd1 vccd1 _12435_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08966__S0 _08941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09902__A _09902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk _12759_/CLK vssd1 vssd1 vccd1 vccd1 _12758_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11978_ _11978_/A _11978_/B vssd1 vssd1 vccd1 vccd1 _11979_/A sky130_fd_sc_hd__and2_1
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10929_ _10932_/B vssd1 vssd1 vccd1 vccd1 _10929_/Y sky130_fd_sc_hd__inv_2
X_13717_ _13717_/A _07048_/X vssd1 vssd1 vccd1 vccd1 _13973_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_32_clk_A _12759_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ _13648_/A _07232_/X vssd1 vssd1 vccd1 vccd1 _14096_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13579_ _13579_/A _07422_/X vssd1 vssd1 vccd1 vccd1 _14027_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08253__A _08266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_47_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09810_ _13524_/A _12379_/Q _09820_/S vssd1 vssd1 vccd1 vccd1 _09811_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09741_ _09776_/A vssd1 vssd1 vccd1 vccd1 _09741_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06953_ _06960_/A _06953_/B vssd1 vssd1 vccd1 vccd1 _06954_/A sky130_fd_sc_hd__or2_1
XFILLER_101_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_105_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09672_ _09711_/S vssd1 vssd1 vccd1 vccd1 _09685_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06884_ _06890_/A _06884_/B _06884_/C vssd1 vssd1 vccd1 vccd1 _06885_/A sky130_fd_sc_hd__or3_1
XFILLER_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08623_ _12426_/Q vssd1 vssd1 vccd1 vccd1 _09997_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_repeater66_A _14102_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_clk _12881_/CLK vssd1 vssd1 vccd1 vccd1 _12923_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _13585_/A vssd1 vssd1 vccd1 vccd1 _08554_/X sky130_fd_sc_hd__buf_2
XFILLER_70_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07505_ _07505_/A vssd1 vssd1 vccd1 vccd1 _07505_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08485_ _11705_/C vssd1 vssd1 vccd1 vccd1 _13365_/A sky130_fd_sc_hd__buf_4
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ _07436_/A vssd1 vssd1 vccd1 vccd1 _07436_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07367_ _07369_/A _07377_/B _07374_/C vssd1 vssd1 vccd1 vccd1 _07368_/A sky130_fd_sc_hd__or3_1
XANTENNA__07986__B _08062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10693__A _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ _11503_/B vssd1 vssd1 vccd1 vccd1 _09967_/B sky130_fd_sc_hd__buf_4
X_06318_ _06320_/A _06323_/B _06323_/C vssd1 vssd1 vccd1 vccd1 _06319_/A sky130_fd_sc_hd__or3_1
XFILLER_136_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07298_ _07307_/A _07303_/B _07300_/C vssd1 vssd1 vccd1 vccd1 _07299_/A sky130_fd_sc_hd__or3_1
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09037_ _09002_/X _09004_/X _09008_/X _09036_/X _08994_/X _08996_/X vssd1 vssd1 vccd1
+ vccd1 _09037_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09762__A1 _09160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07507__A _07507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09940_/A sky130_fd_sc_hd__or2_1
XANTENNA__11029__A _11070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13_0_clk/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__07226__B _07231_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ _12952_/CLK _12950_/D vssd1 vssd1 vccd1 vccd1 _14076_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08948__S0 _08946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11901_ _12896_/Q _13368_/A vssd1 vssd1 vccd1 vccd1 _11905_/A sky130_fd_sc_hd__xor2_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _12881_/CLK _12881_/D vssd1 vssd1 vccd1 vccd1 _14009_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _11832_/A vssd1 vssd1 vccd1 vccd1 _12882_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__A _08338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _12869_/Q _14014_/A _11763_/S vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__mux2_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08057__B _08110_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ hold2/X _07617_/X vssd1 vssd1 vccd1 vccd1 _14110_/Z sky130_fd_sc_hd__ebufn_8
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10720_/A _10714_/B vssd1 vssd1 vccd1 vccd1 _10715_/A sky130_fd_sc_hd__or2_1
XFILLER_41_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11694_/A _11694_/B vssd1 vssd1 vccd1 vccd1 _12850_/D sky130_fd_sc_hd__nor2_1
X_13433_ _13433_/A _07797_/X vssd1 vssd1 vccd1 vccd1 _13625_/Z sky130_fd_sc_hd__ebufn_8
X_10645_ _10645_/A vssd1 vssd1 vccd1 vccd1 _10645_/X sky130_fd_sc_hd__buf_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09169__A _09633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13364_ _13364_/A _08289_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[5] sky130_fd_sc_hd__ebufn_8
XFILLER_154_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10576_ _10585_/A _10576_/B vssd1 vssd1 vccd1 vccd1 _10577_/A sky130_fd_sc_hd__and2_1
X_12315_ _12320_/CLK _12315_/D vssd1 vssd1 vccd1 vccd1 _12315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater134_A peripheralBus_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12246_ _12251_/CLK _12246_/D vssd1 vssd1 vccd1 vccd1 _12246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10899__B1 _10757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ _12177_/A _12177_/B _12177_/C vssd1 vssd1 vccd1 vccd1 _12178_/B sky130_fd_sc_hd__or3_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11128_ _12707_/Q _13948_/A vssd1 vssd1 vccd1 vccd1 _11128_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07417__A _07417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12042__B _13365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ _13818_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11059_/X sky130_fd_sc_hd__or2_1
XFILLER_49_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10497__B _13745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ _08276_/A _08274_/B _08276_/C vssd1 vssd1 vccd1 vccd1 _08271_/A sky130_fd_sc_hd__or3_1
XFILLER_149_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07221_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07221_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater70 peripheralBus_data[6] vssd1 vssd1 vccd1 vccd1 _14069_/Z sky130_fd_sc_hd__buf_12
Xrepeater81 _14126_/Z vssd1 vssd1 vccd1 vccd1 _14030_/Z sky130_fd_sc_hd__buf_12
Xrepeater92 _13994_/Z vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__buf_12
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09079__A _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07152_ _07152_/A _07163_/B _07160_/C vssd1 vssd1 vccd1 vccd1 _07153_/A sky130_fd_sc_hd__or3_1
XFILLER_157_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07083_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07094_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_clk _12917_/CLK vssd1 vssd1 vccd1 vccd1 _12904_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07327__A _07473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07985_ _07999_/A vssd1 vssd1 vccd1 vccd1 _07997_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09724_ _12355_/Q _13565_/A vssd1 vssd1 vccd1 vccd1 _09725_/D sky130_fd_sc_hd__xor2_1
X_06936_ _06936_/A _06941_/B vssd1 vssd1 vccd1 vccd1 _06937_/A sky130_fd_sc_hd__or2_1
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09655_ _14110_/Z _09655_/B vssd1 vssd1 vccd1 vccd1 _09655_/X sky130_fd_sc_hd__or2_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06867_ _06867_/A vssd1 vssd1 vccd1 vccd1 _06867_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10688__A _11457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _09997_/B _09997_/A _12429_/Q _12430_/Q _08575_/X _08576_/X vssd1 vssd1 vccd1
+ vccd1 _08606_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_09586_ _12317_/Q _13560_/A vssd1 vssd1 vccd1 vccd1 _09586_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06798_ _06798_/A vssd1 vssd1 vccd1 vccd1 _06798_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08158__A _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07062__A _07406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08537_ _09377_/A _09382_/A _12272_/Q _12273_/Q _09140_/A _09146_/A vssd1 vssd1 vccd1
+ vccd1 _08537_/X sky130_fd_sc_hd__mux4_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13254__410 vssd1 vssd1 vccd1 vccd1 _13254__410/HI _13925_/A sky130_fd_sc_hd__conb_1
XANTENNA__07997__A _07997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ _08375_/X _08381_/X _08378_/X _08386_/X _08517_/A _08467_/X vssd1 vssd1 vccd1
+ vccd1 _08468_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ _07480_/A vssd1 vssd1 vccd1 vccd1 _07468_/A sky130_fd_sc_hd__buf_2
XANTENNA__10290__A1 _10288_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08399_ _12238_/Q vssd1 vssd1 vccd1 vccd1 _09258_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11312__A _11312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ _13679_/A _12534_/Q _10507_/B vssd1 vssd1 vccd1 vccd1 _10431_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10361_ _12515_/Q _13757_/A vssd1 vssd1 vccd1 vccd1 _10362_/D sky130_fd_sc_hd__xor2_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12100_ _10548_/A _12088_/X _12099_/X _12097_/X vssd1 vssd1 vccd1 vccd1 _12951_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10292_ _09116_/X _10278_/X _10291_/X _10283_/X vssd1 vssd1 vccd1 vccd1 _12499_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _12031_/A vssd1 vssd1 vccd1 vccd1 _12934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11982__A _12033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13982_ _13982_/A _06334_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[15] sky130_fd_sc_hd__ebufn_8
XFILLER_74_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12933_ _12952_/CLK _12933_/D vssd1 vssd1 vccd1 vccd1 _12933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12864_ _12886_/CLK _12864_/D vssd1 vssd1 vccd1 vccd1 _12864_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11815_ _09633_/A _14006_/A _11823_/S vssd1 vssd1 vccd1 vccd1 _11816_/B sky130_fd_sc_hd__mux2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12799_/CLK _12795_/D vssd1 vssd1 vccd1 vccd1 _13969_/A sky130_fd_sc_hd__dfxtp_2
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _11763_/S vssd1 vssd1 vccd1 vccd1 _11760_/S sky130_fd_sc_hd__buf_2
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10281__A1 _09182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11677_ _11677_/A _11677_/B _11677_/C vssd1 vssd1 vccd1 vccd1 _11688_/C sky130_fd_sc_hd__and3_1
X_13038__194 vssd1 vssd1 vccd1 vccd1 _13038__194/HI _13481_/A sky130_fd_sc_hd__conb_1
X_10628_ _12575_/Q _13751_/A vssd1 vssd1 vccd1 vccd1 _10632_/A sky130_fd_sc_hd__xor2_1
X_13416_ _13416_/A _08088_/X vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__12037__B _13370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11579__D _11649_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10559_ _10559_/A vssd1 vssd1 vccd1 vccd1 _12567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09627__A _09640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12229_ _12301_/CLK _12229_/D vssd1 vssd1 vccd1 vccd1 _12229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07147__A _08364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07770_ _07770_/A vssd1 vssd1 vccd1 vccd1 _07770_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06986__A _07979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06721_ _06753_/A vssd1 vssd1 vccd1 vccd1 _06738_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09440_ _09440_/A vssd1 vssd1 vccd1 vccd1 _12285_/D sky130_fd_sc_hd__clkbuf_1
X_06652_ _06652_/A vssd1 vssd1 vccd1 vccd1 _06652_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09371_ _09347_/A _09382_/B _09377_/C vssd1 vssd1 vccd1 vccd1 _09372_/C sky130_fd_sc_hd__a21o_1
XFILLER_52_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06583_ _06583_/A vssd1 vssd1 vccd1 vccd1 _06583_/X sky130_fd_sc_hd__clkbuf_1
X_08322_ _08322_/A vssd1 vssd1 vccd1 vccd1 _08322_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08253_ _08266_/A vssd1 vssd1 vccd1 vccd1 _08264_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_165_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07204_ _07204_/A vssd1 vssd1 vccd1 vccd1 _07204_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08184_ _08184_/A _08184_/B _08184_/C vssd1 vssd1 vccd1 vccd1 _08185_/A sky130_fd_sc_hd__or3_1
X_07135_ _07135_/A _07145_/B _07142_/C vssd1 vssd1 vccd1 vccd1 _07136_/A sky130_fd_sc_hd__or3_1
XANTENNA__10971__A _10971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07066_ _08180_/A _07076_/B _07073_/C vssd1 vssd1 vccd1 vccd1 _07067_/A sky130_fd_sc_hd__or3_1
XFILLER_160_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07968_ _07968_/A vssd1 vssd1 vccd1 vccd1 _07968_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06896__A _07328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ _09836_/A vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06919_ _06923_/A _06929_/B vssd1 vssd1 vccd1 vccd1 _06920_/A sky130_fd_sc_hd__or2_1
X_07899_ _07908_/A _07903_/B _07903_/C vssd1 vssd1 vccd1 vccd1 _07900_/A sky130_fd_sc_hd__or3_1
X_09638_ _09638_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09638_/X sky130_fd_sc_hd__or2_1
XFILLER_82_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11026__B _11026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ _13466_/A _12319_/Q _09575_/S vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__mux2_1
X_11600_ _11631_/B _11595_/X _11505_/B vssd1 vssd1 vccd1 vccd1 _11600_/Y sky130_fd_sc_hd__o21ai_1
X_12580_ _12802_/CLK _12580_/D vssd1 vssd1 vccd1 vccd1 _12580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07520__A _08210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10263__A1 _09756_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ _11626_/D _11625_/C _11531_/C vssd1 vssd1 vccd1 vccd1 _11533_/A sky130_fd_sc_hd__and3_1
XFILLER_156_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11042__A _11070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11462_ _11499_/B vssd1 vssd1 vccd1 vccd1 _11494_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_137_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10413_ _10408_/X _10409_/X _10411_/X _10412_/X vssd1 vssd1 vccd1 vccd1 _12528_/D
+ sky130_fd_sc_hd__o211a_1
X_11393_ _12766_/Q _13941_/A vssd1 vssd1 vccd1 vccd1 _11395_/C sky130_fd_sc_hd__xor2_1
XFILLER_109_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10344_ _10344_/A vssd1 vssd1 vccd1 vccd1 _12514_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08351__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10275_ _09770_/X _10264_/X _10274_/X _10270_/X vssd1 vssd1 vccd1 vccd1 _12493_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12014_ _12014_/A vssd1 vssd1 vccd1 vccd1 _12929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09182__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13965_ _13965_/A _06384_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[30] sky130_fd_sc_hd__ebufn_8
X_12916_ _12918_/CLK _12916_/D vssd1 vssd1 vccd1 vccd1 _14043_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13896_ _13896_/A _06568_/X vssd1 vssd1 vccd1 vccd1 _14120_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_34_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _12850_/CLK _12847_/D vssd1 vssd1 vccd1 vccd1 _12847_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12780_/CLK _12778_/D vssd1 vssd1 vccd1 vccd1 _13904_/A sky130_fd_sc_hd__dfxtp_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10254__A1 _09124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11729_ _11763_/S vssd1 vssd1 vccd1 vccd1 _11743_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_147_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08940_ _12811_/Q vssd1 vssd1 vccd1 vccd1 _11625_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08871_ _12653_/Q vssd1 vssd1 vccd1 vccd1 _10922_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07822_ _07822_/A _07822_/B _07822_/C vssd1 vssd1 vccd1 vccd1 _07823_/A sky130_fd_sc_hd__or3_1
XANTENNA__09092__A _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _07756_/A _07753_/B _07761_/C vssd1 vssd1 vccd1 vccd1 _07754_/A sky130_fd_sc_hd__or3_1
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06704_ _06714_/A _06706_/B _06706_/C vssd1 vssd1 vccd1 vccd1 _06705_/A sky130_fd_sc_hd__or3_1
XANTENNA__10031__A _10101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07684_ _07684_/A vssd1 vssd1 vccd1 vccd1 _07684_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09423_ _09423_/A vssd1 vssd1 vccd1 vccd1 _12280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06635_ _06635_/A vssd1 vssd1 vccd1 vccd1 _06635_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09354_ _09362_/C _09355_/B _09248_/X vssd1 vssd1 vccd1 vccd1 _09356_/A sky130_fd_sc_hd__o21ai_1
XFILLER_80_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06566_ _06566_/A vssd1 vssd1 vccd1 vccd1 _06566_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08305_ _08312_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08306_/A sky130_fd_sc_hd__or2_1
XANTENNA__10245__A1 _13762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _13391_/A _09334_/C _09285_/C _09331_/A vssd1 vssd1 vccd1 vccd1 _09292_/C
+ sky130_fd_sc_hd__and4_1
X_06497_ _06507_/A _06499_/B _06499_/C vssd1 vssd1 vccd1 vccd1 _06498_/A sky130_fd_sc_hd__or3_1
X_08236_ _08236_/A vssd1 vssd1 vccd1 vccd1 _08236_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08167_ _08364_/C vssd1 vssd1 vccd1 vccd1 _08285_/B sky130_fd_sc_hd__clkbuf_1
X_07118_ _07121_/A _07118_/B _07128_/C vssd1 vssd1 vccd1 vccd1 _07119_/A sky130_fd_sc_hd__or3_1
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08171__A _08228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08098_ _08098_/A vssd1 vssd1 vccd1 vccd1 _08098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07049_ _07055_/A _07055_/B vssd1 vssd1 vccd1 vccd1 _07050_/A sky130_fd_sc_hd__or2_1
XFILLER_161_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06403__B _06412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ _10099_/C _10088_/C _10060_/C vssd1 vssd1 vccd1 vccd1 _10064_/B sky130_fd_sc_hd__and3_1
XFILLER_125_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09714__B _13560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10962_ _13812_/A _12666_/Q _10972_/S vssd1 vssd1 vccd1 vccd1 _10963_/B sky130_fd_sc_hd__mux2_1
XFILLER_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13750_ _13750_/A _06966_/X vssd1 vssd1 vccd1 vccd1 _13974_/Z sky130_fd_sc_hd__ebufn_8
XANTENNA__07234__B _07947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ _12704_/CLK _12701_/D vssd1 vssd1 vccd1 vccd1 _12701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10893_ _10897_/C _10891_/B _10908_/A vssd1 vssd1 vccd1 vccd1 _10895_/B sky130_fd_sc_hd__a21oi_1
X_13681_ _13681_/A _07143_/X vssd1 vssd1 vccd1 vccd1 _14097_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12632_ _12634_/CLK _12632_/D vssd1 vssd1 vccd1 vccd1 _12632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12563_ _12565_/CLK _12563_/D vssd1 vssd1 vccd1 vccd1 _13691_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11514_ _11518_/B _11514_/B vssd1 vssd1 vccd1 vccd1 _11517_/A sky130_fd_sc_hd__and2_1
XFILLER_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12494_ _12522_/CLK _12494_/D vssd1 vssd1 vccd1 vccd1 _13624_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ _11189_/X _11438_/X _11442_/X _11444_/X vssd1 vssd1 vccd1 vccd1 _12788_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09177__A _14072_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ _13917_/A _12774_/Q _11381_/S vssd1 vssd1 vccd1 vccd1 _11377_/B sky130_fd_sc_hd__mux2_1
X_10327_ _10348_/S vssd1 vssd1 vccd1 vccd1 _10342_/S sky130_fd_sc_hd__clkbuf_2
X_14095_ _14095_/A _08181_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[0] sky130_fd_sc_hd__ebufn_8
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10258_ _13617_/A _10262_/B vssd1 vssd1 vccd1 vccd1 _10258_/X sky130_fd_sc_hd__or2_1
XFILLER_79_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ _10189_/A vssd1 vssd1 vccd1 vccd1 _12473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07425__A _08131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13948_ _13948_/A _06426_/X vssd1 vssd1 vccd1 vccd1 _14012_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09640__A _09640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13200__356 vssd1 vssd1 vccd1 vccd1 _13200__356/HI _13823_/A sky130_fd_sc_hd__conb_1
XFILLER_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13879_ _13879_/A _06615_/X vssd1 vssd1 vccd1 vccd1 _14007_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11381__S _11381_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06983__B _06983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06420_ _06420_/A vssd1 vssd1 vccd1 vccd1 _06420_/X sky130_fd_sc_hd__clkbuf_1
X_06351_ _06462_/A vssd1 vssd1 vccd1 vccd1 _06362_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_147_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09070_ _08933_/X _09015_/X _09041_/X _09069_/X _08994_/X _08996_/X vssd1 vssd1 vccd1
+ vccd1 _09070_/X sky130_fd_sc_hd__mux4_1
X_06282_ _07603_/A vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__buf_2
XFILLER_147_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ _08021_/A vssd1 vssd1 vccd1 vccd1 _08021_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09972_ _10107_/A _12422_/Q _12421_/Q vssd1 vssd1 vccd1 vccd1 _09972_/X sky130_fd_sc_hd__and3_1
XFILLER_89_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08923_ _12819_/Q _12820_/Q _12821_/Q _12822_/Q _08921_/X _08922_/X vssd1 vssd1 vccd1
+ vccd1 _08923_/X sky130_fd_sc_hd__mux4_2
XANTENNA_repeater96_A _14120_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ _12652_/Q vssd1 vssd1 vccd1 vccd1 _10907_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07335__A _07473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07805_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07805_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08785_ _13776_/A vssd1 vssd1 vccd1 vccd1 _08785_/X sky130_fd_sc_hd__clkbuf_4
X_07736_ _07736_/A vssd1 vssd1 vccd1 vccd1 _07736_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11663__B1 _11576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _07672_/A _07669_/B _07678_/C vssd1 vssd1 vccd1 vccd1 _07668_/A sky130_fd_sc_hd__or3_1
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09406_ _09846_/A vssd1 vssd1 vccd1 vccd1 _11408_/A sky130_fd_sc_hd__buf_6
XFILLER_41_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06618_ _06694_/A vssd1 vssd1 vccd1 vccd1 _06680_/A sky130_fd_sc_hd__buf_2
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07598_ _07601_/A _07598_/B _07608_/C vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__or3_1
XFILLER_71_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09337_ _09343_/C _09343_/D _09236_/X vssd1 vssd1 vccd1 vccd1 _09338_/B sky130_fd_sc_hd__o21ai_1
X_06549_ _06577_/A vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__buf_8
XFILLER_21_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09268_ _09328_/B _09328_/C vssd1 vssd1 vccd1 vccd1 _09285_/C sky130_fd_sc_hd__and2_1
XFILLER_154_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08219_ _08219_/A vssd1 vssd1 vccd1 vccd1 _08219_/X sky130_fd_sc_hd__clkbuf_1
X_09199_ _12228_/Q _09380_/A vssd1 vssd1 vccd1 vccd1 _09200_/A sky130_fd_sc_hd__and2b_1
XFILLER_147_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ _11230_/A vssd1 vssd1 vccd1 vccd1 _12734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06414__A _08338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ _13840_/A _11168_/B vssd1 vssd1 vccd1 vccd1 _11161_/X sky130_fd_sc_hd__or2_1
XANTENNA__08690__S0 _08602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ _10112_/A _10112_/B _10133_/C vssd1 vssd1 vccd1 vccd1 _10137_/C sky130_fd_sc_hd__and3_1
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11092_ _11095_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11093_/A sky130_fd_sc_hd__and2_1
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10043_ _10052_/D _10045_/C _09978_/X vssd1 vssd1 vccd1 vccd1 _10043_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input25_A peripheralBus_oe vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08993__S1 _08947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _13802_/A _06831_/X vssd1 vssd1 vccd1 vccd1 _13994_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_90_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11994_ _11994_/A vssd1 vssd1 vccd1 vccd1 _12923_/D sky130_fd_sc_hd__clkbuf_1
X_13733_ _13733_/A _07008_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[22] sky130_fd_sc_hd__ebufn_8
X_10945_ _13807_/A _12661_/Q _10955_/S vssd1 vssd1 vccd1 vccd1 _10946_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13664_ _13664_/A _07188_/X vssd1 vssd1 vccd1 vccd1 _14048_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10876_ _10876_/A _10876_/B _10876_/C _10876_/D vssd1 vssd1 vccd1 vccd1 _10877_/D
+ sky130_fd_sc_hd__and4_1
X_12615_ _12660_/CLK _12615_/D vssd1 vssd1 vccd1 vccd1 _12615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13595_ _13595_/A _07378_/X vssd1 vssd1 vccd1 vccd1 _14107_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_129_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12546_ _12550_/CLK _12546_/D vssd1 vssd1 vccd1 vccd1 _12546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12477_ _12492_/CLK _12477_/D vssd1 vssd1 vccd1 vccd1 _12477_/Q sky130_fd_sc_hd__dfxtp_1
X_11428_ _11170_/X _11425_/X _11427_/X _11417_/X vssd1 vssd1 vccd1 vccd1 _12782_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ _11381_/S vssd1 vssd1 vccd1 vccd1 _11373_/S sky130_fd_sc_hd__buf_2
XFILLER_113_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14078_ _14078_/A _08034_/X vssd1 vssd1 vccd1 vccd1 _14078_/Z sky130_fd_sc_hd__ebufn_8
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11376__S _11381_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_6_clk_A _12917_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10696__A1 _10377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08570_ _08564_/X _08569_/X _13588_/A vssd1 vssd1 vccd1 vccd1 _09397_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07521_ _08197_/A vssd1 vssd1 vccd1 vccd1 _07531_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__08736__S1 _08735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07452_ _07454_/A _07459_/B vssd1 vssd1 vccd1 vccd1 _07453_/A sky130_fd_sc_hd__or2_1
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06403_ _06403_/A _06412_/B vssd1 vssd1 vccd1 vccd1 _06404_/A sky130_fd_sc_hd__or2_1
X_07383_ _07383_/A vssd1 vssd1 vccd1 vccd1 _07383_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09122_ _09120_/X _09100_/X _09121_/X _09109_/X vssd1 vssd1 vccd1 vccd1 _12213_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06334_ _06334_/A vssd1 vssd1 vccd1 vccd1 _06334_/X sky130_fd_sc_hd__clkbuf_1
X_09053_ _08978_/X _08980_/X _09026_/X _09052_/X _08952_/X _08953_/X vssd1 vssd1 vccd1
+ vccd1 _09053_/X sky130_fd_sc_hd__mux4_1
X_06265_ input12/X input1/X vssd1 vssd1 vccd1 vccd1 _06377_/C sky130_fd_sc_hd__or2_4
XFILLER_163_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08004_ _08004_/A vssd1 vssd1 vccd1 vccd1 _08016_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09955_ _09955_/A vssd1 vssd1 vccd1 vccd1 _12416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07991__C _07993_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ _08825_/X _08855_/X _08879_/X _08905_/X _08831_/X _08876_/X vssd1 vssd1 vccd1
+ vccd1 _08906_/X sky130_fd_sc_hd__mux4_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _13523_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09886_/X sky130_fd_sc_hd__or2_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10687__A1 _10552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08837_ _13779_/A vssd1 vssd1 vccd1 vccd1 _08837_/X sky130_fd_sc_hd__buf_2
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _12627_/Q _12628_/Q _12629_/Q _12630_/Q _08766_/X _08767_/X vssd1 vssd1 vccd1
+ vccd1 _08768_/X sky130_fd_sc_hd__mux4_2
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ _07727_/A _07724_/B _07719_/C vssd1 vssd1 vccd1 vccd1 _07720_/A sky130_fd_sc_hd__or3_1
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _10137_/B _10148_/C _12462_/Q _12463_/Q _08602_/X _08603_/X vssd1 vssd1 vccd1
+ vccd1 _08699_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10730_ _13787_/A _10732_/B vssd1 vssd1 vccd1 vccd1 _10730_/X sky130_fd_sc_hd__or2_1
XFILLER_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10661_ _10659_/X _10655_/X _10660_/X _10650_/X vssd1 vssd1 vccd1 vccd1 _12590_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12400_ _12400_/CLK _12400_/D vssd1 vssd1 vccd1 vccd1 _13528_/A sky130_fd_sc_hd__dfxtp_1
X_13380_ _13380_/A _08328_/X vssd1 vssd1 vccd1 vccd1 peripheralBus_data[21] sky130_fd_sc_hd__ebufn_8
X_10592_ _13721_/A _12577_/Q _10601_/S vssd1 vssd1 vccd1 vccd1 _10593_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12331_ _12331_/CLK _12331_/D vssd1 vssd1 vccd1 vccd1 _13461_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12262_ _12264_/CLK _12262_/D vssd1 vssd1 vccd1 vccd1 _12262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11213_ _13874_/A _12730_/Q _11281_/B vssd1 vssd1 vccd1 vccd1 _11214_/B sky130_fd_sc_hd__mux2_1
XFILLER_5_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14001_ _14001_/A _07987_/X vssd1 vssd1 vccd1 vccd1 _14065_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ _14100_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12193_/X sky130_fd_sc_hd__or2_1
Xoutput30 _13788_/A vssd1 vssd1 vccd1 vccd1 pwm_en[11] sky130_fd_sc_hd__buf_2
Xoutput41 _13596_/A vssd1 vssd1 vccd1 vccd1 pwm_en[7] sky130_fd_sc_hd__buf_2
Xoutput52 _13377_/A vssd1 vssd1 vccd1 vccd1 pwm_out[2] sky130_fd_sc_hd__buf_2
X_11144_ _12699_/Q _13940_/A vssd1 vssd1 vccd1 vccd1 _11148_/A sky130_fd_sc_hd__xor2_1
XFILLER_150_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11075_ _11078_/A _11075_/B vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__and2_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11324__C1 _11319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10026_ _10024_/X _10062_/B _10026_/C vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__and3b_1
XFILLER_76_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10678__A1 _10414_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08966__S1 _08942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11977_ _14110_/Z _14046_/A _11977_/S vssd1 vssd1 vccd1 vccd1 _11978_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13716_ _13716_/A _07050_/X vssd1 vssd1 vccd1 vccd1 _14100_/Z sky130_fd_sc_hd__ebufn_8
X_10928_ _12658_/Q _10928_/B _10928_/C vssd1 vssd1 vccd1 vccd1 _10932_/B sky130_fd_sc_hd__and3_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13271__427 vssd1 vssd1 vccd1 vccd1 _13271__427/HI _13962_/A sky130_fd_sc_hd__conb_1
XFILLER_20_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13647_ _13647_/A _07992_/X vssd1 vssd1 vccd1 vccd1 _13775_/Z sky130_fd_sc_hd__ebufn_8
X_10859_ _10875_/A _10859_/B vssd1 vssd1 vccd1 vccd1 _10860_/C sky130_fd_sc_hd__nand2_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13578_/A _07424_/X vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_8
XFILLER_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09349__B _09372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312__468 vssd1 vssd1 vccd1 vccd1 _13312__468/HI _14049_/A sky130_fd_sc_hd__conb_1
X_12529_ _12583_/CLK _12529_/D vssd1 vssd1 vccd1 vccd1 _13658_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08654__S0 _08556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13165__321 vssd1 vssd1 vccd1 vccd1 _13165__321/HI _13738_/A sky130_fd_sc_hd__conb_1
XANTENNA__09365__A _09380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09740_ _11283_/B _09873_/B _10637_/B vssd1 vssd1 vccd1 vccd1 _09776_/A sky130_fd_sc_hd__or3_4
X_06952_ _06952_/A vssd1 vssd1 vccd1 vccd1 _06952_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
.ends

