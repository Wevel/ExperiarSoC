// This is the unpowered netlist.
module CaravelHost (caravel_uart_rx,
    caravel_uart_tx,
    caravel_wb_ack_i,
    caravel_wb_cyc_o,
    caravel_wb_error_i,
    caravel_wb_stall_i,
    caravel_wb_stb_o,
    caravel_wb_we_o,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    caravel_irq,
    caravel_wb_adr_o,
    caravel_wb_data_i,
    caravel_wb_data_o,
    caravel_wb_sel_o,
    core0Index,
    core1Index,
    la_data_out,
    manufacturerID,
    partID,
    probe_out,
    versionID,
    wbs_adr_i,
    wbs_data_i,
    wbs_data_o,
    wbs_sel_i);
 input caravel_uart_rx;
 output caravel_uart_tx;
 input caravel_wb_ack_i;
 output caravel_wb_cyc_o;
 input caravel_wb_error_i;
 input caravel_wb_stall_i;
 output caravel_wb_stb_o;
 output caravel_wb_we_o;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 output [3:0] caravel_irq;
 output [27:0] caravel_wb_adr_o;
 input [31:0] caravel_wb_data_i;
 output [31:0] caravel_wb_data_o;
 output [3:0] caravel_wb_sel_o;
 output [7:0] core0Index;
 output [7:0] core1Index;
 output [127:0] la_data_out;
 output [10:0] manufacturerID;
 output [15:0] partID;
 input [97:0] probe_out;
 output [3:0] versionID;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_data_i;
 output [31:0] wbs_data_o;
 input [3:0] wbs_sel_i;

 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net722;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net670;
 wire net671;
 wire net700;
 wire net710;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net723;
 wire net728;
 wire net729;
 wire net716;
 wire net717;
 wire net730;
 wire net731;
 wire net711;
 wire net724;
 wire net712;
 wire net725;
 wire net713;
 wire net726;
 wire net714;
 wire net727;
 wire net715;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire \device.configuration[0] ;
 wire \device.configuration[10] ;
 wire \device.configuration[11] ;
 wire \device.configuration[12] ;
 wire \device.configuration[13] ;
 wire \device.configuration[14] ;
 wire \device.configuration[15] ;
 wire \device.configuration[16] ;
 wire \device.configuration[17] ;
 wire \device.configuration[18] ;
 wire \device.configuration[19] ;
 wire \device.configuration[1] ;
 wire \device.configuration[20] ;
 wire \device.configuration[2] ;
 wire \device.configuration[3] ;
 wire \device.configuration[4] ;
 wire \device.configuration[5] ;
 wire \device.configuration[6] ;
 wire \device.configuration[7] ;
 wire \device.configuration[8] ;
 wire \device.configuration[9] ;
 wire \device.rxBuffer.buffer[0][0] ;
 wire \device.rxBuffer.buffer[0][1] ;
 wire \device.rxBuffer.buffer[0][2] ;
 wire \device.rxBuffer.buffer[0][3] ;
 wire \device.rxBuffer.buffer[0][4] ;
 wire \device.rxBuffer.buffer[0][5] ;
 wire \device.rxBuffer.buffer[0][6] ;
 wire \device.rxBuffer.buffer[0][7] ;
 wire \device.rxBuffer.buffer[10][0] ;
 wire \device.rxBuffer.buffer[10][1] ;
 wire \device.rxBuffer.buffer[10][2] ;
 wire \device.rxBuffer.buffer[10][3] ;
 wire \device.rxBuffer.buffer[10][4] ;
 wire \device.rxBuffer.buffer[10][5] ;
 wire \device.rxBuffer.buffer[10][6] ;
 wire \device.rxBuffer.buffer[10][7] ;
 wire \device.rxBuffer.buffer[11][0] ;
 wire \device.rxBuffer.buffer[11][1] ;
 wire \device.rxBuffer.buffer[11][2] ;
 wire \device.rxBuffer.buffer[11][3] ;
 wire \device.rxBuffer.buffer[11][4] ;
 wire \device.rxBuffer.buffer[11][5] ;
 wire \device.rxBuffer.buffer[11][6] ;
 wire \device.rxBuffer.buffer[11][7] ;
 wire \device.rxBuffer.buffer[12][0] ;
 wire \device.rxBuffer.buffer[12][1] ;
 wire \device.rxBuffer.buffer[12][2] ;
 wire \device.rxBuffer.buffer[12][3] ;
 wire \device.rxBuffer.buffer[12][4] ;
 wire \device.rxBuffer.buffer[12][5] ;
 wire \device.rxBuffer.buffer[12][6] ;
 wire \device.rxBuffer.buffer[12][7] ;
 wire \device.rxBuffer.buffer[13][0] ;
 wire \device.rxBuffer.buffer[13][1] ;
 wire \device.rxBuffer.buffer[13][2] ;
 wire \device.rxBuffer.buffer[13][3] ;
 wire \device.rxBuffer.buffer[13][4] ;
 wire \device.rxBuffer.buffer[13][5] ;
 wire \device.rxBuffer.buffer[13][6] ;
 wire \device.rxBuffer.buffer[13][7] ;
 wire \device.rxBuffer.buffer[14][0] ;
 wire \device.rxBuffer.buffer[14][1] ;
 wire \device.rxBuffer.buffer[14][2] ;
 wire \device.rxBuffer.buffer[14][3] ;
 wire \device.rxBuffer.buffer[14][4] ;
 wire \device.rxBuffer.buffer[14][5] ;
 wire \device.rxBuffer.buffer[14][6] ;
 wire \device.rxBuffer.buffer[14][7] ;
 wire \device.rxBuffer.buffer[15][0] ;
 wire \device.rxBuffer.buffer[15][1] ;
 wire \device.rxBuffer.buffer[15][2] ;
 wire \device.rxBuffer.buffer[15][3] ;
 wire \device.rxBuffer.buffer[15][4] ;
 wire \device.rxBuffer.buffer[15][5] ;
 wire \device.rxBuffer.buffer[15][6] ;
 wire \device.rxBuffer.buffer[15][7] ;
 wire \device.rxBuffer.buffer[16][0] ;
 wire \device.rxBuffer.buffer[16][1] ;
 wire \device.rxBuffer.buffer[16][2] ;
 wire \device.rxBuffer.buffer[16][3] ;
 wire \device.rxBuffer.buffer[16][4] ;
 wire \device.rxBuffer.buffer[16][5] ;
 wire \device.rxBuffer.buffer[16][6] ;
 wire \device.rxBuffer.buffer[16][7] ;
 wire \device.rxBuffer.buffer[17][0] ;
 wire \device.rxBuffer.buffer[17][1] ;
 wire \device.rxBuffer.buffer[17][2] ;
 wire \device.rxBuffer.buffer[17][3] ;
 wire \device.rxBuffer.buffer[17][4] ;
 wire \device.rxBuffer.buffer[17][5] ;
 wire \device.rxBuffer.buffer[17][6] ;
 wire \device.rxBuffer.buffer[17][7] ;
 wire \device.rxBuffer.buffer[18][0] ;
 wire \device.rxBuffer.buffer[18][1] ;
 wire \device.rxBuffer.buffer[18][2] ;
 wire \device.rxBuffer.buffer[18][3] ;
 wire \device.rxBuffer.buffer[18][4] ;
 wire \device.rxBuffer.buffer[18][5] ;
 wire \device.rxBuffer.buffer[18][6] ;
 wire \device.rxBuffer.buffer[18][7] ;
 wire \device.rxBuffer.buffer[19][0] ;
 wire \device.rxBuffer.buffer[19][1] ;
 wire \device.rxBuffer.buffer[19][2] ;
 wire \device.rxBuffer.buffer[19][3] ;
 wire \device.rxBuffer.buffer[19][4] ;
 wire \device.rxBuffer.buffer[19][5] ;
 wire \device.rxBuffer.buffer[19][6] ;
 wire \device.rxBuffer.buffer[19][7] ;
 wire \device.rxBuffer.buffer[1][0] ;
 wire \device.rxBuffer.buffer[1][1] ;
 wire \device.rxBuffer.buffer[1][2] ;
 wire \device.rxBuffer.buffer[1][3] ;
 wire \device.rxBuffer.buffer[1][4] ;
 wire \device.rxBuffer.buffer[1][5] ;
 wire \device.rxBuffer.buffer[1][6] ;
 wire \device.rxBuffer.buffer[1][7] ;
 wire \device.rxBuffer.buffer[20][0] ;
 wire \device.rxBuffer.buffer[20][1] ;
 wire \device.rxBuffer.buffer[20][2] ;
 wire \device.rxBuffer.buffer[20][3] ;
 wire \device.rxBuffer.buffer[20][4] ;
 wire \device.rxBuffer.buffer[20][5] ;
 wire \device.rxBuffer.buffer[20][6] ;
 wire \device.rxBuffer.buffer[20][7] ;
 wire \device.rxBuffer.buffer[21][0] ;
 wire \device.rxBuffer.buffer[21][1] ;
 wire \device.rxBuffer.buffer[21][2] ;
 wire \device.rxBuffer.buffer[21][3] ;
 wire \device.rxBuffer.buffer[21][4] ;
 wire \device.rxBuffer.buffer[21][5] ;
 wire \device.rxBuffer.buffer[21][6] ;
 wire \device.rxBuffer.buffer[21][7] ;
 wire \device.rxBuffer.buffer[22][0] ;
 wire \device.rxBuffer.buffer[22][1] ;
 wire \device.rxBuffer.buffer[22][2] ;
 wire \device.rxBuffer.buffer[22][3] ;
 wire \device.rxBuffer.buffer[22][4] ;
 wire \device.rxBuffer.buffer[22][5] ;
 wire \device.rxBuffer.buffer[22][6] ;
 wire \device.rxBuffer.buffer[22][7] ;
 wire \device.rxBuffer.buffer[23][0] ;
 wire \device.rxBuffer.buffer[23][1] ;
 wire \device.rxBuffer.buffer[23][2] ;
 wire \device.rxBuffer.buffer[23][3] ;
 wire \device.rxBuffer.buffer[23][4] ;
 wire \device.rxBuffer.buffer[23][5] ;
 wire \device.rxBuffer.buffer[23][6] ;
 wire \device.rxBuffer.buffer[23][7] ;
 wire \device.rxBuffer.buffer[24][0] ;
 wire \device.rxBuffer.buffer[24][1] ;
 wire \device.rxBuffer.buffer[24][2] ;
 wire \device.rxBuffer.buffer[24][3] ;
 wire \device.rxBuffer.buffer[24][4] ;
 wire \device.rxBuffer.buffer[24][5] ;
 wire \device.rxBuffer.buffer[24][6] ;
 wire \device.rxBuffer.buffer[24][7] ;
 wire \device.rxBuffer.buffer[25][0] ;
 wire \device.rxBuffer.buffer[25][1] ;
 wire \device.rxBuffer.buffer[25][2] ;
 wire \device.rxBuffer.buffer[25][3] ;
 wire \device.rxBuffer.buffer[25][4] ;
 wire \device.rxBuffer.buffer[25][5] ;
 wire \device.rxBuffer.buffer[25][6] ;
 wire \device.rxBuffer.buffer[25][7] ;
 wire \device.rxBuffer.buffer[26][0] ;
 wire \device.rxBuffer.buffer[26][1] ;
 wire \device.rxBuffer.buffer[26][2] ;
 wire \device.rxBuffer.buffer[26][3] ;
 wire \device.rxBuffer.buffer[26][4] ;
 wire \device.rxBuffer.buffer[26][5] ;
 wire \device.rxBuffer.buffer[26][6] ;
 wire \device.rxBuffer.buffer[26][7] ;
 wire \device.rxBuffer.buffer[27][0] ;
 wire \device.rxBuffer.buffer[27][1] ;
 wire \device.rxBuffer.buffer[27][2] ;
 wire \device.rxBuffer.buffer[27][3] ;
 wire \device.rxBuffer.buffer[27][4] ;
 wire \device.rxBuffer.buffer[27][5] ;
 wire \device.rxBuffer.buffer[27][6] ;
 wire \device.rxBuffer.buffer[27][7] ;
 wire \device.rxBuffer.buffer[28][0] ;
 wire \device.rxBuffer.buffer[28][1] ;
 wire \device.rxBuffer.buffer[28][2] ;
 wire \device.rxBuffer.buffer[28][3] ;
 wire \device.rxBuffer.buffer[28][4] ;
 wire \device.rxBuffer.buffer[28][5] ;
 wire \device.rxBuffer.buffer[28][6] ;
 wire \device.rxBuffer.buffer[28][7] ;
 wire \device.rxBuffer.buffer[29][0] ;
 wire \device.rxBuffer.buffer[29][1] ;
 wire \device.rxBuffer.buffer[29][2] ;
 wire \device.rxBuffer.buffer[29][3] ;
 wire \device.rxBuffer.buffer[29][4] ;
 wire \device.rxBuffer.buffer[29][5] ;
 wire \device.rxBuffer.buffer[29][6] ;
 wire \device.rxBuffer.buffer[29][7] ;
 wire \device.rxBuffer.buffer[2][0] ;
 wire \device.rxBuffer.buffer[2][1] ;
 wire \device.rxBuffer.buffer[2][2] ;
 wire \device.rxBuffer.buffer[2][3] ;
 wire \device.rxBuffer.buffer[2][4] ;
 wire \device.rxBuffer.buffer[2][5] ;
 wire \device.rxBuffer.buffer[2][6] ;
 wire \device.rxBuffer.buffer[2][7] ;
 wire \device.rxBuffer.buffer[30][0] ;
 wire \device.rxBuffer.buffer[30][1] ;
 wire \device.rxBuffer.buffer[30][2] ;
 wire \device.rxBuffer.buffer[30][3] ;
 wire \device.rxBuffer.buffer[30][4] ;
 wire \device.rxBuffer.buffer[30][5] ;
 wire \device.rxBuffer.buffer[30][6] ;
 wire \device.rxBuffer.buffer[30][7] ;
 wire \device.rxBuffer.buffer[31][0] ;
 wire \device.rxBuffer.buffer[31][1] ;
 wire \device.rxBuffer.buffer[31][2] ;
 wire \device.rxBuffer.buffer[31][3] ;
 wire \device.rxBuffer.buffer[31][4] ;
 wire \device.rxBuffer.buffer[31][5] ;
 wire \device.rxBuffer.buffer[31][6] ;
 wire \device.rxBuffer.buffer[31][7] ;
 wire \device.rxBuffer.buffer[3][0] ;
 wire \device.rxBuffer.buffer[3][1] ;
 wire \device.rxBuffer.buffer[3][2] ;
 wire \device.rxBuffer.buffer[3][3] ;
 wire \device.rxBuffer.buffer[3][4] ;
 wire \device.rxBuffer.buffer[3][5] ;
 wire \device.rxBuffer.buffer[3][6] ;
 wire \device.rxBuffer.buffer[3][7] ;
 wire \device.rxBuffer.buffer[4][0] ;
 wire \device.rxBuffer.buffer[4][1] ;
 wire \device.rxBuffer.buffer[4][2] ;
 wire \device.rxBuffer.buffer[4][3] ;
 wire \device.rxBuffer.buffer[4][4] ;
 wire \device.rxBuffer.buffer[4][5] ;
 wire \device.rxBuffer.buffer[4][6] ;
 wire \device.rxBuffer.buffer[4][7] ;
 wire \device.rxBuffer.buffer[5][0] ;
 wire \device.rxBuffer.buffer[5][1] ;
 wire \device.rxBuffer.buffer[5][2] ;
 wire \device.rxBuffer.buffer[5][3] ;
 wire \device.rxBuffer.buffer[5][4] ;
 wire \device.rxBuffer.buffer[5][5] ;
 wire \device.rxBuffer.buffer[5][6] ;
 wire \device.rxBuffer.buffer[5][7] ;
 wire \device.rxBuffer.buffer[6][0] ;
 wire \device.rxBuffer.buffer[6][1] ;
 wire \device.rxBuffer.buffer[6][2] ;
 wire \device.rxBuffer.buffer[6][3] ;
 wire \device.rxBuffer.buffer[6][4] ;
 wire \device.rxBuffer.buffer[6][5] ;
 wire \device.rxBuffer.buffer[6][6] ;
 wire \device.rxBuffer.buffer[6][7] ;
 wire \device.rxBuffer.buffer[7][0] ;
 wire \device.rxBuffer.buffer[7][1] ;
 wire \device.rxBuffer.buffer[7][2] ;
 wire \device.rxBuffer.buffer[7][3] ;
 wire \device.rxBuffer.buffer[7][4] ;
 wire \device.rxBuffer.buffer[7][5] ;
 wire \device.rxBuffer.buffer[7][6] ;
 wire \device.rxBuffer.buffer[7][7] ;
 wire \device.rxBuffer.buffer[8][0] ;
 wire \device.rxBuffer.buffer[8][1] ;
 wire \device.rxBuffer.buffer[8][2] ;
 wire \device.rxBuffer.buffer[8][3] ;
 wire \device.rxBuffer.buffer[8][4] ;
 wire \device.rxBuffer.buffer[8][5] ;
 wire \device.rxBuffer.buffer[8][6] ;
 wire \device.rxBuffer.buffer[8][7] ;
 wire \device.rxBuffer.buffer[9][0] ;
 wire \device.rxBuffer.buffer[9][1] ;
 wire \device.rxBuffer.buffer[9][2] ;
 wire \device.rxBuffer.buffer[9][3] ;
 wire \device.rxBuffer.buffer[9][4] ;
 wire \device.rxBuffer.buffer[9][5] ;
 wire \device.rxBuffer.buffer[9][6] ;
 wire \device.rxBuffer.buffer[9][7] ;
 wire \device.rxBuffer.dataIn_buffered[0] ;
 wire \device.rxBuffer.dataIn_buffered[1] ;
 wire \device.rxBuffer.dataIn_buffered[2] ;
 wire \device.rxBuffer.dataIn_buffered[3] ;
 wire \device.rxBuffer.dataIn_buffered[4] ;
 wire \device.rxBuffer.dataIn_buffered[5] ;
 wire \device.rxBuffer.dataIn_buffered[6] ;
 wire \device.rxBuffer.dataIn_buffered[7] ;
 wire \device.rxBuffer.dataOut[0] ;
 wire \device.rxBuffer.dataOut[1] ;
 wire \device.rxBuffer.dataOut[2] ;
 wire \device.rxBuffer.dataOut[3] ;
 wire \device.rxBuffer.dataOut[4] ;
 wire \device.rxBuffer.dataOut[5] ;
 wire \device.rxBuffer.dataOut[6] ;
 wire \device.rxBuffer.dataOut[7] ;
 wire \device.rxBuffer.endPointer[0] ;
 wire \device.rxBuffer.endPointer[1] ;
 wire \device.rxBuffer.endPointer[2] ;
 wire \device.rxBuffer.endPointer[3] ;
 wire \device.rxBuffer.endPointer[4] ;
 wire \device.rxBuffer.lastWriteLostData ;
 wire \device.rxBuffer.oe_buffered ;
 wire \device.rxBuffer.startPointer[0] ;
 wire \device.rxBuffer.startPointer[1] ;
 wire \device.rxBuffer.startPointer[2] ;
 wire \device.rxBuffer.startPointer[3] ;
 wire \device.rxBuffer.startPointer[4] ;
 wire \device.rxBuffer.we_buffered ;
 wire \device.rxBufferFullBuffered ;
 wire \device.rxDataAvailableBuffered ;
 wire \device.rxDataLostBuffered ;
 wire \device.rxRegister.baseReadData[0] ;
 wire \device.rxRegister.baseReadData[1] ;
 wire \device.rxRegister.baseReadData[2] ;
 wire \device.rxRegister.baseReadData[3] ;
 wire \device.rxRegister.baseReadData[4] ;
 wire \device.rxRegister.baseReadData[5] ;
 wire \device.rxRegister.baseReadData[6] ;
 wire \device.rxRegister.baseReadData[7] ;
 wire \device.statusRegister.baseReadData[0] ;
 wire \device.statusRegister.baseReadData[1] ;
 wire \device.statusRegister.baseReadData[2] ;
 wire \device.statusRegister.baseReadData[3] ;
 wire \device.statusRegister.baseReadData[4] ;
 wire \device.statusRegister.baseReadData[5] ;
 wire \device.txBuffer.buffer[0][0] ;
 wire \device.txBuffer.buffer[0][1] ;
 wire \device.txBuffer.buffer[0][2] ;
 wire \device.txBuffer.buffer[0][3] ;
 wire \device.txBuffer.buffer[0][4] ;
 wire \device.txBuffer.buffer[0][5] ;
 wire \device.txBuffer.buffer[0][6] ;
 wire \device.txBuffer.buffer[0][7] ;
 wire \device.txBuffer.buffer[10][0] ;
 wire \device.txBuffer.buffer[10][1] ;
 wire \device.txBuffer.buffer[10][2] ;
 wire \device.txBuffer.buffer[10][3] ;
 wire \device.txBuffer.buffer[10][4] ;
 wire \device.txBuffer.buffer[10][5] ;
 wire \device.txBuffer.buffer[10][6] ;
 wire \device.txBuffer.buffer[10][7] ;
 wire \device.txBuffer.buffer[11][0] ;
 wire \device.txBuffer.buffer[11][1] ;
 wire \device.txBuffer.buffer[11][2] ;
 wire \device.txBuffer.buffer[11][3] ;
 wire \device.txBuffer.buffer[11][4] ;
 wire \device.txBuffer.buffer[11][5] ;
 wire \device.txBuffer.buffer[11][6] ;
 wire \device.txBuffer.buffer[11][7] ;
 wire \device.txBuffer.buffer[12][0] ;
 wire \device.txBuffer.buffer[12][1] ;
 wire \device.txBuffer.buffer[12][2] ;
 wire \device.txBuffer.buffer[12][3] ;
 wire \device.txBuffer.buffer[12][4] ;
 wire \device.txBuffer.buffer[12][5] ;
 wire \device.txBuffer.buffer[12][6] ;
 wire \device.txBuffer.buffer[12][7] ;
 wire \device.txBuffer.buffer[13][0] ;
 wire \device.txBuffer.buffer[13][1] ;
 wire \device.txBuffer.buffer[13][2] ;
 wire \device.txBuffer.buffer[13][3] ;
 wire \device.txBuffer.buffer[13][4] ;
 wire \device.txBuffer.buffer[13][5] ;
 wire \device.txBuffer.buffer[13][6] ;
 wire \device.txBuffer.buffer[13][7] ;
 wire \device.txBuffer.buffer[14][0] ;
 wire \device.txBuffer.buffer[14][1] ;
 wire \device.txBuffer.buffer[14][2] ;
 wire \device.txBuffer.buffer[14][3] ;
 wire \device.txBuffer.buffer[14][4] ;
 wire \device.txBuffer.buffer[14][5] ;
 wire \device.txBuffer.buffer[14][6] ;
 wire \device.txBuffer.buffer[14][7] ;
 wire \device.txBuffer.buffer[15][0] ;
 wire \device.txBuffer.buffer[15][1] ;
 wire \device.txBuffer.buffer[15][2] ;
 wire \device.txBuffer.buffer[15][3] ;
 wire \device.txBuffer.buffer[15][4] ;
 wire \device.txBuffer.buffer[15][5] ;
 wire \device.txBuffer.buffer[15][6] ;
 wire \device.txBuffer.buffer[15][7] ;
 wire \device.txBuffer.buffer[16][0] ;
 wire \device.txBuffer.buffer[16][1] ;
 wire \device.txBuffer.buffer[16][2] ;
 wire \device.txBuffer.buffer[16][3] ;
 wire \device.txBuffer.buffer[16][4] ;
 wire \device.txBuffer.buffer[16][5] ;
 wire \device.txBuffer.buffer[16][6] ;
 wire \device.txBuffer.buffer[16][7] ;
 wire \device.txBuffer.buffer[17][0] ;
 wire \device.txBuffer.buffer[17][1] ;
 wire \device.txBuffer.buffer[17][2] ;
 wire \device.txBuffer.buffer[17][3] ;
 wire \device.txBuffer.buffer[17][4] ;
 wire \device.txBuffer.buffer[17][5] ;
 wire \device.txBuffer.buffer[17][6] ;
 wire \device.txBuffer.buffer[17][7] ;
 wire \device.txBuffer.buffer[18][0] ;
 wire \device.txBuffer.buffer[18][1] ;
 wire \device.txBuffer.buffer[18][2] ;
 wire \device.txBuffer.buffer[18][3] ;
 wire \device.txBuffer.buffer[18][4] ;
 wire \device.txBuffer.buffer[18][5] ;
 wire \device.txBuffer.buffer[18][6] ;
 wire \device.txBuffer.buffer[18][7] ;
 wire \device.txBuffer.buffer[19][0] ;
 wire \device.txBuffer.buffer[19][1] ;
 wire \device.txBuffer.buffer[19][2] ;
 wire \device.txBuffer.buffer[19][3] ;
 wire \device.txBuffer.buffer[19][4] ;
 wire \device.txBuffer.buffer[19][5] ;
 wire \device.txBuffer.buffer[19][6] ;
 wire \device.txBuffer.buffer[19][7] ;
 wire \device.txBuffer.buffer[1][0] ;
 wire \device.txBuffer.buffer[1][1] ;
 wire \device.txBuffer.buffer[1][2] ;
 wire \device.txBuffer.buffer[1][3] ;
 wire \device.txBuffer.buffer[1][4] ;
 wire \device.txBuffer.buffer[1][5] ;
 wire \device.txBuffer.buffer[1][6] ;
 wire \device.txBuffer.buffer[1][7] ;
 wire \device.txBuffer.buffer[20][0] ;
 wire \device.txBuffer.buffer[20][1] ;
 wire \device.txBuffer.buffer[20][2] ;
 wire \device.txBuffer.buffer[20][3] ;
 wire \device.txBuffer.buffer[20][4] ;
 wire \device.txBuffer.buffer[20][5] ;
 wire \device.txBuffer.buffer[20][6] ;
 wire \device.txBuffer.buffer[20][7] ;
 wire \device.txBuffer.buffer[21][0] ;
 wire \device.txBuffer.buffer[21][1] ;
 wire \device.txBuffer.buffer[21][2] ;
 wire \device.txBuffer.buffer[21][3] ;
 wire \device.txBuffer.buffer[21][4] ;
 wire \device.txBuffer.buffer[21][5] ;
 wire \device.txBuffer.buffer[21][6] ;
 wire \device.txBuffer.buffer[21][7] ;
 wire \device.txBuffer.buffer[22][0] ;
 wire \device.txBuffer.buffer[22][1] ;
 wire \device.txBuffer.buffer[22][2] ;
 wire \device.txBuffer.buffer[22][3] ;
 wire \device.txBuffer.buffer[22][4] ;
 wire \device.txBuffer.buffer[22][5] ;
 wire \device.txBuffer.buffer[22][6] ;
 wire \device.txBuffer.buffer[22][7] ;
 wire \device.txBuffer.buffer[23][0] ;
 wire \device.txBuffer.buffer[23][1] ;
 wire \device.txBuffer.buffer[23][2] ;
 wire \device.txBuffer.buffer[23][3] ;
 wire \device.txBuffer.buffer[23][4] ;
 wire \device.txBuffer.buffer[23][5] ;
 wire \device.txBuffer.buffer[23][6] ;
 wire \device.txBuffer.buffer[23][7] ;
 wire \device.txBuffer.buffer[24][0] ;
 wire \device.txBuffer.buffer[24][1] ;
 wire \device.txBuffer.buffer[24][2] ;
 wire \device.txBuffer.buffer[24][3] ;
 wire \device.txBuffer.buffer[24][4] ;
 wire \device.txBuffer.buffer[24][5] ;
 wire \device.txBuffer.buffer[24][6] ;
 wire \device.txBuffer.buffer[24][7] ;
 wire \device.txBuffer.buffer[25][0] ;
 wire \device.txBuffer.buffer[25][1] ;
 wire \device.txBuffer.buffer[25][2] ;
 wire \device.txBuffer.buffer[25][3] ;
 wire \device.txBuffer.buffer[25][4] ;
 wire \device.txBuffer.buffer[25][5] ;
 wire \device.txBuffer.buffer[25][6] ;
 wire \device.txBuffer.buffer[25][7] ;
 wire \device.txBuffer.buffer[26][0] ;
 wire \device.txBuffer.buffer[26][1] ;
 wire \device.txBuffer.buffer[26][2] ;
 wire \device.txBuffer.buffer[26][3] ;
 wire \device.txBuffer.buffer[26][4] ;
 wire \device.txBuffer.buffer[26][5] ;
 wire \device.txBuffer.buffer[26][6] ;
 wire \device.txBuffer.buffer[26][7] ;
 wire \device.txBuffer.buffer[27][0] ;
 wire \device.txBuffer.buffer[27][1] ;
 wire \device.txBuffer.buffer[27][2] ;
 wire \device.txBuffer.buffer[27][3] ;
 wire \device.txBuffer.buffer[27][4] ;
 wire \device.txBuffer.buffer[27][5] ;
 wire \device.txBuffer.buffer[27][6] ;
 wire \device.txBuffer.buffer[27][7] ;
 wire \device.txBuffer.buffer[28][0] ;
 wire \device.txBuffer.buffer[28][1] ;
 wire \device.txBuffer.buffer[28][2] ;
 wire \device.txBuffer.buffer[28][3] ;
 wire \device.txBuffer.buffer[28][4] ;
 wire \device.txBuffer.buffer[28][5] ;
 wire \device.txBuffer.buffer[28][6] ;
 wire \device.txBuffer.buffer[28][7] ;
 wire \device.txBuffer.buffer[29][0] ;
 wire \device.txBuffer.buffer[29][1] ;
 wire \device.txBuffer.buffer[29][2] ;
 wire \device.txBuffer.buffer[29][3] ;
 wire \device.txBuffer.buffer[29][4] ;
 wire \device.txBuffer.buffer[29][5] ;
 wire \device.txBuffer.buffer[29][6] ;
 wire \device.txBuffer.buffer[29][7] ;
 wire \device.txBuffer.buffer[2][0] ;
 wire \device.txBuffer.buffer[2][1] ;
 wire \device.txBuffer.buffer[2][2] ;
 wire \device.txBuffer.buffer[2][3] ;
 wire \device.txBuffer.buffer[2][4] ;
 wire \device.txBuffer.buffer[2][5] ;
 wire \device.txBuffer.buffer[2][6] ;
 wire \device.txBuffer.buffer[2][7] ;
 wire \device.txBuffer.buffer[30][0] ;
 wire \device.txBuffer.buffer[30][1] ;
 wire \device.txBuffer.buffer[30][2] ;
 wire \device.txBuffer.buffer[30][3] ;
 wire \device.txBuffer.buffer[30][4] ;
 wire \device.txBuffer.buffer[30][5] ;
 wire \device.txBuffer.buffer[30][6] ;
 wire \device.txBuffer.buffer[30][7] ;
 wire \device.txBuffer.buffer[31][0] ;
 wire \device.txBuffer.buffer[31][1] ;
 wire \device.txBuffer.buffer[31][2] ;
 wire \device.txBuffer.buffer[31][3] ;
 wire \device.txBuffer.buffer[31][4] ;
 wire \device.txBuffer.buffer[31][5] ;
 wire \device.txBuffer.buffer[31][6] ;
 wire \device.txBuffer.buffer[31][7] ;
 wire \device.txBuffer.buffer[3][0] ;
 wire \device.txBuffer.buffer[3][1] ;
 wire \device.txBuffer.buffer[3][2] ;
 wire \device.txBuffer.buffer[3][3] ;
 wire \device.txBuffer.buffer[3][4] ;
 wire \device.txBuffer.buffer[3][5] ;
 wire \device.txBuffer.buffer[3][6] ;
 wire \device.txBuffer.buffer[3][7] ;
 wire \device.txBuffer.buffer[4][0] ;
 wire \device.txBuffer.buffer[4][1] ;
 wire \device.txBuffer.buffer[4][2] ;
 wire \device.txBuffer.buffer[4][3] ;
 wire \device.txBuffer.buffer[4][4] ;
 wire \device.txBuffer.buffer[4][5] ;
 wire \device.txBuffer.buffer[4][6] ;
 wire \device.txBuffer.buffer[4][7] ;
 wire \device.txBuffer.buffer[5][0] ;
 wire \device.txBuffer.buffer[5][1] ;
 wire \device.txBuffer.buffer[5][2] ;
 wire \device.txBuffer.buffer[5][3] ;
 wire \device.txBuffer.buffer[5][4] ;
 wire \device.txBuffer.buffer[5][5] ;
 wire \device.txBuffer.buffer[5][6] ;
 wire \device.txBuffer.buffer[5][7] ;
 wire \device.txBuffer.buffer[6][0] ;
 wire \device.txBuffer.buffer[6][1] ;
 wire \device.txBuffer.buffer[6][2] ;
 wire \device.txBuffer.buffer[6][3] ;
 wire \device.txBuffer.buffer[6][4] ;
 wire \device.txBuffer.buffer[6][5] ;
 wire \device.txBuffer.buffer[6][6] ;
 wire \device.txBuffer.buffer[6][7] ;
 wire \device.txBuffer.buffer[7][0] ;
 wire \device.txBuffer.buffer[7][1] ;
 wire \device.txBuffer.buffer[7][2] ;
 wire \device.txBuffer.buffer[7][3] ;
 wire \device.txBuffer.buffer[7][4] ;
 wire \device.txBuffer.buffer[7][5] ;
 wire \device.txBuffer.buffer[7][6] ;
 wire \device.txBuffer.buffer[7][7] ;
 wire \device.txBuffer.buffer[8][0] ;
 wire \device.txBuffer.buffer[8][1] ;
 wire \device.txBuffer.buffer[8][2] ;
 wire \device.txBuffer.buffer[8][3] ;
 wire \device.txBuffer.buffer[8][4] ;
 wire \device.txBuffer.buffer[8][5] ;
 wire \device.txBuffer.buffer[8][6] ;
 wire \device.txBuffer.buffer[8][7] ;
 wire \device.txBuffer.buffer[9][0] ;
 wire \device.txBuffer.buffer[9][1] ;
 wire \device.txBuffer.buffer[9][2] ;
 wire \device.txBuffer.buffer[9][3] ;
 wire \device.txBuffer.buffer[9][4] ;
 wire \device.txBuffer.buffer[9][5] ;
 wire \device.txBuffer.buffer[9][6] ;
 wire \device.txBuffer.buffer[9][7] ;
 wire \device.txBuffer.dataIn_buffered[0] ;
 wire \device.txBuffer.dataIn_buffered[1] ;
 wire \device.txBuffer.dataIn_buffered[2] ;
 wire \device.txBuffer.dataIn_buffered[3] ;
 wire \device.txBuffer.dataIn_buffered[4] ;
 wire \device.txBuffer.dataIn_buffered[5] ;
 wire \device.txBuffer.dataIn_buffered[6] ;
 wire \device.txBuffer.dataIn_buffered[7] ;
 wire \device.txBuffer.dataOut[0] ;
 wire \device.txBuffer.dataOut[1] ;
 wire \device.txBuffer.dataOut[2] ;
 wire \device.txBuffer.dataOut[3] ;
 wire \device.txBuffer.dataOut[4] ;
 wire \device.txBuffer.dataOut[5] ;
 wire \device.txBuffer.dataOut[6] ;
 wire \device.txBuffer.dataOut[7] ;
 wire \device.txBuffer.endPointer[0] ;
 wire \device.txBuffer.endPointer[1] ;
 wire \device.txBuffer.endPointer[2] ;
 wire \device.txBuffer.endPointer[3] ;
 wire \device.txBuffer.endPointer[4] ;
 wire \device.txBuffer.lastWriteLostData ;
 wire \device.txBuffer.oe_buffered ;
 wire \device.txBuffer.startPointer[0] ;
 wire \device.txBuffer.startPointer[1] ;
 wire \device.txBuffer.startPointer[2] ;
 wire \device.txBuffer.startPointer[3] ;
 wire \device.txBuffer.startPointer[4] ;
 wire \device.txBuffer.we_buffered ;
 wire \device.txBufferFullBuffered ;
 wire \device.txDataAvailableBuffered ;
 wire \device.txDataLostBuffered ;
 wire \device.txSendBusy ;
 wire \device.uartRx.bitCounter[0] ;
 wire \device.uartRx.bitCounter[1] ;
 wire \device.uartRx.bitCounter[2] ;
 wire \device.uartRx.delayCounter[0] ;
 wire \device.uartRx.delayCounter[10] ;
 wire \device.uartRx.delayCounter[11] ;
 wire \device.uartRx.delayCounter[12] ;
 wire \device.uartRx.delayCounter[13] ;
 wire \device.uartRx.delayCounter[14] ;
 wire \device.uartRx.delayCounter[15] ;
 wire \device.uartRx.delayCounter[1] ;
 wire \device.uartRx.delayCounter[2] ;
 wire \device.uartRx.delayCounter[3] ;
 wire \device.uartRx.delayCounter[4] ;
 wire \device.uartRx.delayCounter[5] ;
 wire \device.uartRx.delayCounter[6] ;
 wire \device.uartRx.delayCounter[7] ;
 wire \device.uartRx.delayCounter[8] ;
 wire \device.uartRx.delayCounter[9] ;
 wire \device.uartRx.newData ;
 wire \device.uartRx.savedData[0] ;
 wire \device.uartRx.savedData[1] ;
 wire \device.uartRx.savedData[2] ;
 wire \device.uartRx.savedData[3] ;
 wire \device.uartRx.savedData[4] ;
 wire \device.uartRx.savedData[5] ;
 wire \device.uartRx.savedData[6] ;
 wire \device.uartRx.savedData[7] ;
 wire \device.uartRx.state[0] ;
 wire \device.uartRx.state[1] ;
 wire \device.uartTx.bitCounter[0] ;
 wire \device.uartTx.bitCounter[1] ;
 wire \device.uartTx.bitCounter[2] ;
 wire \device.uartTx.delayCounter[0] ;
 wire \device.uartTx.delayCounter[10] ;
 wire \device.uartTx.delayCounter[11] ;
 wire \device.uartTx.delayCounter[12] ;
 wire \device.uartTx.delayCounter[13] ;
 wire \device.uartTx.delayCounter[14] ;
 wire \device.uartTx.delayCounter[15] ;
 wire \device.uartTx.delayCounter[1] ;
 wire \device.uartTx.delayCounter[2] ;
 wire \device.uartTx.delayCounter[3] ;
 wire \device.uartTx.delayCounter[4] ;
 wire \device.uartTx.delayCounter[5] ;
 wire \device.uartTx.delayCounter[6] ;
 wire \device.uartTx.delayCounter[7] ;
 wire \device.uartTx.delayCounter[8] ;
 wire \device.uartTx.delayCounter[9] ;
 wire \device.uartTx.savedData[0] ;
 wire \device.uartTx.savedData[1] ;
 wire \device.uartTx.savedData[2] ;
 wire \device.uartTx.savedData[3] ;
 wire \device.uartTx.savedData[4] ;
 wire \device.uartTx.savedData[5] ;
 wire \device.uartTx.savedData[6] ;
 wire \device.uartTx.savedData[7] ;
 wire \device.uartTx.state[0] ;
 wire \device.uartTx.state[1] ;
 wire hostConfigLatch;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net152;
 wire net1521;
 wire net1524;
 wire net1526;
 wire net1527;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1534;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1543;
 wire net1546;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1608;
 wire net1609;
 wire net161;
 wire net162;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1648;
 wire net165;
 wire net1652;
 wire net1653;
 wire net1655;
 wire net1658;
 wire net166;
 wire net1660;
 wire net1664;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1689;
 wire net169;
 wire net1696;
 wire net1697;
 wire net17;
 wire net170;
 wire net1706;
 wire net1707;
 wire net171;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1718;
 wire net172;
 wire net1722;
 wire net1726;
 wire net173;
 wire net1730;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1744;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1755;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1774;
 wire net1775;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net179;
 wire net1793;
 wire net1798;
 wire net18;
 wire net180;
 wire net1802;
 wire net1803;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net181;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net182;
 wire net1822;
 wire net1823;
 wire net1829;
 wire net183;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net184;
 wire net1841;
 wire net1842;
 wire net185;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1865;
 wire net1866;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net188;
 wire net1880;
 wire net189;
 wire net19;
 wire net190;
 wire net1909;
 wire net191;
 wire net192;
 wire net1922;
 wire net193;
 wire net194;
 wire net1943;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net196;
 wire net1963;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1977;
 wire net198;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1998;
 wire net2;
 wire net20;
 wire net200;
 wire net2004;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2029;
 wire net203;
 wire net2035;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2047;
 wire net205;
 wire net2055;
 wire net206;
 wire net2063;
 wire net2067;
 wire net2068;
 wire net207;
 wire net2074;
 wire net208;
 wire net2080;
 wire net2084;
 wire net2085;
 wire net209;
 wire net2091;
 wire net2097;
 wire net21;
 wire net210;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net211;
 wire net2114;
 wire net212;
 wire net2122;
 wire net2123;
 wire net2129;
 wire net213;
 wire net2133;
 wire net2134;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2143;
 wire net2144;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net216;
 wire net2160;
 wire net217;
 wire net218;
 wire net2184;
 wire net219;
 wire net2190;
 wire net22;
 wire net220;
 wire net221;
 wire net2210;
 wire net222;
 wire net223;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2346;
 wire net2347;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2366;
 wire net2367;
 wire net237;
 wire net2373;
 wire net2374;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2387;
 wire net2388;
 wire net239;
 wire net2394;
 wire net2395;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net241;
 wire net2413;
 wire net2414;
 wire net242;
 wire net2420;
 wire net2421;
 wire net243;
 wire net2432;
 wire net2433;
 wire net2438;
 wire net2439;
 wire net244;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net245;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net246;
 wire net2460;
 wire net2466;
 wire net2467;
 wire net247;
 wire net2473;
 wire net2474;
 wire net2478;
 wire net2479;
 wire net248;
 wire net2480;
 wire net2481;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net249;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2499;
 wire net25;
 wire net250;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net251;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net252;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2528;
 wire net2529;
 wire net253;
 wire net2535;
 wire net2536;
 wire net254;
 wire net2542;
 wire net2543;
 wire net2549;
 wire net255;
 wire net2550;
 wire net2556;
 wire net2557;
 wire net256;
 wire net2563;
 wire net2564;
 wire net257;
 wire net2570;
 wire net2571;
 wire net2574;
 wire net2575;
 wire net2579;
 wire net258;
 wire net2580;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net259;
 wire net2595;
 wire net2596;
 wire net26;
 wire net260;
 wire net2604;
 wire net2605;
 wire net2608;
 wire net2609;
 wire net261;
 wire net2612;
 wire net2613;
 wire net2616;
 wire net2617;
 wire net262;
 wire net2620;
 wire net2621;
 wire net2624;
 wire net2625;
 wire net263;
 wire net2633;
 wire net2634;
 wire net2637;
 wire net2638;
 wire net264;
 wire net2641;
 wire net2642;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net265;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net266;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net267;
 wire net2670;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net268;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net269;
 wire net2694;
 wire net2695;
 wire net2699;
 wire net27;
 wire net270;
 wire net2700;
 wire net2704;
 wire net2705;
 wire net2709;
 wire net271;
 wire net2710;
 wire net2714;
 wire net2715;
 wire net2719;
 wire net272;
 wire net2720;
 wire net2724;
 wire net2725;
 wire net2728;
 wire net2729;
 wire net273;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2736;
 wire net2737;
 wire net274;
 wire net2740;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net275;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net276;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net277;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net278;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net279;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net28;
 wire net280;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net281;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net282;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net283;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net284;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net285;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net286;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net287;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net288;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net289;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net29;
 wire net290;
 wire net2900;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2909;
 wire net291;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net292;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net293;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2938;
 wire net2939;
 wire net294;
 wire net2940;
 wire net2941;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net295;
 wire net2950;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net296;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net297;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net298;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net299;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2999;
 wire net3;
 wire net30;
 wire net300;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3008;
 wire net3009;
 wire net301;
 wire net3010;
 wire net3011;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net302;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net303;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net304;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net305;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net306;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net307;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3079;
 wire net308;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3088;
 wire net3089;
 wire net309;
 wire net3090;
 wire net3091;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net31;
 wire net310;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net311;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net312;
 wire net3120;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net313;
 wire net3130;
 wire net3131;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net314;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net315;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net316;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net317;
 wire net3170;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net318;
 wire net3180;
 wire net3181;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net319;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net32;
 wire net320;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net321;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3218;
 wire net3219;
 wire net322;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3229;
 wire net323;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net324;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net325;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net326;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net327;
 wire net3270;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3279;
 wire net328;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net329;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net33;
 wire net330;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3308;
 wire net3309;
 wire net331;
 wire net3310;
 wire net3311;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net332;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net333;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net334;
 wire net3340;
 wire net3348;
 wire net3349;
 wire net335;
 wire net3350;
 wire net3351;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net336;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3369;
 wire net337;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net338;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net339;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net34;
 wire net340;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net341;
 wire net3410;
 wire net3411;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net342;
 wire net3420;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net343;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net344;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net345;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net346;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net347;
 wire net3470;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net348;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net349;
 wire net3490;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net35;
 wire net350;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net351;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net352;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net353;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net354;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net355;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net356;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net357;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net358;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net359;
 wire net3590;
 wire net3591;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net36;
 wire net360;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net361;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net362;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net363;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net364;
 wire net3640;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net365;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3659;
 wire net366;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net367;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net368;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net369;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net37;
 wire net370;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net371;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net372;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net373;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net374;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net375;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net376;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net377;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3778;
 wire net3779;
 wire net378;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net379;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net38;
 wire net380;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net381;
 wire net3810;
 wire net3811;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net382;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net383;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net384;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net385;
 wire net3850;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net386;
 wire net3860;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net387;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net388;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net389;
 wire net3890;
 wire net3898;
 wire net3899;
 wire net39;
 wire net390;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net391;
 wire net3910;
 wire net3911;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net392;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net393;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net394;
 wire net3940;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net395;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3959;
 wire net396;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net397;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net398;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net399;
 wire net3990;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3998;
 wire net4;
 wire net40;
 wire net400;
 wire net4001;
 wire net401;
 wire net4011;
 wire net4012;
 wire net4016;
 wire net4017;
 wire net402;
 wire net4020;
 wire net4021;
 wire net4025;
 wire net4029;
 wire net403;
 wire net4033;
 wire net4037;
 wire net404;
 wire net4041;
 wire net4045;
 wire net4049;
 wire net405;
 wire net4053;
 wire net4059;
 wire net406;
 wire net4068;
 wire net4069;
 wire net407;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net408;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net409;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net41;
 wire net410;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4106;
 wire net4107;
 wire net411;
 wire net4112;
 wire net4113;
 wire net4119;
 wire net412;
 wire net4125;
 wire net413;
 wire net4131;
 wire net4137;
 wire net414;
 wire net4143;
 wire net4149;
 wire net415;
 wire net4150;
 wire net4156;
 wire net416;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net417;
 wire net4170;
 wire net4171;
 wire net4174;
 wire net4175;
 wire net4178;
 wire net4179;
 wire net418;
 wire net4180;
 wire net4181;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \wbAddressExtension.acknowledge ;
 wire \wbAddressExtension.currentAddress[0] ;
 wire \wbAddressExtension.currentAddress[10] ;
 wire \wbAddressExtension.currentAddress[11] ;
 wire \wbAddressExtension.currentAddress[12] ;
 wire \wbAddressExtension.currentAddress[13] ;
 wire \wbAddressExtension.currentAddress[14] ;
 wire \wbAddressExtension.currentAddress[15] ;
 wire \wbAddressExtension.currentAddress[16] ;
 wire \wbAddressExtension.currentAddress[17] ;
 wire \wbAddressExtension.currentAddress[18] ;
 wire \wbAddressExtension.currentAddress[19] ;
 wire \wbAddressExtension.currentAddress[1] ;
 wire \wbAddressExtension.currentAddress[20] ;
 wire \wbAddressExtension.currentAddress[21] ;
 wire \wbAddressExtension.currentAddress[22] ;
 wire \wbAddressExtension.currentAddress[23] ;
 wire \wbAddressExtension.currentAddress[24] ;
 wire \wbAddressExtension.currentAddress[25] ;
 wire \wbAddressExtension.currentAddress[26] ;
 wire \wbAddressExtension.currentAddress[27] ;
 wire \wbAddressExtension.currentAddress[28] ;
 wire \wbAddressExtension.currentAddress[29] ;
 wire \wbAddressExtension.currentAddress[2] ;
 wire \wbAddressExtension.currentAddress[30] ;
 wire \wbAddressExtension.currentAddress[31] ;
 wire \wbAddressExtension.currentAddress[3] ;
 wire \wbAddressExtension.currentAddress[4] ;
 wire \wbAddressExtension.currentAddress[5] ;
 wire \wbAddressExtension.currentAddress[6] ;
 wire \wbAddressExtension.currentAddress[7] ;
 wire \wbAddressExtension.currentAddress[8] ;
 wire \wbAddressExtension.currentAddress[9] ;
 wire \wbAddressExtension.dataRead_buffered[0] ;
 wire \wbAddressExtension.dataRead_buffered[10] ;
 wire \wbAddressExtension.dataRead_buffered[11] ;
 wire \wbAddressExtension.dataRead_buffered[12] ;
 wire \wbAddressExtension.dataRead_buffered[13] ;
 wire \wbAddressExtension.dataRead_buffered[14] ;
 wire \wbAddressExtension.dataRead_buffered[15] ;
 wire \wbAddressExtension.dataRead_buffered[16] ;
 wire \wbAddressExtension.dataRead_buffered[17] ;
 wire \wbAddressExtension.dataRead_buffered[18] ;
 wire \wbAddressExtension.dataRead_buffered[19] ;
 wire \wbAddressExtension.dataRead_buffered[1] ;
 wire \wbAddressExtension.dataRead_buffered[20] ;
 wire \wbAddressExtension.dataRead_buffered[21] ;
 wire \wbAddressExtension.dataRead_buffered[22] ;
 wire \wbAddressExtension.dataRead_buffered[23] ;
 wire \wbAddressExtension.dataRead_buffered[24] ;
 wire \wbAddressExtension.dataRead_buffered[25] ;
 wire \wbAddressExtension.dataRead_buffered[26] ;
 wire \wbAddressExtension.dataRead_buffered[27] ;
 wire \wbAddressExtension.dataRead_buffered[28] ;
 wire \wbAddressExtension.dataRead_buffered[29] ;
 wire \wbAddressExtension.dataRead_buffered[2] ;
 wire \wbAddressExtension.dataRead_buffered[30] ;
 wire \wbAddressExtension.dataRead_buffered[31] ;
 wire \wbAddressExtension.dataRead_buffered[3] ;
 wire \wbAddressExtension.dataRead_buffered[4] ;
 wire \wbAddressExtension.dataRead_buffered[5] ;
 wire \wbAddressExtension.dataRead_buffered[6] ;
 wire \wbAddressExtension.dataRead_buffered[7] ;
 wire \wbAddressExtension.dataRead_buffered[8] ;
 wire \wbAddressExtension.dataRead_buffered[9] ;
 wire \wbAddressExtension.state[0] ;
 wire \wbAddressExtension.state[1] ;
 wire \wbPeripheralBusInterface.acknowledge ;
 wire \wbPeripheralBusInterface.currentAddress[10] ;
 wire \wbPeripheralBusInterface.currentAddress[11] ;
 wire \wbPeripheralBusInterface.currentAddress[12] ;
 wire \wbPeripheralBusInterface.currentAddress[13] ;
 wire \wbPeripheralBusInterface.currentAddress[14] ;
 wire \wbPeripheralBusInterface.currentAddress[15] ;
 wire \wbPeripheralBusInterface.currentAddress[16] ;
 wire \wbPeripheralBusInterface.currentAddress[17] ;
 wire \wbPeripheralBusInterface.currentAddress[18] ;
 wire \wbPeripheralBusInterface.currentAddress[19] ;
 wire \wbPeripheralBusInterface.currentAddress[20] ;
 wire \wbPeripheralBusInterface.currentAddress[21] ;
 wire \wbPeripheralBusInterface.currentAddress[22] ;
 wire \wbPeripheralBusInterface.currentAddress[23] ;
 wire \wbPeripheralBusInterface.currentAddress[2] ;
 wire \wbPeripheralBusInterface.currentAddress[3] ;
 wire \wbPeripheralBusInterface.currentAddress[4] ;
 wire \wbPeripheralBusInterface.currentAddress[5] ;
 wire \wbPeripheralBusInterface.currentAddress[6] ;
 wire \wbPeripheralBusInterface.currentAddress[7] ;
 wire \wbPeripheralBusInterface.currentAddress[8] ;
 wire \wbPeripheralBusInterface.currentAddress[9] ;
 wire \wbPeripheralBusInterface.currentByteSelect[0] ;
 wire \wbPeripheralBusInterface.currentByteSelect[1] ;
 wire \wbPeripheralBusInterface.currentByteSelect[2] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[0] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[10] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[11] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[12] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[13] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[14] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[15] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[16] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[17] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[18] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[19] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[1] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[20] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[21] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[2] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[3] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[4] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[5] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[6] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[7] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[8] ;
 wire \wbPeripheralBusInterface.dataRead_buffered[9] ;
 wire \wbPeripheralBusInterface.state[0] ;
 wire \wbPeripheralBusInterface.state[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(wbs_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(wbs_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(wbs_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net2796));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net2853));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net3530));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net3542));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net3550));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net3713));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_1781_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_1808_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\device.txDataAvailableBuffered ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\wbPeripheralBusInterface.currentByteSelect[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(wbs_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(wbs_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(wbs_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1980_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net1283));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net2261));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net3520));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net3548));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net3672));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\device.rxBuffer.dataIn_buffered[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\device.rxBuffer.dataIn_buffered[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\device.txBuffer.dataIn_buffered[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(wbs_adr_i[3]));
 sky130_fd_sc_hd__conb_1 CaravelHost_651 (.LO(net651));
 sky130_fd_sc_hd__conb_1 CaravelHost_652 (.LO(net652));
 sky130_fd_sc_hd__conb_1 CaravelHost_653 (.LO(net653));
 sky130_fd_sc_hd__conb_1 CaravelHost_654 (.LO(net654));
 sky130_fd_sc_hd__conb_1 CaravelHost_655 (.LO(net655));
 sky130_fd_sc_hd__conb_1 CaravelHost_656 (.LO(net656));
 sky130_fd_sc_hd__conb_1 CaravelHost_657 (.LO(net657));
 sky130_fd_sc_hd__conb_1 CaravelHost_658 (.LO(net658));
 sky130_fd_sc_hd__conb_1 CaravelHost_659 (.LO(net659));
 sky130_fd_sc_hd__conb_1 CaravelHost_660 (.LO(net660));
 sky130_fd_sc_hd__conb_1 CaravelHost_661 (.LO(net661));
 sky130_fd_sc_hd__conb_1 CaravelHost_662 (.LO(net662));
 sky130_fd_sc_hd__conb_1 CaravelHost_663 (.LO(net663));
 sky130_fd_sc_hd__conb_1 CaravelHost_664 (.LO(net664));
 sky130_fd_sc_hd__conb_1 CaravelHost_665 (.LO(net665));
 sky130_fd_sc_hd__conb_1 CaravelHost_666 (.LO(net666));
 sky130_fd_sc_hd__conb_1 CaravelHost_667 (.LO(net667));
 sky130_fd_sc_hd__conb_1 CaravelHost_668 (.LO(net668));
 sky130_fd_sc_hd__conb_1 CaravelHost_669 (.LO(net669));
 sky130_fd_sc_hd__conb_1 CaravelHost_670 (.LO(net670));
 sky130_fd_sc_hd__conb_1 CaravelHost_671 (.LO(net671));
 sky130_fd_sc_hd__conb_1 CaravelHost_672 (.LO(net672));
 sky130_fd_sc_hd__conb_1 CaravelHost_673 (.LO(net673));
 sky130_fd_sc_hd__conb_1 CaravelHost_674 (.LO(net674));
 sky130_fd_sc_hd__conb_1 CaravelHost_675 (.LO(net675));
 sky130_fd_sc_hd__conb_1 CaravelHost_676 (.LO(net676));
 sky130_fd_sc_hd__conb_1 CaravelHost_677 (.LO(net677));
 sky130_fd_sc_hd__conb_1 CaravelHost_678 (.LO(net678));
 sky130_fd_sc_hd__conb_1 CaravelHost_679 (.LO(net679));
 sky130_fd_sc_hd__conb_1 CaravelHost_680 (.LO(net680));
 sky130_fd_sc_hd__conb_1 CaravelHost_681 (.LO(net681));
 sky130_fd_sc_hd__conb_1 CaravelHost_682 (.LO(net682));
 sky130_fd_sc_hd__conb_1 CaravelHost_683 (.LO(net683));
 sky130_fd_sc_hd__conb_1 CaravelHost_684 (.LO(net684));
 sky130_fd_sc_hd__conb_1 CaravelHost_685 (.LO(net685));
 sky130_fd_sc_hd__conb_1 CaravelHost_686 (.LO(net686));
 sky130_fd_sc_hd__conb_1 CaravelHost_687 (.LO(net687));
 sky130_fd_sc_hd__conb_1 CaravelHost_688 (.LO(net688));
 sky130_fd_sc_hd__conb_1 CaravelHost_689 (.LO(net689));
 sky130_fd_sc_hd__conb_1 CaravelHost_690 (.LO(net690));
 sky130_fd_sc_hd__conb_1 CaravelHost_691 (.LO(net691));
 sky130_fd_sc_hd__conb_1 CaravelHost_692 (.LO(net692));
 sky130_fd_sc_hd__conb_1 CaravelHost_693 (.LO(net693));
 sky130_fd_sc_hd__conb_1 CaravelHost_694 (.LO(net694));
 sky130_fd_sc_hd__conb_1 CaravelHost_695 (.LO(net695));
 sky130_fd_sc_hd__conb_1 CaravelHost_696 (.LO(net696));
 sky130_fd_sc_hd__conb_1 CaravelHost_697 (.LO(net697));
 sky130_fd_sc_hd__conb_1 CaravelHost_698 (.LO(net698));
 sky130_fd_sc_hd__conb_1 CaravelHost_699 (.LO(net699));
 sky130_fd_sc_hd__conb_1 CaravelHost_700 (.LO(net700));
 sky130_fd_sc_hd__conb_1 CaravelHost_701 (.LO(net701));
 sky130_fd_sc_hd__conb_1 CaravelHost_702 (.LO(net702));
 sky130_fd_sc_hd__conb_1 CaravelHost_703 (.LO(net703));
 sky130_fd_sc_hd__conb_1 CaravelHost_704 (.LO(net704));
 sky130_fd_sc_hd__conb_1 CaravelHost_705 (.LO(net705));
 sky130_fd_sc_hd__conb_1 CaravelHost_706 (.LO(net706));
 sky130_fd_sc_hd__conb_1 CaravelHost_707 (.LO(net707));
 sky130_fd_sc_hd__conb_1 CaravelHost_708 (.LO(net708));
 sky130_fd_sc_hd__conb_1 CaravelHost_709 (.LO(net709));
 sky130_fd_sc_hd__conb_1 CaravelHost_710 (.LO(net710));
 sky130_fd_sc_hd__conb_1 CaravelHost_711 (.LO(net711));
 sky130_fd_sc_hd__conb_1 CaravelHost_712 (.LO(net712));
 sky130_fd_sc_hd__conb_1 CaravelHost_713 (.LO(net713));
 sky130_fd_sc_hd__conb_1 CaravelHost_714 (.LO(net714));
 sky130_fd_sc_hd__conb_1 CaravelHost_715 (.LO(net715));
 sky130_fd_sc_hd__conb_1 CaravelHost_716 (.LO(net716));
 sky130_fd_sc_hd__conb_1 CaravelHost_717 (.LO(net717));
 sky130_fd_sc_hd__conb_1 CaravelHost_718 (.LO(net718));
 sky130_fd_sc_hd__conb_1 CaravelHost_719 (.LO(net719));
 sky130_fd_sc_hd__conb_1 CaravelHost_720 (.LO(net720));
 sky130_fd_sc_hd__conb_1 CaravelHost_721 (.LO(net721));
 sky130_fd_sc_hd__conb_1 CaravelHost_722 (.HI(net722));
 sky130_fd_sc_hd__conb_1 CaravelHost_723 (.HI(net723));
 sky130_fd_sc_hd__conb_1 CaravelHost_724 (.HI(net724));
 sky130_fd_sc_hd__conb_1 CaravelHost_725 (.HI(net725));
 sky130_fd_sc_hd__conb_1 CaravelHost_726 (.HI(net726));
 sky130_fd_sc_hd__conb_1 CaravelHost_727 (.HI(net727));
 sky130_fd_sc_hd__conb_1 CaravelHost_728 (.HI(net728));
 sky130_fd_sc_hd__conb_1 CaravelHost_729 (.HI(net729));
 sky130_fd_sc_hd__conb_1 CaravelHost_730 (.HI(net730));
 sky130_fd_sc_hd__conb_1 CaravelHost_731 (.HI(net731));
 sky130_fd_sc_hd__fill_2 FILLER_0_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_94 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkinv_4 _2433_ (.A(\device.configuration[7] ),
    .Y(_1340_));
 sky130_fd_sc_hd__inv_2 _2434_ (.A(\device.configuration[14] ),
    .Y(_1341_));
 sky130_fd_sc_hd__inv_2 _2435_ (.A(\device.configuration[16] ),
    .Y(_1342_));
 sky130_fd_sc_hd__inv_2 _2436_ (.A(\device.configuration[17] ),
    .Y(_1343_));
 sky130_fd_sc_hd__inv_2 _2437_ (.A(\device.uartRx.bitCounter[2] ),
    .Y(_1344_));
 sky130_fd_sc_hd__inv_2 _2438_ (.A(\device.uartRx.bitCounter[0] ),
    .Y(_1345_));
 sky130_fd_sc_hd__inv_2 _2439_ (.A(\device.uartRx.delayCounter[14] ),
    .Y(_1346_));
 sky130_fd_sc_hd__inv_2 _2440_ (.A(\device.uartRx.delayCounter[13] ),
    .Y(_1347_));
 sky130_fd_sc_hd__inv_2 _2441_ (.A(\device.uartRx.delayCounter[12] ),
    .Y(_1348_));
 sky130_fd_sc_hd__inv_2 _2442_ (.A(\device.uartRx.delayCounter[11] ),
    .Y(_1349_));
 sky130_fd_sc_hd__inv_2 _2443_ (.A(\device.uartRx.delayCounter[10] ),
    .Y(_1350_));
 sky130_fd_sc_hd__inv_2 _2444_ (.A(\device.uartRx.delayCounter[9] ),
    .Y(_1351_));
 sky130_fd_sc_hd__inv_2 _2445_ (.A(\device.uartRx.delayCounter[8] ),
    .Y(_1352_));
 sky130_fd_sc_hd__inv_2 _2446_ (.A(\device.uartRx.delayCounter[7] ),
    .Y(_1353_));
 sky130_fd_sc_hd__inv_2 _2447_ (.A(\device.uartRx.delayCounter[6] ),
    .Y(_1354_));
 sky130_fd_sc_hd__inv_2 _2448_ (.A(\device.uartRx.delayCounter[5] ),
    .Y(_1355_));
 sky130_fd_sc_hd__inv_2 _2449_ (.A(\device.uartRx.delayCounter[4] ),
    .Y(_1356_));
 sky130_fd_sc_hd__inv_2 _2450_ (.A(\device.uartRx.delayCounter[3] ),
    .Y(_1357_));
 sky130_fd_sc_hd__inv_2 _2451_ (.A(\device.uartRx.delayCounter[2] ),
    .Y(_1358_));
 sky130_fd_sc_hd__inv_2 _2452_ (.A(\device.uartRx.delayCounter[1] ),
    .Y(_1359_));
 sky130_fd_sc_hd__inv_2 _2453_ (.A(\device.uartRx.delayCounter[0] ),
    .Y(_1360_));
 sky130_fd_sc_hd__inv_2 _2454_ (.A(\device.uartTx.bitCounter[1] ),
    .Y(_1361_));
 sky130_fd_sc_hd__inv_2 _2455_ (.A(\device.uartTx.delayCounter[11] ),
    .Y(_1362_));
 sky130_fd_sc_hd__inv_2 _2456_ (.A(\device.uartTx.delayCounter[9] ),
    .Y(_1363_));
 sky130_fd_sc_hd__inv_2 _2457_ (.A(\device.uartTx.state[1] ),
    .Y(_1364_));
 sky130_fd_sc_hd__clkinv_2 _2458_ (.A(net511),
    .Y(_1365_));
 sky130_fd_sc_hd__inv_2 _2459_ (.A(\device.rxBuffer.endPointer[0] ),
    .Y(_1366_));
 sky130_fd_sc_hd__clkinv_2 _2460_ (.A(net514),
    .Y(_1367_));
 sky130_fd_sc_hd__inv_2 _2461_ (.A(\device.txBuffer.endPointer[3] ),
    .Y(_1368_));
 sky130_fd_sc_hd__inv_2 _2462_ (.A(\device.txBuffer.endPointer[0] ),
    .Y(_1369_));
 sky130_fd_sc_hd__inv_2 _2463_ (.A(\device.txBuffer.startPointer[3] ),
    .Y(_1370_));
 sky130_fd_sc_hd__inv_2 _2464_ (.A(net530),
    .Y(_1371_));
 sky130_fd_sc_hd__inv_4 _2465_ (.A(net630),
    .Y(_1372_));
 sky130_fd_sc_hd__inv_2 _2466_ (.A(net638),
    .Y(_1373_));
 sky130_fd_sc_hd__inv_4 _2467_ (.A(net3998),
    .Y(_1374_));
 sky130_fd_sc_hd__inv_2 _2468_ (.A(net628),
    .Y(_1375_));
 sky130_fd_sc_hd__clkinv_4 _2469_ (.A(\device.txBuffer.oe_buffered ),
    .Y(_1376_));
 sky130_fd_sc_hd__inv_2 _2470_ (.A(\device.rxBuffer.oe_buffered ),
    .Y(_1377_));
 sky130_fd_sc_hd__inv_2 _2471__1 (.A(clknet_leaf_35_wb_clk_i),
    .Y(net732));
 sky130_fd_sc_hd__or3b_4 _2472_ (.A(net529),
    .B(_1368_),
    .C_N(\device.txBuffer.endPointer[4] ),
    .X(_1378_));
 sky130_fd_sc_hd__xor2_1 _2473_ (.A(\device.txBuffer.endPointer[1] ),
    .B(net536),
    .X(_1379_));
 sky130_fd_sc_hd__or2_1 _2474_ (.A(_1369_),
    .B(net542),
    .X(_1380_));
 sky130_fd_sc_hd__nand2_1 _2475_ (.A(_1369_),
    .B(net542),
    .Y(_1381_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(_1381_),
    .A1(_1380_),
    .S(_1379_),
    .X(_1382_));
 sky130_fd_sc_hd__xnor2_2 _2477_ (.A(\device.txBuffer.endPointer[4] ),
    .B(\device.txBuffer.startPointer[4] ),
    .Y(_1383_));
 sky130_fd_sc_hd__nand2_4 _2478_ (.A(\device.txBuffer.endPointer[1] ),
    .B(\device.txBuffer.endPointer[0] ),
    .Y(_1384_));
 sky130_fd_sc_hd__and3_1 _2479_ (.A(\device.txBuffer.endPointer[2] ),
    .B(\device.txBuffer.endPointer[1] ),
    .C(\device.txBuffer.endPointer[0] ),
    .X(_1385_));
 sky130_fd_sc_hd__xor2_1 _2480_ (.A(\device.txBuffer.endPointer[3] ),
    .B(\device.txBuffer.startPointer[3] ),
    .X(_1386_));
 sky130_fd_sc_hd__o211a_1 _2481_ (.A1(\device.txBuffer.endPointer[3] ),
    .A2(_1370_),
    .B1(_1383_),
    .C1(_1385_),
    .X(_1387_));
 sky130_fd_sc_hd__xor2_2 _2482_ (.A(net529),
    .B(net531),
    .X(_1388_));
 sky130_fd_sc_hd__a31o_1 _2483_ (.A1(\device.txBuffer.endPointer[3] ),
    .A2(_1370_),
    .A3(_1385_),
    .B1(_1383_),
    .X(_1389_));
 sky130_fd_sc_hd__o21ai_1 _2484_ (.A1(_1384_),
    .A2(_1388_),
    .B1(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__a21oi_1 _2485_ (.A1(_1384_),
    .A2(_1388_),
    .B1(_1386_),
    .Y(_1391_));
 sky130_fd_sc_hd__nor2_1 _2486_ (.A(_1385_),
    .B(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__or4_4 _2487_ (.A(_1382_),
    .B(_1387_),
    .C(_1390_),
    .D(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__nand2_8 _2488_ (.A(\device.txBuffer.we_buffered ),
    .B(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__nor2_1 _2489_ (.A(_1369_),
    .B(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__and2_4 _2490_ (.A(_1372_),
    .B(net631),
    .X(_1396_));
 sky130_fd_sc_hd__nand2_4 _2491_ (.A(_1372_),
    .B(\wbPeripheralBusInterface.state[0] ),
    .Y(_1397_));
 sky130_fd_sc_hd__or4_2 _2492_ (.A(net145),
    .B(net144),
    .C(net148),
    .D(net147),
    .X(_1398_));
 sky130_fd_sc_hd__or3b_4 _2493_ (.A(net159),
    .B(net158),
    .C_N(net167),
    .X(_1399_));
 sky130_fd_sc_hd__or4bb_1 _2494_ (.A(net154),
    .B(net153),
    .C_N(net155),
    .D_N(net156),
    .X(_1400_));
 sky130_fd_sc_hd__or4_1 _2495_ (.A(net150),
    .B(net149),
    .C(net152),
    .D(net151),
    .X(_1401_));
 sky130_fd_sc_hd__or3_4 _2496_ (.A(_1399_),
    .B(_1400_),
    .C(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__nor4_4 _2497_ (.A(net143),
    .B(net142),
    .C(_1398_),
    .D(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__and2_4 _2498_ (.A(net638),
    .B(net502),
    .X(_1404_));
 sky130_fd_sc_hd__and3_4 _2499_ (.A(net193),
    .B(net509),
    .C(net484),
    .X(_1405_));
 sky130_fd_sc_hd__nor2_2 _2500_ (.A(net630),
    .B(net631),
    .Y(_1406_));
 sky130_fd_sc_hd__or2_2 _2501_ (.A(net630),
    .B(net631),
    .X(_1407_));
 sky130_fd_sc_hd__nand2_4 _2502_ (.A(net628),
    .B(net559),
    .Y(_1408_));
 sky130_fd_sc_hd__or4_2 _2503_ (.A(\wbPeripheralBusInterface.currentAddress[6] ),
    .B(\wbPeripheralBusInterface.currentAddress[7] ),
    .C(\wbPeripheralBusInterface.currentAddress[8] ),
    .D(\wbPeripheralBusInterface.currentAddress[9] ),
    .X(_1409_));
 sky130_fd_sc_hd__or3_4 _2504_ (.A(\wbPeripheralBusInterface.currentAddress[4] ),
    .B(\wbPeripheralBusInterface.currentAddress[5] ),
    .C(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__or4_4 _2505_ (.A(\wbPeripheralBusInterface.currentAddress[16] ),
    .B(\wbPeripheralBusInterface.currentAddress[17] ),
    .C(\wbPeripheralBusInterface.currentAddress[18] ),
    .D(\wbPeripheralBusInterface.currentAddress[19] ),
    .X(_1411_));
 sky130_fd_sc_hd__or4_4 _2506_ (.A(\wbPeripheralBusInterface.currentAddress[20] ),
    .B(\wbPeripheralBusInterface.currentAddress[21] ),
    .C(\wbPeripheralBusInterface.currentAddress[22] ),
    .D(\wbPeripheralBusInterface.currentAddress[23] ),
    .X(_1412_));
 sky130_fd_sc_hd__or4b_4 _2507_ (.A(\wbPeripheralBusInterface.currentAddress[13] ),
    .B(\wbPeripheralBusInterface.currentAddress[14] ),
    .C(\wbPeripheralBusInterface.currentAddress[15] ),
    .D_N(\wbPeripheralBusInterface.currentAddress[12] ),
    .X(_1413_));
 sky130_fd_sc_hd__or4_2 _2508_ (.A(_1406_),
    .B(_1411_),
    .C(_1412_),
    .D(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__or4b_1 _2509_ (.A(\wbPeripheralBusInterface.currentAddress[10] ),
    .B(\wbPeripheralBusInterface.currentAddress[11] ),
    .C(_1406_),
    .D_N(\wbPeripheralBusInterface.currentAddress[2] ),
    .X(_1415_));
 sky130_fd_sc_hd__or3_4 _2510_ (.A(\wbPeripheralBusInterface.currentAddress[3] ),
    .B(_1414_),
    .C(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__nor3_2 _2511_ (.A(_1408_),
    .B(_1410_),
    .C(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__or4_1 _2512_ (.A(_1406_),
    .B(_1411_),
    .C(_1412_),
    .D(_1413_),
    .X(_1418_));
 sky130_fd_sc_hd__a21oi_4 _2513_ (.A1(_1405_),
    .A2(_1417_),
    .B1(net642),
    .Y(_1419_));
 sky130_fd_sc_hd__or4b_4 _2514_ (.A(\device.txBuffer.endPointer[1] ),
    .B(_1369_),
    .C(_1394_),
    .D_N(net442),
    .X(_1420_));
 sky130_fd_sc_hd__or2_4 _2515_ (.A(_1378_),
    .B(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(net563),
    .A1(\device.txBuffer.buffer[25][7] ),
    .S(_1421_),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(net567),
    .A1(\device.txBuffer.buffer[25][6] ),
    .S(_1421_),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(net570),
    .A1(\device.txBuffer.buffer[25][5] ),
    .S(_1421_),
    .X(_0919_));
 sky130_fd_sc_hd__mux2_1 _2519_ (.A0(net574),
    .A1(\device.txBuffer.buffer[25][4] ),
    .S(_1421_),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(net577),
    .A1(\device.txBuffer.buffer[25][3] ),
    .S(_1421_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _2521_ (.A0(net581),
    .A1(\device.txBuffer.buffer[25][2] ),
    .S(_1421_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(net585),
    .A1(\device.txBuffer.buffer[25][1] ),
    .S(_1421_),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(net589),
    .A1(\device.txBuffer.buffer[25][0] ),
    .S(_1421_),
    .X(_0914_));
 sky130_fd_sc_hd__or3_4 _2524_ (.A(\device.txBuffer.endPointer[4] ),
    .B(_1368_),
    .C(net529),
    .X(_1422_));
 sky130_fd_sc_hd__or2_4 _2525_ (.A(_1420_),
    .B(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(net560),
    .A1(\device.txBuffer.buffer[9][7] ),
    .S(_1423_),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(net564),
    .A1(\device.txBuffer.buffer[9][6] ),
    .S(_1423_),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _2528_ (.A0(net568),
    .A1(\device.txBuffer.buffer[9][5] ),
    .S(_1423_),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _2529_ (.A0(net572),
    .A1(\device.txBuffer.buffer[9][4] ),
    .S(_1423_),
    .X(_0910_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(net576),
    .A1(\device.txBuffer.buffer[9][3] ),
    .S(_1423_),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(net580),
    .A1(\device.txBuffer.buffer[9][2] ),
    .S(_1423_),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(\device.txBuffer.dataIn_buffered[1] ),
    .A1(\device.txBuffer.buffer[9][1] ),
    .S(_1423_),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _2533_ (.A0(net588),
    .A1(\device.txBuffer.buffer[9][0] ),
    .S(_1423_),
    .X(_0906_));
 sky130_fd_sc_hd__or4b_4 _2534_ (.A(\device.txBuffer.endPointer[1] ),
    .B(\device.txBuffer.endPointer[0] ),
    .C(_1394_),
    .D_N(net442),
    .X(_1424_));
 sky130_fd_sc_hd__or2_4 _2535_ (.A(_1378_),
    .B(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(net563),
    .A1(\device.txBuffer.buffer[24][7] ),
    .S(_1425_),
    .X(_0905_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(net567),
    .A1(\device.txBuffer.buffer[24][6] ),
    .S(_1425_),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(net570),
    .A1(\device.txBuffer.buffer[24][5] ),
    .S(_1425_),
    .X(_0903_));
 sky130_fd_sc_hd__mux2_1 _2539_ (.A0(net574),
    .A1(\device.txBuffer.buffer[24][4] ),
    .S(_1425_),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(net577),
    .A1(\device.txBuffer.buffer[24][3] ),
    .S(_1425_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _2541_ (.A0(net582),
    .A1(\device.txBuffer.buffer[24][2] ),
    .S(_1425_),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(net585),
    .A1(\device.txBuffer.buffer[24][1] ),
    .S(_1425_),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _2543_ (.A0(net589),
    .A1(\device.txBuffer.buffer[24][0] ),
    .S(_1425_),
    .X(_0898_));
 sky130_fd_sc_hd__or3b_4 _2544_ (.A(\device.txBuffer.endPointer[4] ),
    .B(_1368_),
    .C_N(\device.txBuffer.endPointer[2] ),
    .X(_1426_));
 sky130_fd_sc_hd__nor2_8 _2545_ (.A(_1384_),
    .B(_1394_),
    .Y(_1427_));
 sky130_fd_sc_hd__nand2_8 _2546_ (.A(net442),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__nor2_8 _2547_ (.A(_1426_),
    .B(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(\device.txBuffer.buffer[15][7] ),
    .A1(net561),
    .S(_1429_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _2549_ (.A0(\device.txBuffer.buffer[15][6] ),
    .A1(net564),
    .S(_1429_),
    .X(_0859_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(\device.txBuffer.buffer[15][5] ),
    .A1(net568),
    .S(_1429_),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(\device.txBuffer.buffer[15][4] ),
    .A1(\device.txBuffer.dataIn_buffered[4] ),
    .S(_1429_),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(\device.txBuffer.buffer[15][3] ),
    .A1(net576),
    .S(_1429_),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_1 _2553_ (.A0(\device.txBuffer.buffer[15][2] ),
    .A1(net580),
    .S(_1429_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(\device.txBuffer.buffer[15][1] ),
    .A1(net584),
    .S(_1429_),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(\device.txBuffer.buffer[15][0] ),
    .A1(net588),
    .S(_1429_),
    .X(_0853_));
 sky130_fd_sc_hd__or3b_4 _2556_ (.A(\device.txBuffer.endPointer[3] ),
    .B(net529),
    .C_N(\device.txBuffer.endPointer[4] ),
    .X(_1430_));
 sky130_fd_sc_hd__or2_4 _2557_ (.A(_1424_),
    .B(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_1 _2558_ (.A0(net562),
    .A1(\device.txBuffer.buffer[16][7] ),
    .S(_1431_),
    .X(_0852_));
 sky130_fd_sc_hd__mux2_1 _2559_ (.A0(net566),
    .A1(\device.txBuffer.buffer[16][6] ),
    .S(_1431_),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(net569),
    .A1(\device.txBuffer.buffer[16][5] ),
    .S(_1431_),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(net573),
    .A1(\device.txBuffer.buffer[16][4] ),
    .S(_1431_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(net577),
    .A1(\device.txBuffer.buffer[16][3] ),
    .S(_1431_),
    .X(_0848_));
 sky130_fd_sc_hd__mux2_1 _2563_ (.A0(net581),
    .A1(\device.txBuffer.buffer[16][2] ),
    .S(_1431_),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_1 _2564_ (.A0(net586),
    .A1(\device.txBuffer.buffer[16][1] ),
    .S(_1431_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(net589),
    .A1(\device.txBuffer.buffer[16][0] ),
    .S(_1431_),
    .X(_0845_));
 sky130_fd_sc_hd__or2_4 _2566_ (.A(_1420_),
    .B(_1430_),
    .X(_1432_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(net562),
    .A1(\device.txBuffer.buffer[17][7] ),
    .S(_1432_),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_1 _2568_ (.A0(net566),
    .A1(\device.txBuffer.buffer[17][6] ),
    .S(_1432_),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(net569),
    .A1(\device.txBuffer.buffer[17][5] ),
    .S(_1432_),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(net573),
    .A1(\device.txBuffer.buffer[17][4] ),
    .S(_1432_),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _2571_ (.A0(net577),
    .A1(\device.txBuffer.buffer[17][3] ),
    .S(_1432_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(net581),
    .A1(\device.txBuffer.buffer[17][2] ),
    .S(_1432_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(net586),
    .A1(\device.txBuffer.buffer[17][1] ),
    .S(_1432_),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(net589),
    .A1(\device.txBuffer.buffer[17][0] ),
    .S(_1432_),
    .X(_0837_));
 sky130_fd_sc_hd__or4bb_4 _2575_ (.A(\device.txBuffer.endPointer[0] ),
    .B(_1394_),
    .C_N(net442),
    .D_N(\device.txBuffer.endPointer[1] ),
    .X(_1433_));
 sky130_fd_sc_hd__or2_4 _2576_ (.A(_1430_),
    .B(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__mux2_4 _2577_ (.A0(net562),
    .A1(\device.txBuffer.buffer[18][7] ),
    .S(_1434_),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_4 _2578_ (.A0(net566),
    .A1(\device.txBuffer.buffer[18][6] ),
    .S(_1434_),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _2579_ (.A0(net569),
    .A1(\device.txBuffer.buffer[18][5] ),
    .S(_1434_),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(net573),
    .A1(\device.txBuffer.buffer[18][4] ),
    .S(_1434_),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _2581_ (.A0(net577),
    .A1(\device.txBuffer.buffer[18][3] ),
    .S(_1434_),
    .X(_0832_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(net581),
    .A1(\device.txBuffer.buffer[18][2] ),
    .S(_1434_),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_4 _2583_ (.A0(net586),
    .A1(\device.txBuffer.buffer[18][1] ),
    .S(_1434_),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_4 _2584_ (.A0(net590),
    .A1(\device.txBuffer.buffer[18][0] ),
    .S(_1434_),
    .X(_0829_));
 sky130_fd_sc_hd__or3_4 _2585_ (.A(\device.txBuffer.endPointer[4] ),
    .B(\device.txBuffer.endPointer[3] ),
    .C(net529),
    .X(_1435_));
 sky130_fd_sc_hd__or2_4 _2586_ (.A(_1420_),
    .B(_1435_),
    .X(_1436_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(net560),
    .A1(\device.txBuffer.buffer[1][7] ),
    .S(_1436_),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _2588_ (.A0(net564),
    .A1(\device.txBuffer.buffer[1][6] ),
    .S(_1436_),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_1 _2589_ (.A0(net568),
    .A1(\device.txBuffer.buffer[1][5] ),
    .S(_1436_),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _2590_ (.A0(net572),
    .A1(\device.txBuffer.buffer[1][4] ),
    .S(_1436_),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_1 _2591_ (.A0(net576),
    .A1(\device.txBuffer.buffer[1][3] ),
    .S(_1436_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _2592_ (.A0(\device.txBuffer.dataIn_buffered[2] ),
    .A1(\device.txBuffer.buffer[1][2] ),
    .S(_1436_),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _2593_ (.A0(net584),
    .A1(\device.txBuffer.buffer[1][1] ),
    .S(_1436_),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _2594_ (.A0(net588),
    .A1(\device.txBuffer.buffer[1][0] ),
    .S(_1436_),
    .X(_0821_));
 sky130_fd_sc_hd__nand3_4 _2595_ (.A(\device.txBuffer.endPointer[4] ),
    .B(_1368_),
    .C(net529),
    .Y(_1437_));
 sky130_fd_sc_hd__or2_4 _2596_ (.A(_1424_),
    .B(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(net562),
    .A1(\device.txBuffer.buffer[20][7] ),
    .S(_1438_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _2598_ (.A0(net566),
    .A1(\device.txBuffer.buffer[20][6] ),
    .S(_1438_),
    .X(_0819_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(net569),
    .A1(\device.txBuffer.buffer[20][5] ),
    .S(_1438_),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(net573),
    .A1(\device.txBuffer.buffer[20][4] ),
    .S(_1438_),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_1 _2601_ (.A0(net578),
    .A1(\device.txBuffer.buffer[20][3] ),
    .S(_1438_),
    .X(_0816_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(net581),
    .A1(\device.txBuffer.buffer[20][2] ),
    .S(_1438_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _2603_ (.A0(net585),
    .A1(\device.txBuffer.buffer[20][1] ),
    .S(_1438_),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _2604_ (.A0(net591),
    .A1(\device.txBuffer.buffer[20][0] ),
    .S(_1438_),
    .X(_0813_));
 sky130_fd_sc_hd__or2_4 _2605_ (.A(_1420_),
    .B(_1437_),
    .X(_1439_));
 sky130_fd_sc_hd__mux2_1 _2606_ (.A0(net562),
    .A1(\device.txBuffer.buffer[21][7] ),
    .S(_1439_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(net566),
    .A1(\device.txBuffer.buffer[21][6] ),
    .S(_1439_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _2608_ (.A0(net569),
    .A1(\device.txBuffer.buffer[21][5] ),
    .S(_1439_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(net573),
    .A1(\device.txBuffer.buffer[21][4] ),
    .S(_1439_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _2610_ (.A0(net578),
    .A1(\device.txBuffer.buffer[21][3] ),
    .S(_1439_),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(net581),
    .A1(\device.txBuffer.buffer[21][2] ),
    .S(_1439_),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _2612_ (.A0(net585),
    .A1(\device.txBuffer.buffer[21][1] ),
    .S(_1439_),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(net591),
    .A1(\device.txBuffer.buffer[21][0] ),
    .S(_1439_),
    .X(_0805_));
 sky130_fd_sc_hd__nand3_4 _2614_ (.A(\device.rxBuffer.endPointer[4] ),
    .B(_1365_),
    .C(net512),
    .Y(_1440_));
 sky130_fd_sc_hd__nor4_4 _2615_ (.A(_1397_),
    .B(_1408_),
    .C(_1410_),
    .D(_1416_),
    .Y(_1441_));
 sky130_fd_sc_hd__a31oi_4 _2616_ (.A1(net190),
    .A2(net486),
    .A3(_1441_),
    .B1(net645),
    .Y(_1442_));
 sky130_fd_sc_hd__xor2_2 _2617_ (.A(\device.rxBuffer.endPointer[1] ),
    .B(net517),
    .X(_1443_));
 sky130_fd_sc_hd__or2_1 _2618_ (.A(_1366_),
    .B(net521),
    .X(_1444_));
 sky130_fd_sc_hd__xor2_4 _2619_ (.A(net512),
    .B(net513),
    .X(_1445_));
 sky130_fd_sc_hd__inv_2 _2620_ (.A(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__a21o_1 _2621_ (.A1(\device.rxBuffer.endPointer[1] ),
    .A2(_1446_),
    .B1(_1444_),
    .X(_1447_));
 sky130_fd_sc_hd__xnor2_2 _2622_ (.A(\device.rxBuffer.endPointer[4] ),
    .B(\device.rxBuffer.startPointer[4] ),
    .Y(_1448_));
 sky130_fd_sc_hd__nand2_2 _2623_ (.A(\device.rxBuffer.endPointer[1] ),
    .B(\device.rxBuffer.endPointer[0] ),
    .Y(_1449_));
 sky130_fd_sc_hd__nand3_2 _2624_ (.A(net512),
    .B(\device.rxBuffer.endPointer[1] ),
    .C(\device.rxBuffer.endPointer[0] ),
    .Y(_1450_));
 sky130_fd_sc_hd__or3_1 _2625_ (.A(_1365_),
    .B(\device.rxBuffer.startPointer[3] ),
    .C(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__a21oi_1 _2626_ (.A1(_1365_),
    .A2(\device.rxBuffer.startPointer[3] ),
    .B1(_1450_),
    .Y(_1452_));
 sky130_fd_sc_hd__mux2_1 _2627_ (.A0(_1451_),
    .A1(_1452_),
    .S(_1448_),
    .X(_1453_));
 sky130_fd_sc_hd__xor2_1 _2628_ (.A(net511),
    .B(\device.rxBuffer.startPointer[3] ),
    .X(_1454_));
 sky130_fd_sc_hd__a21oi_1 _2629_ (.A1(_1366_),
    .A2(net521),
    .B1(_1443_),
    .Y(_1455_));
 sky130_fd_sc_hd__a221o_1 _2630_ (.A1(_1445_),
    .A2(_1449_),
    .B1(_1450_),
    .B2(_1454_),
    .C1(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__a211o_4 _2631_ (.A1(_1443_),
    .A2(_1447_),
    .B1(_1453_),
    .C1(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__and2_1 _2632_ (.A(\device.rxBuffer.we_buffered ),
    .B(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__nand2_4 _2633_ (.A(\device.rxBuffer.we_buffered ),
    .B(_1457_),
    .Y(_1459_));
 sky130_fd_sc_hd__nand2_1 _2634_ (.A(net438),
    .B(_1458_),
    .Y(_1460_));
 sky130_fd_sc_hd__or3_4 _2635_ (.A(\device.rxBuffer.endPointer[1] ),
    .B(\device.rxBuffer.endPointer[0] ),
    .C(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__nor2_8 _2636_ (.A(_1440_),
    .B(net405),
    .Y(_1462_));
 sky130_fd_sc_hd__mux2_1 _2637_ (.A0(\device.rxBuffer.buffer[20][7] ),
    .A1(net594),
    .S(_1462_),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _2638_ (.A0(\device.rxBuffer.buffer[20][6] ),
    .A1(net599),
    .S(_1462_),
    .X(_0803_));
 sky130_fd_sc_hd__mux2_1 _2639_ (.A0(\device.rxBuffer.buffer[20][5] ),
    .A1(net604),
    .S(_1462_),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _2640_ (.A0(\device.rxBuffer.buffer[20][4] ),
    .A1(net606),
    .S(_1462_),
    .X(_0801_));
 sky130_fd_sc_hd__mux2_1 _2641_ (.A0(\device.rxBuffer.buffer[20][3] ),
    .A1(net612),
    .S(_1462_),
    .X(_0800_));
 sky130_fd_sc_hd__mux2_1 _2642_ (.A0(\device.rxBuffer.buffer[20][2] ),
    .A1(net616),
    .S(_1462_),
    .X(_0799_));
 sky130_fd_sc_hd__mux2_1 _2643_ (.A0(\device.rxBuffer.buffer[20][1] ),
    .A1(net620),
    .S(_1462_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _2644_ (.A0(\device.rxBuffer.buffer[20][0] ),
    .A1(net624),
    .S(_1462_),
    .X(_0797_));
 sky130_fd_sc_hd__nor2_8 _2645_ (.A(_1433_),
    .B(_1437_),
    .Y(_1463_));
 sky130_fd_sc_hd__mux2_1 _2646_ (.A0(\device.txBuffer.buffer[22][7] ),
    .A1(net562),
    .S(_1463_),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _2647_ (.A0(\device.txBuffer.buffer[22][6] ),
    .A1(net566),
    .S(_1463_),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _2648_ (.A0(\device.txBuffer.buffer[22][5] ),
    .A1(net569),
    .S(_1463_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _2649_ (.A0(\device.txBuffer.buffer[22][4] ),
    .A1(net573),
    .S(_1463_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _2650_ (.A0(\device.txBuffer.buffer[22][3] ),
    .A1(net577),
    .S(_1463_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _2651_ (.A0(\device.txBuffer.buffer[22][2] ),
    .A1(net581),
    .S(_1463_),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _2652_ (.A0(\device.txBuffer.buffer[22][1] ),
    .A1(net585),
    .S(_1463_),
    .X(_0790_));
 sky130_fd_sc_hd__mux2_1 _2653_ (.A0(\device.txBuffer.buffer[22][0] ),
    .A1(net590),
    .S(_1463_),
    .X(_0789_));
 sky130_fd_sc_hd__or3_4 _2654_ (.A(\device.rxBuffer.endPointer[1] ),
    .B(_1366_),
    .C(_1460_),
    .X(_1464_));
 sky130_fd_sc_hd__or2_4 _2655_ (.A(_1440_),
    .B(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__mux2_1 _2656_ (.A0(net594),
    .A1(\device.rxBuffer.buffer[21][7] ),
    .S(_1465_),
    .X(_0788_));
 sky130_fd_sc_hd__mux2_1 _2657_ (.A0(net599),
    .A1(\device.rxBuffer.buffer[21][6] ),
    .S(_1465_),
    .X(_0787_));
 sky130_fd_sc_hd__mux2_1 _2658_ (.A0(net604),
    .A1(\device.rxBuffer.buffer[21][5] ),
    .S(_1465_),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(net607),
    .A1(\device.rxBuffer.buffer[21][4] ),
    .S(_1465_),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _2660_ (.A0(net612),
    .A1(\device.rxBuffer.buffer[21][3] ),
    .S(_1465_),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(net616),
    .A1(\device.rxBuffer.buffer[21][2] ),
    .S(_1465_),
    .X(_0783_));
 sky130_fd_sc_hd__mux2_1 _2662_ (.A0(net620),
    .A1(\device.rxBuffer.buffer[21][1] ),
    .S(_1465_),
    .X(_0782_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(net624),
    .A1(\device.rxBuffer.buffer[21][0] ),
    .S(_1465_),
    .X(_0781_));
 sky130_fd_sc_hd__nor2_8 _2664_ (.A(_1428_),
    .B(_1437_),
    .Y(_1466_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(\device.txBuffer.buffer[23][7] ),
    .A1(net562),
    .S(_1466_),
    .X(_0780_));
 sky130_fd_sc_hd__mux2_1 _2666_ (.A0(\device.txBuffer.buffer[23][6] ),
    .A1(net566),
    .S(_1466_),
    .X(_0779_));
 sky130_fd_sc_hd__mux2_1 _2667_ (.A0(\device.txBuffer.buffer[23][5] ),
    .A1(net570),
    .S(_1466_),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_1 _2668_ (.A0(\device.txBuffer.buffer[23][4] ),
    .A1(net573),
    .S(_1466_),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _2669_ (.A0(\device.txBuffer.buffer[23][3] ),
    .A1(net577),
    .S(_1466_),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_1 _2670_ (.A0(\device.txBuffer.buffer[23][2] ),
    .A1(net581),
    .S(_1466_),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _2671_ (.A0(\device.txBuffer.buffer[23][1] ),
    .A1(net585),
    .S(_1466_),
    .X(_0774_));
 sky130_fd_sc_hd__mux2_1 _2672_ (.A0(\device.txBuffer.buffer[23][0] ),
    .A1(net590),
    .S(_1466_),
    .X(_0773_));
 sky130_fd_sc_hd__or3b_4 _2673_ (.A(\device.rxBuffer.endPointer[0] ),
    .B(_1460_),
    .C_N(\device.rxBuffer.endPointer[1] ),
    .X(_1467_));
 sky130_fd_sc_hd__or2_4 _2674_ (.A(_1440_),
    .B(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_1 _2675_ (.A0(net594),
    .A1(\device.rxBuffer.buffer[22][7] ),
    .S(_1468_),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _2676_ (.A0(net599),
    .A1(\device.rxBuffer.buffer[22][6] ),
    .S(_1468_),
    .X(_0771_));
 sky130_fd_sc_hd__mux2_1 _2677_ (.A0(net604),
    .A1(\device.rxBuffer.buffer[22][5] ),
    .S(_1468_),
    .X(_0770_));
 sky130_fd_sc_hd__mux2_1 _2678_ (.A0(net607),
    .A1(\device.rxBuffer.buffer[22][4] ),
    .S(_1468_),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_1 _2679_ (.A0(net613),
    .A1(\device.rxBuffer.buffer[22][3] ),
    .S(_1468_),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_1 _2680_ (.A0(net617),
    .A1(\device.rxBuffer.buffer[22][2] ),
    .S(_1468_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _2681_ (.A0(net621),
    .A1(\device.rxBuffer.buffer[22][1] ),
    .S(_1468_),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _2682_ (.A0(net623),
    .A1(\device.rxBuffer.buffer[22][0] ),
    .S(_1468_),
    .X(_0765_));
 sky130_fd_sc_hd__or3b_4 _2683_ (.A(net511),
    .B(net512),
    .C_N(\device.rxBuffer.endPointer[4] ),
    .X(_1469_));
 sky130_fd_sc_hd__or2_4 _2684_ (.A(_1467_),
    .B(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_1 _2685_ (.A0(net594),
    .A1(\device.rxBuffer.buffer[18][7] ),
    .S(_1470_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _2686_ (.A0(net599),
    .A1(\device.rxBuffer.buffer[18][6] ),
    .S(_1470_),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _2687_ (.A0(net604),
    .A1(\device.rxBuffer.buffer[18][5] ),
    .S(_1470_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _2688_ (.A0(net607),
    .A1(\device.rxBuffer.buffer[18][4] ),
    .S(_1470_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _2689_ (.A0(net612),
    .A1(\device.rxBuffer.buffer[18][3] ),
    .S(_1470_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _2690_ (.A0(net616),
    .A1(\device.rxBuffer.buffer[18][2] ),
    .S(_1470_),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _2691_ (.A0(net620),
    .A1(\device.rxBuffer.buffer[18][1] ),
    .S(_1470_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _2692_ (.A0(net622),
    .A1(\device.rxBuffer.buffer[18][0] ),
    .S(_1470_),
    .X(_0729_));
 sky130_fd_sc_hd__nand3_4 _2693_ (.A(\device.txBuffer.endPointer[4] ),
    .B(\device.txBuffer.endPointer[3] ),
    .C(net529),
    .Y(_1471_));
 sky130_fd_sc_hd__nor2_8 _2694_ (.A(_1428_),
    .B(_1471_),
    .Y(_1472_));
 sky130_fd_sc_hd__mux2_1 _2695_ (.A0(\device.txBuffer.buffer[31][7] ),
    .A1(net563),
    .S(_1472_),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(\device.txBuffer.buffer[31][6] ),
    .A1(net566),
    .S(_1472_),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _2697_ (.A0(\device.txBuffer.buffer[31][5] ),
    .A1(net571),
    .S(_1472_),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _2698_ (.A0(\device.txBuffer.buffer[31][4] ),
    .A1(net574),
    .S(_1472_),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _2699_ (.A0(\device.txBuffer.buffer[31][3] ),
    .A1(net579),
    .S(_1472_),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _2700_ (.A0(\device.txBuffer.buffer[31][2] ),
    .A1(net582),
    .S(_1472_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _2701_ (.A0(\device.txBuffer.buffer[31][1] ),
    .A1(net585),
    .S(_1472_),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _2702_ (.A0(\device.txBuffer.buffer[31][0] ),
    .A1(net589),
    .S(_1472_),
    .X(_0719_));
 sky130_fd_sc_hd__or2_4 _2703_ (.A(_1428_),
    .B(_1435_),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_1 _2704_ (.A0(net560),
    .A1(\device.txBuffer.buffer[3][7] ),
    .S(_1473_),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _2705_ (.A0(net564),
    .A1(\device.txBuffer.buffer[3][6] ),
    .S(_1473_),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _2706_ (.A0(net568),
    .A1(\device.txBuffer.buffer[3][5] ),
    .S(_1473_),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _2707_ (.A0(net572),
    .A1(\device.txBuffer.buffer[3][4] ),
    .S(_1473_),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _2708_ (.A0(net576),
    .A1(\device.txBuffer.buffer[3][3] ),
    .S(_1473_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(net580),
    .A1(\device.txBuffer.buffer[3][2] ),
    .S(_1473_),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _2710_ (.A0(net584),
    .A1(\device.txBuffer.buffer[3][1] ),
    .S(_1473_),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _2711_ (.A0(net588),
    .A1(\device.txBuffer.buffer[3][0] ),
    .S(_1473_),
    .X(_0711_));
 sky130_fd_sc_hd__or3b_4 _2712_ (.A(\device.txBuffer.endPointer[4] ),
    .B(\device.txBuffer.endPointer[3] ),
    .C_N(net529),
    .X(_1474_));
 sky130_fd_sc_hd__or2_4 _2713_ (.A(_1424_),
    .B(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__mux2_1 _2714_ (.A0(net560),
    .A1(\device.txBuffer.buffer[4][7] ),
    .S(_1475_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _2715_ (.A0(net565),
    .A1(\device.txBuffer.buffer[4][6] ),
    .S(_1475_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _2716_ (.A0(net569),
    .A1(\device.txBuffer.buffer[4][5] ),
    .S(_1475_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _2717_ (.A0(net575),
    .A1(\device.txBuffer.buffer[4][4] ),
    .S(_1475_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _2718_ (.A0(net578),
    .A1(\device.txBuffer.buffer[4][3] ),
    .S(_1475_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _2719_ (.A0(net583),
    .A1(\device.txBuffer.buffer[4][2] ),
    .S(_1475_),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _2720_ (.A0(net587),
    .A1(\device.txBuffer.buffer[4][1] ),
    .S(_1475_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(net591),
    .A1(\device.txBuffer.buffer[4][0] ),
    .S(_1475_),
    .X(_0703_));
 sky130_fd_sc_hd__or2_4 _2722_ (.A(_1420_),
    .B(_1474_),
    .X(_1476_));
 sky130_fd_sc_hd__mux2_1 _2723_ (.A0(net562),
    .A1(\device.txBuffer.buffer[5][7] ),
    .S(_1476_),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _2724_ (.A0(net565),
    .A1(\device.txBuffer.buffer[5][6] ),
    .S(_1476_),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _2725_ (.A0(net569),
    .A1(\device.txBuffer.buffer[5][5] ),
    .S(_1476_),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _2726_ (.A0(net575),
    .A1(\device.txBuffer.buffer[5][4] ),
    .S(_1476_),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _2727_ (.A0(net578),
    .A1(\device.txBuffer.buffer[5][3] ),
    .S(_1476_),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _2728_ (.A0(net583),
    .A1(\device.txBuffer.buffer[5][2] ),
    .S(_1476_),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _2729_ (.A0(net587),
    .A1(\device.txBuffer.buffer[5][1] ),
    .S(_1476_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _2730_ (.A0(net591),
    .A1(\device.txBuffer.buffer[5][0] ),
    .S(_1476_),
    .X(_0695_));
 sky130_fd_sc_hd__or2_4 _2731_ (.A(_1433_),
    .B(_1474_),
    .X(_1477_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(net562),
    .A1(\device.txBuffer.buffer[6][7] ),
    .S(_1477_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _2733_ (.A0(net565),
    .A1(\device.txBuffer.buffer[6][6] ),
    .S(_1477_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(net569),
    .A1(\device.txBuffer.buffer[6][5] ),
    .S(_1477_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(net575),
    .A1(\device.txBuffer.buffer[6][4] ),
    .S(_1477_),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _2736_ (.A0(net578),
    .A1(\device.txBuffer.buffer[6][3] ),
    .S(_1477_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _2737_ (.A0(net583),
    .A1(\device.txBuffer.buffer[6][2] ),
    .S(_1477_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(net587),
    .A1(\device.txBuffer.buffer[6][1] ),
    .S(_1477_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _2739_ (.A0(net591),
    .A1(\device.txBuffer.buffer[6][0] ),
    .S(_1477_),
    .X(_0687_));
 sky130_fd_sc_hd__or2_4 _2740_ (.A(_1428_),
    .B(_1474_),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _2741_ (.A0(net561),
    .A1(\device.txBuffer.buffer[7][7] ),
    .S(_1478_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _2742_ (.A0(net565),
    .A1(\device.txBuffer.buffer[7][6] ),
    .S(_1478_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _2743_ (.A0(net569),
    .A1(\device.txBuffer.buffer[7][5] ),
    .S(_1478_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _2744_ (.A0(net575),
    .A1(\device.txBuffer.buffer[7][4] ),
    .S(_1478_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _2745_ (.A0(net578),
    .A1(\device.txBuffer.buffer[7][3] ),
    .S(_1478_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _2746_ (.A0(net583),
    .A1(\device.txBuffer.buffer[7][2] ),
    .S(_1478_),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(net587),
    .A1(\device.txBuffer.buffer[7][1] ),
    .S(_1478_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(net591),
    .A1(\device.txBuffer.buffer[7][0] ),
    .S(_1478_),
    .X(_0679_));
 sky130_fd_sc_hd__or2_4 _2749_ (.A(_1422_),
    .B(_1424_),
    .X(_1479_));
 sky130_fd_sc_hd__mux2_1 _2750_ (.A0(net560),
    .A1(\device.txBuffer.buffer[8][7] ),
    .S(_1479_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(net564),
    .A1(\device.txBuffer.buffer[8][6] ),
    .S(_1479_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _2752_ (.A0(net568),
    .A1(\device.txBuffer.buffer[8][5] ),
    .S(_1479_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _2753_ (.A0(net572),
    .A1(\device.txBuffer.buffer[8][4] ),
    .S(_1479_),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _2754_ (.A0(net579),
    .A1(\device.txBuffer.buffer[8][3] ),
    .S(_1479_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _2755_ (.A0(net580),
    .A1(\device.txBuffer.buffer[8][2] ),
    .S(_1479_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _2756_ (.A0(net584),
    .A1(\device.txBuffer.buffer[8][1] ),
    .S(_1479_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(net588),
    .A1(\device.txBuffer.buffer[8][0] ),
    .S(_1479_),
    .X(_0671_));
 sky130_fd_sc_hd__or2_4 _2758_ (.A(_1424_),
    .B(_1435_),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_1 _2759_ (.A0(net560),
    .A1(\device.txBuffer.buffer[0][7] ),
    .S(_1480_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _2760_ (.A0(net564),
    .A1(\device.txBuffer.buffer[0][6] ),
    .S(_1480_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _2761_ (.A0(net568),
    .A1(\device.txBuffer.buffer[0][5] ),
    .S(_1480_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _2762_ (.A0(net572),
    .A1(\device.txBuffer.buffer[0][4] ),
    .S(_1480_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(net576),
    .A1(\device.txBuffer.buffer[0][3] ),
    .S(_1480_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _2764_ (.A0(\device.txBuffer.dataIn_buffered[2] ),
    .A1(\device.txBuffer.buffer[0][2] ),
    .S(_1480_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _2765_ (.A0(net584),
    .A1(\device.txBuffer.buffer[0][1] ),
    .S(_1480_),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _2766_ (.A0(net588),
    .A1(\device.txBuffer.buffer[0][0] ),
    .S(_1480_),
    .X(_0663_));
 sky130_fd_sc_hd__or2_4 _2767_ (.A(_1422_),
    .B(_1433_),
    .X(_1481_));
 sky130_fd_sc_hd__mux2_1 _2768_ (.A0(net560),
    .A1(\device.txBuffer.buffer[10][7] ),
    .S(_1481_),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _2769_ (.A0(net565),
    .A1(\device.txBuffer.buffer[10][6] ),
    .S(_1481_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _2770_ (.A0(net571),
    .A1(\device.txBuffer.buffer[10][5] ),
    .S(_1481_),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _2771_ (.A0(net572),
    .A1(\device.txBuffer.buffer[10][4] ),
    .S(_1481_),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _2772_ (.A0(net576),
    .A1(\device.txBuffer.buffer[10][3] ),
    .S(_1481_),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _2773_ (.A0(net580),
    .A1(\device.txBuffer.buffer[10][2] ),
    .S(_1481_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _2774_ (.A0(net584),
    .A1(\device.txBuffer.buffer[10][1] ),
    .S(_1481_),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(net588),
    .A1(\device.txBuffer.buffer[10][0] ),
    .S(_1481_),
    .X(_0655_));
 sky130_fd_sc_hd__nor2_1 _2776_ (.A(_1366_),
    .B(_1459_),
    .Y(_1482_));
 sky130_fd_sc_hd__nor2_4 _2777_ (.A(_1449_),
    .B(_1459_),
    .Y(_1483_));
 sky130_fd_sc_hd__nand2_8 _2778_ (.A(net438),
    .B(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__nor2_8 _2779_ (.A(_1440_),
    .B(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__mux2_1 _2780_ (.A0(\device.rxBuffer.buffer[23][7] ),
    .A1(net594),
    .S(_1485_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _2781_ (.A0(\device.rxBuffer.buffer[23][6] ),
    .A1(net599),
    .S(_1485_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _2782_ (.A0(\device.rxBuffer.buffer[23][5] ),
    .A1(net604),
    .S(_1485_),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _2783_ (.A0(\device.rxBuffer.buffer[23][4] ),
    .A1(net607),
    .S(_1485_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _2784_ (.A0(\device.rxBuffer.buffer[23][3] ),
    .A1(net613),
    .S(_1485_),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _2785_ (.A0(\device.rxBuffer.buffer[23][2] ),
    .A1(net617),
    .S(_1485_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _2786_ (.A0(\device.rxBuffer.buffer[23][1] ),
    .A1(net621),
    .S(_1485_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _2787_ (.A0(\device.rxBuffer.buffer[23][0] ),
    .A1(net624),
    .S(_1485_),
    .X(_0647_));
 sky130_fd_sc_hd__or2_4 _2788_ (.A(_1422_),
    .B(_1428_),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_1 _2789_ (.A0(net561),
    .A1(\device.txBuffer.buffer[11][7] ),
    .S(_1486_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _2790_ (.A0(net565),
    .A1(\device.txBuffer.buffer[11][6] ),
    .S(_1486_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _2791_ (.A0(net571),
    .A1(\device.txBuffer.buffer[11][5] ),
    .S(_1486_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _2792_ (.A0(net572),
    .A1(\device.txBuffer.buffer[11][4] ),
    .S(_1486_),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _2793_ (.A0(net576),
    .A1(\device.txBuffer.buffer[11][3] ),
    .S(_1486_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _2794_ (.A0(net580),
    .A1(\device.txBuffer.buffer[11][2] ),
    .S(_1486_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _2795_ (.A0(net584),
    .A1(\device.txBuffer.buffer[11][1] ),
    .S(_1486_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(net588),
    .A1(\device.txBuffer.buffer[11][0] ),
    .S(_1486_),
    .X(_0639_));
 sky130_fd_sc_hd__nand3b_4 _2797_ (.A_N(\device.rxBuffer.endPointer[2] ),
    .B(net511),
    .C(\device.rxBuffer.endPointer[4] ),
    .Y(_1487_));
 sky130_fd_sc_hd__nor2_8 _2798_ (.A(_1461_),
    .B(_1487_),
    .Y(_1488_));
 sky130_fd_sc_hd__mux2_1 _2799_ (.A0(\device.rxBuffer.buffer[24][7] ),
    .A1(net595),
    .S(_1488_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _2800_ (.A0(\device.rxBuffer.buffer[24][6] ),
    .A1(net600),
    .S(_1488_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _2801_ (.A0(\device.rxBuffer.buffer[24][5] ),
    .A1(net604),
    .S(_1488_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(\device.rxBuffer.buffer[24][4] ),
    .A1(net609),
    .S(_1488_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _2803_ (.A0(\device.rxBuffer.buffer[24][3] ),
    .A1(net613),
    .S(_1488_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _2804_ (.A0(\device.rxBuffer.buffer[24][2] ),
    .A1(net617),
    .S(_1488_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _2805_ (.A0(\device.rxBuffer.buffer[24][1] ),
    .A1(net621),
    .S(_1488_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _2806_ (.A0(\device.rxBuffer.buffer[24][0] ),
    .A1(net625),
    .S(_1488_),
    .X(_0631_));
 sky130_fd_sc_hd__or2_4 _2807_ (.A(_1464_),
    .B(_1487_),
    .X(_1489_));
 sky130_fd_sc_hd__mux2_1 _2808_ (.A0(net595),
    .A1(\device.rxBuffer.buffer[25][7] ),
    .S(_1489_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _2809_ (.A0(net600),
    .A1(\device.rxBuffer.buffer[25][6] ),
    .S(_1489_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _2810_ (.A0(net604),
    .A1(\device.rxBuffer.buffer[25][5] ),
    .S(_1489_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _2811_ (.A0(net609),
    .A1(\device.rxBuffer.buffer[25][4] ),
    .S(_1489_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _2812_ (.A0(net613),
    .A1(\device.rxBuffer.buffer[25][3] ),
    .S(_1489_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _2813_ (.A0(net617),
    .A1(\device.rxBuffer.buffer[25][2] ),
    .S(_1489_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _2814_ (.A0(net621),
    .A1(\device.rxBuffer.buffer[25][1] ),
    .S(_1489_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _2815_ (.A0(net625),
    .A1(\device.rxBuffer.buffer[25][0] ),
    .S(_1489_),
    .X(_0623_));
 sky130_fd_sc_hd__or2_4 _2816_ (.A(_1424_),
    .B(_1426_),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _2817_ (.A0(net560),
    .A1(\device.txBuffer.buffer[12][7] ),
    .S(_1490_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _2818_ (.A0(net564),
    .A1(\device.txBuffer.buffer[12][6] ),
    .S(_1490_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _2819_ (.A0(net568),
    .A1(\device.txBuffer.buffer[12][5] ),
    .S(_1490_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _2820_ (.A0(net572),
    .A1(\device.txBuffer.buffer[12][4] ),
    .S(_1490_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _2821_ (.A0(net576),
    .A1(\device.txBuffer.buffer[12][3] ),
    .S(_1490_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _2822_ (.A0(net580),
    .A1(\device.txBuffer.buffer[12][2] ),
    .S(_1490_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _2823_ (.A0(net584),
    .A1(\device.txBuffer.buffer[12][1] ),
    .S(_1490_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _2824_ (.A0(\device.txBuffer.dataIn_buffered[0] ),
    .A1(\device.txBuffer.buffer[12][0] ),
    .S(_1490_),
    .X(_0615_));
 sky130_fd_sc_hd__or2_4 _2825_ (.A(_1420_),
    .B(_1426_),
    .X(_1491_));
 sky130_fd_sc_hd__mux2_1 _2826_ (.A0(net560),
    .A1(\device.txBuffer.buffer[13][7] ),
    .S(_1491_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _2827_ (.A0(net564),
    .A1(\device.txBuffer.buffer[13][6] ),
    .S(_1491_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _2828_ (.A0(net568),
    .A1(\device.txBuffer.buffer[13][5] ),
    .S(_1491_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _2829_ (.A0(net572),
    .A1(\device.txBuffer.buffer[13][4] ),
    .S(_1491_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _2830_ (.A0(net576),
    .A1(\device.txBuffer.buffer[13][3] ),
    .S(_1491_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _2831_ (.A0(net580),
    .A1(\device.txBuffer.buffer[13][2] ),
    .S(_1491_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _2832_ (.A0(\device.txBuffer.dataIn_buffered[1] ),
    .A1(\device.txBuffer.buffer[13][1] ),
    .S(_1491_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _2833_ (.A0(\device.txBuffer.dataIn_buffered[0] ),
    .A1(\device.txBuffer.buffer[13][0] ),
    .S(_1491_),
    .X(_0607_));
 sky130_fd_sc_hd__or2_4 _2834_ (.A(_1467_),
    .B(_1487_),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(net595),
    .A1(\device.rxBuffer.buffer[26][7] ),
    .S(_1492_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _2836_ (.A0(net600),
    .A1(\device.rxBuffer.buffer[26][6] ),
    .S(_1492_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _2837_ (.A0(net605),
    .A1(\device.rxBuffer.buffer[26][5] ),
    .S(_1492_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _2838_ (.A0(net609),
    .A1(\device.rxBuffer.buffer[26][4] ),
    .S(_1492_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _2839_ (.A0(net613),
    .A1(\device.rxBuffer.buffer[26][3] ),
    .S(_1492_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _2840_ (.A0(net617),
    .A1(\device.rxBuffer.buffer[26][2] ),
    .S(_1492_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _2841_ (.A0(net621),
    .A1(\device.rxBuffer.buffer[26][1] ),
    .S(_1492_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _2842_ (.A0(net625),
    .A1(\device.rxBuffer.buffer[26][0] ),
    .S(_1492_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_8 _2843_ (.A(_1484_),
    .B(_1487_),
    .Y(_1493_));
 sky130_fd_sc_hd__mux2_1 _2844_ (.A0(\device.rxBuffer.buffer[27][7] ),
    .A1(net595),
    .S(_1493_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _2845_ (.A0(\device.rxBuffer.buffer[27][6] ),
    .A1(net600),
    .S(_1493_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(\device.rxBuffer.buffer[27][5] ),
    .A1(net605),
    .S(_1493_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _2847_ (.A0(\device.rxBuffer.buffer[27][4] ),
    .A1(\device.rxBuffer.dataIn_buffered[4] ),
    .S(_1493_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _2848_ (.A0(\device.rxBuffer.buffer[27][3] ),
    .A1(net613),
    .S(_1493_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(\device.rxBuffer.buffer[27][2] ),
    .A1(net617),
    .S(_1493_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _2850_ (.A0(\device.rxBuffer.buffer[27][1] ),
    .A1(net621),
    .S(_1493_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(\device.rxBuffer.buffer[27][0] ),
    .A1(net625),
    .S(_1493_),
    .X(_0591_));
 sky130_fd_sc_hd__nor2_8 _2852_ (.A(_1426_),
    .B(_1433_),
    .Y(_1494_));
 sky130_fd_sc_hd__mux2_1 _2853_ (.A0(\device.txBuffer.buffer[14][7] ),
    .A1(net561),
    .S(_1494_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _2854_ (.A0(\device.txBuffer.buffer[14][6] ),
    .A1(net564),
    .S(_1494_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _2855_ (.A0(\device.txBuffer.buffer[14][5] ),
    .A1(net568),
    .S(_1494_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _2856_ (.A0(\device.txBuffer.buffer[14][4] ),
    .A1(\device.txBuffer.dataIn_buffered[4] ),
    .S(_1494_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _2857_ (.A0(\device.txBuffer.buffer[14][3] ),
    .A1(net579),
    .S(_1494_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _2858_ (.A0(\device.txBuffer.buffer[14][2] ),
    .A1(net580),
    .S(_1494_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _2859_ (.A0(\device.txBuffer.buffer[14][1] ),
    .A1(net584),
    .S(_1494_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _2860_ (.A0(\device.txBuffer.buffer[14][0] ),
    .A1(net588),
    .S(_1494_),
    .X(_0583_));
 sky130_fd_sc_hd__nor2_1 _2861_ (.A(_1445_),
    .B(_1454_),
    .Y(_1495_));
 sky130_fd_sc_hd__and4_4 _2862_ (.A(_1444_),
    .B(_1448_),
    .C(_1455_),
    .D(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__nor2_1 _2863_ (.A(_1377_),
    .B(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__nand2_2 _2864_ (.A(net517),
    .B(net522),
    .Y(_1498_));
 sky130_fd_sc_hd__or2_1 _2865_ (.A(net517),
    .B(net522),
    .X(_1499_));
 sky130_fd_sc_hd__nand2_1 _2866_ (.A(_1498_),
    .B(net499),
    .Y(_1500_));
 sky130_fd_sc_hd__and3_4 _2867_ (.A(net513),
    .B(net517),
    .C(net521),
    .X(_1501_));
 sky130_fd_sc_hd__a21oi_2 _2868_ (.A1(net518),
    .A2(net525),
    .B1(\device.rxBuffer.startPointer[2] ),
    .Y(_1502_));
 sky130_fd_sc_hd__nor2_1 _2869_ (.A(_1501_),
    .B(net497),
    .Y(_1503_));
 sky130_fd_sc_hd__or2_1 _2870_ (.A(_1501_),
    .B(net497),
    .X(_1504_));
 sky130_fd_sc_hd__mux4_2 _2871_ (.A0(\device.rxBuffer.buffer[5][7] ),
    .A1(\device.rxBuffer.buffer[6][7] ),
    .A2(\device.rxBuffer.buffer[7][7] ),
    .A3(\device.rxBuffer.buffer[4][7] ),
    .S0(net523),
    .S1(net515),
    .X(_1505_));
 sky130_fd_sc_hd__and2_4 _2872_ (.A(\device.rxBuffer.startPointer[3] ),
    .B(_1501_),
    .X(_1506_));
 sky130_fd_sc_hd__nor2_1 _2873_ (.A(\device.rxBuffer.startPointer[3] ),
    .B(_1501_),
    .Y(_1507_));
 sky130_fd_sc_hd__nor2_2 _2874_ (.A(_1506_),
    .B(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__or2_4 _2875_ (.A(_1506_),
    .B(_1507_),
    .X(_1509_));
 sky130_fd_sc_hd__mux4_1 _2876_ (.A0(\device.rxBuffer.buffer[1][7] ),
    .A1(\device.rxBuffer.buffer[3][7] ),
    .A2(\device.rxBuffer.buffer[2][7] ),
    .A3(\device.rxBuffer.buffer[0][7] ),
    .S0(net515),
    .S1(net520),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_1 _2877_ (.A0(_1505_),
    .A1(_1510_),
    .S(net473),
    .X(_1511_));
 sky130_fd_sc_hd__mux4_2 _2878_ (.A0(\device.rxBuffer.buffer[13][7] ),
    .A1(\device.rxBuffer.buffer[14][7] ),
    .A2(\device.rxBuffer.buffer[15][7] ),
    .A3(\device.rxBuffer.buffer[12][7] ),
    .S0(net523),
    .S1(net516),
    .X(_1512_));
 sky130_fd_sc_hd__mux4_2 _2879_ (.A0(\device.rxBuffer.buffer[9][7] ),
    .A1(\device.rxBuffer.buffer[11][7] ),
    .A2(\device.rxBuffer.buffer[10][7] ),
    .A3(\device.rxBuffer.buffer[8][7] ),
    .S0(net515),
    .S1(net520),
    .X(_1513_));
 sky130_fd_sc_hd__a21o_1 _2880_ (.A1(net473),
    .A2(_1513_),
    .B1(net454),
    .X(_1514_));
 sky130_fd_sc_hd__a21o_1 _2881_ (.A1(net476),
    .A2(_1512_),
    .B1(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__xnor2_4 _2882_ (.A(\device.rxBuffer.startPointer[4] ),
    .B(_1506_),
    .Y(_1516_));
 sky130_fd_sc_hd__xor2_4 _2883_ (.A(\device.rxBuffer.startPointer[4] ),
    .B(_1506_),
    .X(_1517_));
 sky130_fd_sc_hd__o211a_1 _2884_ (.A1(net456),
    .A2(_1511_),
    .B1(_1515_),
    .C1(_1516_),
    .X(_1518_));
 sky130_fd_sc_hd__mux4_2 _2885_ (.A0(\device.rxBuffer.buffer[21][7] ),
    .A1(\device.rxBuffer.buffer[22][7] ),
    .A2(\device.rxBuffer.buffer[23][7] ),
    .A3(\device.rxBuffer.buffer[20][7] ),
    .S0(net526),
    .S1(net518),
    .X(_1519_));
 sky130_fd_sc_hd__mux4_1 _2886_ (.A0(\device.rxBuffer.buffer[17][7] ),
    .A1(\device.rxBuffer.buffer[19][7] ),
    .A2(\device.rxBuffer.buffer[18][7] ),
    .A3(\device.rxBuffer.buffer[16][7] ),
    .S0(net518),
    .S1(net526),
    .X(_1520_));
 sky130_fd_sc_hd__a21o_1 _2887_ (.A1(net478),
    .A2(_1519_),
    .B1(net456),
    .X(_1521_));
 sky130_fd_sc_hd__a21o_1 _2888_ (.A1(net474),
    .A2(_1520_),
    .B1(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__mux4_2 _2889_ (.A0(\device.rxBuffer.buffer[29][7] ),
    .A1(\device.rxBuffer.buffer[31][7] ),
    .A2(\device.rxBuffer.buffer[30][7] ),
    .A3(\device.rxBuffer.buffer[28][7] ),
    .S0(net519),
    .S1(net525),
    .X(_1523_));
 sky130_fd_sc_hd__mux4_1 _2890_ (.A0(\device.rxBuffer.buffer[25][7] ),
    .A1(\device.rxBuffer.buffer[26][7] ),
    .A2(\device.rxBuffer.buffer[27][7] ),
    .A3(\device.rxBuffer.buffer[24][7] ),
    .S0(net526),
    .S1(net519),
    .X(_1524_));
 sky130_fd_sc_hd__a21o_1 _2891_ (.A1(net474),
    .A2(_1524_),
    .B1(net454),
    .X(_1525_));
 sky130_fd_sc_hd__a21o_2 _2892_ (.A1(net478),
    .A2(_1523_),
    .B1(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__a31o_2 _2893_ (.A1(_1517_),
    .A2(_1522_),
    .A3(_1526_),
    .B1(_1518_),
    .X(_1527_));
 sky130_fd_sc_hd__and2_4 _2894_ (.A(\device.rxBuffer.we_buffered ),
    .B(_1496_),
    .X(_1528_));
 sky130_fd_sc_hd__nand2_4 _2895_ (.A(\device.rxBuffer.we_buffered ),
    .B(_1496_),
    .Y(_1529_));
 sky130_fd_sc_hd__a221o_1 _2896_ (.A1(_1377_),
    .A2(\device.rxBuffer.dataOut[7] ),
    .B1(net435),
    .B2(_1527_),
    .C1(_1528_),
    .X(_1530_));
 sky130_fd_sc_hd__o211a_1 _2897_ (.A1(net596),
    .A2(_1529_),
    .B1(_1530_),
    .C1(net437),
    .X(_0580_));
 sky130_fd_sc_hd__mux4_1 _2898_ (.A0(\device.rxBuffer.buffer[1][6] ),
    .A1(\device.rxBuffer.buffer[3][6] ),
    .A2(\device.rxBuffer.buffer[2][6] ),
    .A3(\device.rxBuffer.buffer[0][6] ),
    .S0(net515),
    .S1(net520),
    .X(_1531_));
 sky130_fd_sc_hd__mux4_1 _2899_ (.A0(\device.rxBuffer.buffer[5][6] ),
    .A1(\device.rxBuffer.buffer[6][6] ),
    .A2(\device.rxBuffer.buffer[7][6] ),
    .A3(\device.rxBuffer.buffer[4][6] ),
    .S0(net523),
    .S1(net515),
    .X(_1532_));
 sky130_fd_sc_hd__mux2_1 _2900_ (.A0(_1531_),
    .A1(_1532_),
    .S(net476),
    .X(_1533_));
 sky130_fd_sc_hd__mux4_2 _2901_ (.A0(\device.rxBuffer.buffer[13][6] ),
    .A1(\device.rxBuffer.buffer[14][6] ),
    .A2(\device.rxBuffer.buffer[15][6] ),
    .A3(\device.rxBuffer.buffer[12][6] ),
    .S0(net523),
    .S1(net516),
    .X(_1534_));
 sky130_fd_sc_hd__mux4_2 _2902_ (.A0(\device.rxBuffer.buffer[9][6] ),
    .A1(\device.rxBuffer.buffer[11][6] ),
    .A2(\device.rxBuffer.buffer[10][6] ),
    .A3(\device.rxBuffer.buffer[8][6] ),
    .S0(net515),
    .S1(net520),
    .X(_1535_));
 sky130_fd_sc_hd__a21o_1 _2903_ (.A1(net473),
    .A2(_1535_),
    .B1(net454),
    .X(_1536_));
 sky130_fd_sc_hd__a21o_1 _2904_ (.A1(net476),
    .A2(_1534_),
    .B1(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__o211a_2 _2905_ (.A1(net456),
    .A2(_1533_),
    .B1(_1537_),
    .C1(_1516_),
    .X(_1538_));
 sky130_fd_sc_hd__mux4_2 _2906_ (.A0(\device.rxBuffer.buffer[21][6] ),
    .A1(\device.rxBuffer.buffer[22][6] ),
    .A2(\device.rxBuffer.buffer[23][6] ),
    .A3(\device.rxBuffer.buffer[20][6] ),
    .S0(net526),
    .S1(net518),
    .X(_1539_));
 sky130_fd_sc_hd__mux4_1 _2907_ (.A0(\device.rxBuffer.buffer[17][6] ),
    .A1(\device.rxBuffer.buffer[19][6] ),
    .A2(\device.rxBuffer.buffer[18][6] ),
    .A3(\device.rxBuffer.buffer[16][6] ),
    .S0(net518),
    .S1(net526),
    .X(_1540_));
 sky130_fd_sc_hd__a21o_1 _2908_ (.A1(net478),
    .A2(_1539_),
    .B1(net456),
    .X(_1541_));
 sky130_fd_sc_hd__a21o_1 _2909_ (.A1(net474),
    .A2(_1540_),
    .B1(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__mux4_1 _2910_ (.A0(\device.rxBuffer.buffer[29][6] ),
    .A1(\device.rxBuffer.buffer[31][6] ),
    .A2(\device.rxBuffer.buffer[30][6] ),
    .A3(\device.rxBuffer.buffer[28][6] ),
    .S0(net518),
    .S1(net525),
    .X(_1543_));
 sky130_fd_sc_hd__mux4_2 _2911_ (.A0(\device.rxBuffer.buffer[25][6] ),
    .A1(\device.rxBuffer.buffer[26][6] ),
    .A2(\device.rxBuffer.buffer[27][6] ),
    .A3(\device.rxBuffer.buffer[24][6] ),
    .S0(net527),
    .S1(net519),
    .X(_1544_));
 sky130_fd_sc_hd__a21o_1 _2912_ (.A1(net474),
    .A2(_1544_),
    .B1(net454),
    .X(_1545_));
 sky130_fd_sc_hd__a21o_2 _2913_ (.A1(net479),
    .A2(_1543_),
    .B1(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__a31o_2 _2914_ (.A1(_1517_),
    .A2(_1542_),
    .A3(_1546_),
    .B1(_1538_),
    .X(_1547_));
 sky130_fd_sc_hd__a221o_1 _2915_ (.A1(_1377_),
    .A2(\device.rxBuffer.dataOut[6] ),
    .B1(net435),
    .B2(_1547_),
    .C1(_1528_),
    .X(_1548_));
 sky130_fd_sc_hd__o211a_1 _2916_ (.A1(net601),
    .A2(_1529_),
    .B1(_1548_),
    .C1(net437),
    .X(_0579_));
 sky130_fd_sc_hd__mux4_2 _2917_ (.A0(\device.rxBuffer.buffer[1][5] ),
    .A1(\device.rxBuffer.buffer[3][5] ),
    .A2(\device.rxBuffer.buffer[2][5] ),
    .A3(\device.rxBuffer.buffer[0][5] ),
    .S0(net515),
    .S1(net521),
    .X(_1549_));
 sky130_fd_sc_hd__mux4_1 _2918_ (.A0(\device.rxBuffer.buffer[5][5] ),
    .A1(\device.rxBuffer.buffer[6][5] ),
    .A2(\device.rxBuffer.buffer[7][5] ),
    .A3(\device.rxBuffer.buffer[4][5] ),
    .S0(net523),
    .S1(net516),
    .X(_1550_));
 sky130_fd_sc_hd__nand2_1 _2919_ (.A(net436),
    .B(net454),
    .Y(_1551_));
 sky130_fd_sc_hd__mux4_2 _2920_ (.A0(\device.rxBuffer.buffer[21][5] ),
    .A1(\device.rxBuffer.buffer[22][5] ),
    .A2(\device.rxBuffer.buffer[23][5] ),
    .A3(\device.rxBuffer.buffer[20][5] ),
    .S0(net526),
    .S1(net518),
    .X(_1552_));
 sky130_fd_sc_hd__mux4_1 _2921_ (.A0(\device.rxBuffer.buffer[17][5] ),
    .A1(\device.rxBuffer.buffer[19][5] ),
    .A2(\device.rxBuffer.buffer[18][5] ),
    .A3(\device.rxBuffer.buffer[16][5] ),
    .S0(net518),
    .S1(net526),
    .X(_1553_));
 sky130_fd_sc_hd__mux4_2 _2922_ (.A0(\device.rxBuffer.buffer[13][5] ),
    .A1(\device.rxBuffer.buffer[14][5] ),
    .A2(\device.rxBuffer.buffer[15][5] ),
    .A3(\device.rxBuffer.buffer[12][5] ),
    .S0(net523),
    .S1(net516),
    .X(_1554_));
 sky130_fd_sc_hd__mux4_2 _2923_ (.A0(\device.rxBuffer.buffer[9][5] ),
    .A1(\device.rxBuffer.buffer[11][5] ),
    .A2(\device.rxBuffer.buffer[10][5] ),
    .A3(\device.rxBuffer.buffer[8][5] ),
    .S0(net515),
    .S1(net520),
    .X(_1555_));
 sky130_fd_sc_hd__and2_1 _2924_ (.A(net473),
    .B(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__mux4_2 _2925_ (.A0(\device.rxBuffer.buffer[29][5] ),
    .A1(\device.rxBuffer.buffer[31][5] ),
    .A2(\device.rxBuffer.buffer[30][5] ),
    .A3(\device.rxBuffer.buffer[28][5] ),
    .S0(net518),
    .S1(net525),
    .X(_1557_));
 sky130_fd_sc_hd__mux4_1 _2926_ (.A0(\device.rxBuffer.buffer[25][5] ),
    .A1(\device.rxBuffer.buffer[26][5] ),
    .A2(\device.rxBuffer.buffer[27][5] ),
    .A3(\device.rxBuffer.buffer[24][5] ),
    .S0(net527),
    .S1(net519),
    .X(_1558_));
 sky130_fd_sc_hd__a21o_1 _2927_ (.A1(net476),
    .A2(_1554_),
    .B1(net454),
    .X(_1559_));
 sky130_fd_sc_hd__mux2_1 _2928_ (.A0(_1549_),
    .A1(_1550_),
    .S(net476),
    .X(_1560_));
 sky130_fd_sc_hd__o221a_2 _2929_ (.A1(_1556_),
    .A2(_1559_),
    .B1(_1560_),
    .B2(net456),
    .C1(_1516_),
    .X(_1561_));
 sky130_fd_sc_hd__a21o_1 _2930_ (.A1(net478),
    .A2(_1552_),
    .B1(net457),
    .X(_1562_));
 sky130_fd_sc_hd__a21o_1 _2931_ (.A1(net474),
    .A2(_1553_),
    .B1(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__a21o_1 _2932_ (.A1(net479),
    .A2(_1557_),
    .B1(net455),
    .X(_1564_));
 sky130_fd_sc_hd__a21o_2 _2933_ (.A1(net474),
    .A2(_1558_),
    .B1(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__a31o_2 _2934_ (.A1(_1517_),
    .A2(_1563_),
    .A3(_1565_),
    .B1(_1561_),
    .X(_1566_));
 sky130_fd_sc_hd__a221o_1 _2935_ (.A1(_1377_),
    .A2(\device.rxBuffer.dataOut[5] ),
    .B1(net435),
    .B2(_1566_),
    .C1(_1528_),
    .X(_1567_));
 sky130_fd_sc_hd__o211a_1 _2936_ (.A1(net602),
    .A2(_1529_),
    .B1(_1567_),
    .C1(net437),
    .X(_0578_));
 sky130_fd_sc_hd__mux4_1 _2937_ (.A0(\device.rxBuffer.buffer[1][4] ),
    .A1(\device.rxBuffer.buffer[3][4] ),
    .A2(\device.rxBuffer.buffer[2][4] ),
    .A3(\device.rxBuffer.buffer[0][4] ),
    .S0(net515),
    .S1(net521),
    .X(_1568_));
 sky130_fd_sc_hd__mux4_2 _2938_ (.A0(\device.rxBuffer.buffer[5][4] ),
    .A1(\device.rxBuffer.buffer[6][4] ),
    .A2(\device.rxBuffer.buffer[7][4] ),
    .A3(\device.rxBuffer.buffer[4][4] ),
    .S0(net523),
    .S1(net516),
    .X(_1569_));
 sky130_fd_sc_hd__mux4_2 _2939_ (.A0(\device.rxBuffer.buffer[21][4] ),
    .A1(\device.rxBuffer.buffer[22][4] ),
    .A2(\device.rxBuffer.buffer[23][4] ),
    .A3(\device.rxBuffer.buffer[20][4] ),
    .S0(net522),
    .S1(net517),
    .X(_1570_));
 sky130_fd_sc_hd__mux4_1 _2940_ (.A0(\device.rxBuffer.buffer[17][4] ),
    .A1(\device.rxBuffer.buffer[19][4] ),
    .A2(\device.rxBuffer.buffer[18][4] ),
    .A3(\device.rxBuffer.buffer[16][4] ),
    .S0(net517),
    .S1(net522),
    .X(_1571_));
 sky130_fd_sc_hd__mux4_1 _2941_ (.A0(\device.rxBuffer.buffer[29][4] ),
    .A1(\device.rxBuffer.buffer[31][4] ),
    .A2(\device.rxBuffer.buffer[30][4] ),
    .A3(\device.rxBuffer.buffer[28][4] ),
    .S0(net518),
    .S1(net525),
    .X(_1572_));
 sky130_fd_sc_hd__mux4_2 _2942_ (.A0(\device.rxBuffer.buffer[25][4] ),
    .A1(\device.rxBuffer.buffer[26][4] ),
    .A2(\device.rxBuffer.buffer[27][4] ),
    .A3(\device.rxBuffer.buffer[24][4] ),
    .S0(net527),
    .S1(net519),
    .X(_1573_));
 sky130_fd_sc_hd__mux4_2 _2943_ (.A0(\device.rxBuffer.buffer[13][4] ),
    .A1(\device.rxBuffer.buffer[14][4] ),
    .A2(\device.rxBuffer.buffer[15][4] ),
    .A3(\device.rxBuffer.buffer[12][4] ),
    .S0(net523),
    .S1(net516),
    .X(_1574_));
 sky130_fd_sc_hd__mux4_2 _2944_ (.A0(\device.rxBuffer.buffer[9][4] ),
    .A1(\device.rxBuffer.buffer[11][4] ),
    .A2(\device.rxBuffer.buffer[10][4] ),
    .A3(\device.rxBuffer.buffer[8][4] ),
    .S0(net515),
    .S1(net520),
    .X(_1575_));
 sky130_fd_sc_hd__and2_1 _2945_ (.A(net473),
    .B(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__a21o_1 _2946_ (.A1(net476),
    .A2(_1574_),
    .B1(net454),
    .X(_1577_));
 sky130_fd_sc_hd__mux2_1 _2947_ (.A0(_1568_),
    .A1(_1569_),
    .S(net476),
    .X(_1578_));
 sky130_fd_sc_hd__o221a_2 _2948_ (.A1(_1576_),
    .A2(_1577_),
    .B1(_1578_),
    .B2(net456),
    .C1(_1516_),
    .X(_1579_));
 sky130_fd_sc_hd__a21o_1 _2949_ (.A1(net477),
    .A2(_1570_),
    .B1(net457),
    .X(_1580_));
 sky130_fd_sc_hd__a21o_1 _2950_ (.A1(net473),
    .A2(_1571_),
    .B1(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__a21o_1 _2951_ (.A1(net479),
    .A2(_1572_),
    .B1(net455),
    .X(_1582_));
 sky130_fd_sc_hd__a21o_2 _2952_ (.A1(net474),
    .A2(_1573_),
    .B1(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__a31o_2 _2953_ (.A1(_1517_),
    .A2(_1581_),
    .A3(_1583_),
    .B1(_1579_),
    .X(_1584_));
 sky130_fd_sc_hd__a221o_1 _2954_ (.A1(_1377_),
    .A2(\device.rxBuffer.dataOut[4] ),
    .B1(net435),
    .B2(_1584_),
    .C1(_1528_),
    .X(_1585_));
 sky130_fd_sc_hd__o211a_1 _2955_ (.A1(net608),
    .A2(_1529_),
    .B1(_1585_),
    .C1(net437),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _2956_ (.A0(\device.rxBuffer.buffer[7][3] ),
    .A1(\device.rxBuffer.buffer[6][3] ),
    .S(net522),
    .X(_1586_));
 sky130_fd_sc_hd__o221a_1 _2957_ (.A1(net513),
    .A2(\device.rxBuffer.buffer[4][3] ),
    .B1(net498),
    .B2(\device.rxBuffer.buffer[5][3] ),
    .C1(net477),
    .X(_1587_));
 sky130_fd_sc_hd__o21a_1 _2958_ (.A1(net480),
    .A2(_1586_),
    .B1(_1587_),
    .X(_1588_));
 sky130_fd_sc_hd__mux2_1 _2959_ (.A0(\device.rxBuffer.buffer[3][3] ),
    .A1(\device.rxBuffer.buffer[2][3] ),
    .S(net524),
    .X(_1589_));
 sky130_fd_sc_hd__o22a_1 _2960_ (.A1(\device.rxBuffer.buffer[0][3] ),
    .A2(net497),
    .B1(_1589_),
    .B2(net480),
    .X(_1590_));
 sky130_fd_sc_hd__o211a_1 _2961_ (.A1(\device.rxBuffer.buffer[1][3] ),
    .A2(net498),
    .B1(net473),
    .C1(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_1 _2962_ (.A0(\device.rxBuffer.buffer[23][3] ),
    .A1(\device.rxBuffer.buffer[22][3] ),
    .S(net526),
    .X(_1592_));
 sky130_fd_sc_hd__o221a_1 _2963_ (.A1(\device.rxBuffer.buffer[20][3] ),
    .A2(net514),
    .B1(net500),
    .B2(\device.rxBuffer.buffer[21][3] ),
    .C1(net478),
    .X(_1593_));
 sky130_fd_sc_hd__o21a_1 _2964_ (.A1(net482),
    .A2(_1592_),
    .B1(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(\device.rxBuffer.buffer[19][3] ),
    .A1(\device.rxBuffer.buffer[18][3] ),
    .S(net525),
    .X(_1595_));
 sky130_fd_sc_hd__o22a_1 _2966_ (.A1(\device.rxBuffer.buffer[16][3] ),
    .A2(net497),
    .B1(_1595_),
    .B2(net482),
    .X(_1596_));
 sky130_fd_sc_hd__o211a_1 _2967_ (.A1(\device.rxBuffer.buffer[17][3] ),
    .A2(net500),
    .B1(net474),
    .C1(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__mux2_1 _2968_ (.A0(\device.rxBuffer.buffer[15][3] ),
    .A1(\device.rxBuffer.buffer[14][3] ),
    .S(net524),
    .X(_1598_));
 sky130_fd_sc_hd__o221a_1 _2969_ (.A1(net513),
    .A2(\device.rxBuffer.buffer[12][3] ),
    .B1(net498),
    .B2(\device.rxBuffer.buffer[13][3] ),
    .C1(net477),
    .X(_1599_));
 sky130_fd_sc_hd__o21a_1 _2970_ (.A1(net480),
    .A2(_1598_),
    .B1(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__a21o_1 _2971_ (.A1(\device.rxBuffer.buffer[8][3] ),
    .A2(_1501_),
    .B1(net497),
    .X(_1601_));
 sky130_fd_sc_hd__mux2_1 _2972_ (.A0(\device.rxBuffer.buffer[11][3] ),
    .A1(\device.rxBuffer.buffer[10][3] ),
    .S(net524),
    .X(_1602_));
 sky130_fd_sc_hd__o22a_1 _2973_ (.A1(\device.rxBuffer.buffer[9][3] ),
    .A2(net498),
    .B1(net480),
    .B2(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__mux2_1 _2974_ (.A0(\device.rxBuffer.buffer[27][3] ),
    .A1(\device.rxBuffer.buffer[26][3] ),
    .S(net527),
    .X(_1604_));
 sky130_fd_sc_hd__o22a_1 _2975_ (.A1(\device.rxBuffer.buffer[24][3] ),
    .A2(_1367_),
    .B1(net501),
    .B2(\device.rxBuffer.buffer[25][3] ),
    .X(_1605_));
 sky130_fd_sc_hd__o211a_1 _2976_ (.A1(net482),
    .A2(_1604_),
    .B1(_1605_),
    .C1(net475),
    .X(_1606_));
 sky130_fd_sc_hd__mux2_1 _2977_ (.A0(\device.rxBuffer.buffer[31][3] ),
    .A1(\device.rxBuffer.buffer[30][3] ),
    .S(net528),
    .X(_1607_));
 sky130_fd_sc_hd__or2_1 _2978_ (.A(net482),
    .B(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__o221a_1 _2979_ (.A1(net514),
    .A2(\device.rxBuffer.buffer[28][3] ),
    .B1(\device.rxBuffer.buffer[29][3] ),
    .B2(net500),
    .C1(net478),
    .X(_1609_));
 sky130_fd_sc_hd__a211o_1 _2980_ (.A1(_1601_),
    .A2(_1603_),
    .B1(net454),
    .C1(_1600_),
    .X(_1610_));
 sky130_fd_sc_hd__or3_1 _2981_ (.A(net456),
    .B(_1588_),
    .C(_1591_),
    .X(_1611_));
 sky130_fd_sc_hd__a211o_1 _2982_ (.A1(_1608_),
    .A2(_1609_),
    .B1(net455),
    .C1(_1606_),
    .X(_1612_));
 sky130_fd_sc_hd__o311a_2 _2983_ (.A1(net457),
    .A2(_1594_),
    .A3(_1597_),
    .B1(_1612_),
    .C1(_1517_),
    .X(_1613_));
 sky130_fd_sc_hd__a31o_1 _2984_ (.A1(_1516_),
    .A2(_1610_),
    .A3(_1611_),
    .B1(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__a221o_1 _2985_ (.A1(_1377_),
    .A2(\device.rxBuffer.dataOut[3] ),
    .B1(net435),
    .B2(_1614_),
    .C1(_1528_),
    .X(_1615_));
 sky130_fd_sc_hd__o211a_1 _2986_ (.A1(net610),
    .A2(_1529_),
    .B1(_1615_),
    .C1(net437),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(\device.rxBuffer.buffer[7][2] ),
    .A1(\device.rxBuffer.buffer[6][2] ),
    .S(net523),
    .X(_1616_));
 sky130_fd_sc_hd__o221a_1 _2988_ (.A1(net513),
    .A2(\device.rxBuffer.buffer[4][2] ),
    .B1(net498),
    .B2(\device.rxBuffer.buffer[5][2] ),
    .C1(net477),
    .X(_1617_));
 sky130_fd_sc_hd__o21a_1 _2989_ (.A1(net480),
    .A2(_1616_),
    .B1(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__mux2_1 _2990_ (.A0(\device.rxBuffer.buffer[3][2] ),
    .A1(\device.rxBuffer.buffer[2][2] ),
    .S(net520),
    .X(_1619_));
 sky130_fd_sc_hd__o22a_1 _2991_ (.A1(\device.rxBuffer.buffer[0][2] ),
    .A2(net497),
    .B1(_1619_),
    .B2(net480),
    .X(_1620_));
 sky130_fd_sc_hd__o211a_1 _2992_ (.A1(\device.rxBuffer.buffer[1][2] ),
    .A2(net498),
    .B1(net473),
    .C1(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__mux2_1 _2993_ (.A0(\device.rxBuffer.buffer[19][2] ),
    .A1(\device.rxBuffer.buffer[18][2] ),
    .S(net525),
    .X(_1622_));
 sky130_fd_sc_hd__o22a_1 _2994_ (.A1(\device.rxBuffer.buffer[16][2] ),
    .A2(net497),
    .B1(_1622_),
    .B2(net482),
    .X(_1623_));
 sky130_fd_sc_hd__o211a_1 _2995_ (.A1(\device.rxBuffer.buffer[17][2] ),
    .A2(net501),
    .B1(net474),
    .C1(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(\device.rxBuffer.buffer[23][2] ),
    .A1(\device.rxBuffer.buffer[22][2] ),
    .S(net526),
    .X(_1625_));
 sky130_fd_sc_hd__o221a_1 _2997_ (.A1(\device.rxBuffer.buffer[20][2] ),
    .A2(net514),
    .B1(net500),
    .B2(\device.rxBuffer.buffer[21][2] ),
    .C1(net478),
    .X(_1626_));
 sky130_fd_sc_hd__o21a_1 _2998_ (.A1(net482),
    .A2(_1625_),
    .B1(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__mux2_1 _2999_ (.A0(\device.rxBuffer.buffer[27][2] ),
    .A1(\device.rxBuffer.buffer[26][2] ),
    .S(net527),
    .X(_1628_));
 sky130_fd_sc_hd__o22a_1 _3000_ (.A1(\device.rxBuffer.buffer[24][2] ),
    .A2(_1367_),
    .B1(net501),
    .B2(\device.rxBuffer.buffer[25][2] ),
    .X(_1629_));
 sky130_fd_sc_hd__o211a_1 _3001_ (.A1(net483),
    .A2(_1628_),
    .B1(_1629_),
    .C1(net475),
    .X(_1630_));
 sky130_fd_sc_hd__mux2_1 _3002_ (.A0(\device.rxBuffer.buffer[31][2] ),
    .A1(\device.rxBuffer.buffer[30][2] ),
    .S(net528),
    .X(_1631_));
 sky130_fd_sc_hd__or2_1 _3003_ (.A(net482),
    .B(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__o221a_1 _3004_ (.A1(net514),
    .A2(\device.rxBuffer.buffer[28][2] ),
    .B1(\device.rxBuffer.buffer[29][2] ),
    .B2(net500),
    .C1(net479),
    .X(_1633_));
 sky130_fd_sc_hd__mux2_1 _3005_ (.A0(\device.rxBuffer.buffer[15][2] ),
    .A1(\device.rxBuffer.buffer[14][2] ),
    .S(net524),
    .X(_1634_));
 sky130_fd_sc_hd__o221a_1 _3006_ (.A1(net513),
    .A2(\device.rxBuffer.buffer[12][2] ),
    .B1(net499),
    .B2(\device.rxBuffer.buffer[13][2] ),
    .C1(net476),
    .X(_1635_));
 sky130_fd_sc_hd__o21a_1 _3007_ (.A1(net481),
    .A2(_1634_),
    .B1(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__a21o_1 _3008_ (.A1(\device.rxBuffer.buffer[8][2] ),
    .A2(_1501_),
    .B1(net497),
    .X(_1637_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(\device.rxBuffer.buffer[11][2] ),
    .A1(\device.rxBuffer.buffer[10][2] ),
    .S(net520),
    .X(_1638_));
 sky130_fd_sc_hd__o22a_1 _3010_ (.A1(\device.rxBuffer.buffer[9][2] ),
    .A2(net498),
    .B1(net480),
    .B2(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__a211o_1 _3011_ (.A1(_1637_),
    .A2(_1639_),
    .B1(net454),
    .C1(_1636_),
    .X(_1640_));
 sky130_fd_sc_hd__or3_1 _3012_ (.A(net456),
    .B(_1618_),
    .C(_1621_),
    .X(_1641_));
 sky130_fd_sc_hd__a211o_1 _3013_ (.A1(_1632_),
    .A2(_1633_),
    .B1(net455),
    .C1(_1630_),
    .X(_1642_));
 sky130_fd_sc_hd__o311a_2 _3014_ (.A1(net457),
    .A2(_1624_),
    .A3(_1627_),
    .B1(_1642_),
    .C1(_1517_),
    .X(_1643_));
 sky130_fd_sc_hd__a31o_1 _3015_ (.A1(_1516_),
    .A2(_1640_),
    .A3(_1641_),
    .B1(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__a221o_1 _3016_ (.A1(_1377_),
    .A2(\device.rxBuffer.dataOut[2] ),
    .B1(net435),
    .B2(_1644_),
    .C1(_1528_),
    .X(_1645_));
 sky130_fd_sc_hd__o211a_1 _3017_ (.A1(net614),
    .A2(_1529_),
    .B1(_1645_),
    .C1(net437),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(\device.rxBuffer.buffer[7][1] ),
    .A1(\device.rxBuffer.buffer[6][1] ),
    .S(net522),
    .X(_1646_));
 sky130_fd_sc_hd__o221a_1 _3019_ (.A1(net513),
    .A2(\device.rxBuffer.buffer[4][1] ),
    .B1(net498),
    .B2(\device.rxBuffer.buffer[5][1] ),
    .C1(net476),
    .X(_1647_));
 sky130_fd_sc_hd__o21a_1 _3020_ (.A1(net480),
    .A2(_1646_),
    .B1(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__mux2_1 _3021_ (.A0(\device.rxBuffer.buffer[3][1] ),
    .A1(\device.rxBuffer.buffer[2][1] ),
    .S(net520),
    .X(_1649_));
 sky130_fd_sc_hd__o22a_1 _3022_ (.A1(\device.rxBuffer.buffer[0][1] ),
    .A2(net497),
    .B1(_1649_),
    .B2(net480),
    .X(_1650_));
 sky130_fd_sc_hd__o211a_1 _3023_ (.A1(\device.rxBuffer.buffer[1][1] ),
    .A2(net498),
    .B1(net473),
    .C1(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(\device.rxBuffer.buffer[23][1] ),
    .A1(\device.rxBuffer.buffer[22][1] ),
    .S(net526),
    .X(_1652_));
 sky130_fd_sc_hd__o221a_1 _3025_ (.A1(\device.rxBuffer.buffer[20][1] ),
    .A2(\device.rxBuffer.startPointer[2] ),
    .B1(net500),
    .B2(\device.rxBuffer.buffer[21][1] ),
    .C1(net478),
    .X(_1653_));
 sky130_fd_sc_hd__o21a_1 _3026_ (.A1(net482),
    .A2(_1652_),
    .B1(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__mux2_1 _3027_ (.A0(\device.rxBuffer.buffer[19][1] ),
    .A1(\device.rxBuffer.buffer[18][1] ),
    .S(net525),
    .X(_1655_));
 sky130_fd_sc_hd__o22a_1 _3028_ (.A1(\device.rxBuffer.buffer[16][1] ),
    .A2(_1502_),
    .B1(_1655_),
    .B2(net482),
    .X(_1656_));
 sky130_fd_sc_hd__o211a_1 _3029_ (.A1(\device.rxBuffer.buffer[17][1] ),
    .A2(net500),
    .B1(net474),
    .C1(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__mux2_1 _3030_ (.A0(\device.rxBuffer.buffer[27][1] ),
    .A1(\device.rxBuffer.buffer[26][1] ),
    .S(net527),
    .X(_1658_));
 sky130_fd_sc_hd__o22a_1 _3031_ (.A1(\device.rxBuffer.buffer[24][1] ),
    .A2(_1367_),
    .B1(net501),
    .B2(\device.rxBuffer.buffer[25][1] ),
    .X(_1659_));
 sky130_fd_sc_hd__o211a_1 _3032_ (.A1(net483),
    .A2(_1658_),
    .B1(_1659_),
    .C1(net475),
    .X(_1660_));
 sky130_fd_sc_hd__mux2_1 _3033_ (.A0(\device.rxBuffer.buffer[31][1] ),
    .A1(\device.rxBuffer.buffer[30][1] ),
    .S(net525),
    .X(_1661_));
 sky130_fd_sc_hd__or2_1 _3034_ (.A(net482),
    .B(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__o221a_1 _3035_ (.A1(net514),
    .A2(\device.rxBuffer.buffer[28][1] ),
    .B1(\device.rxBuffer.buffer[29][1] ),
    .B2(net500),
    .C1(net478),
    .X(_1663_));
 sky130_fd_sc_hd__mux2_1 _3036_ (.A0(\device.rxBuffer.buffer[15][1] ),
    .A1(\device.rxBuffer.buffer[14][1] ),
    .S(net523),
    .X(_1664_));
 sky130_fd_sc_hd__o221a_1 _3037_ (.A1(net513),
    .A2(\device.rxBuffer.buffer[12][1] ),
    .B1(net499),
    .B2(\device.rxBuffer.buffer[13][1] ),
    .C1(net476),
    .X(_1665_));
 sky130_fd_sc_hd__o21a_1 _3038_ (.A1(net481),
    .A2(_1664_),
    .B1(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__a21o_1 _3039_ (.A1(\device.rxBuffer.buffer[8][1] ),
    .A2(_1501_),
    .B1(net497),
    .X(_1667_));
 sky130_fd_sc_hd__mux2_1 _3040_ (.A0(\device.rxBuffer.buffer[11][1] ),
    .A1(\device.rxBuffer.buffer[10][1] ),
    .S(net520),
    .X(_1668_));
 sky130_fd_sc_hd__o22a_1 _3041_ (.A1(\device.rxBuffer.buffer[9][1] ),
    .A2(net498),
    .B1(net480),
    .B2(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__a211o_1 _3042_ (.A1(_1667_),
    .A2(_1669_),
    .B1(net454),
    .C1(_1666_),
    .X(_1670_));
 sky130_fd_sc_hd__or3_1 _3043_ (.A(net456),
    .B(_1648_),
    .C(_1651_),
    .X(_1671_));
 sky130_fd_sc_hd__a211o_1 _3044_ (.A1(_1662_),
    .A2(_1663_),
    .B1(net455),
    .C1(_1660_),
    .X(_1672_));
 sky130_fd_sc_hd__o311a_2 _3045_ (.A1(net457),
    .A2(_1654_),
    .A3(_1657_),
    .B1(_1672_),
    .C1(_1517_),
    .X(_1673_));
 sky130_fd_sc_hd__a31o_1 _3046_ (.A1(_1516_),
    .A2(_1670_),
    .A3(_1671_),
    .B1(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__a221o_1 _3047_ (.A1(_1377_),
    .A2(\device.rxBuffer.dataOut[1] ),
    .B1(net435),
    .B2(_1674_),
    .C1(_1528_),
    .X(_1675_));
 sky130_fd_sc_hd__o211a_1 _3048_ (.A1(net618),
    .A2(_1529_),
    .B1(_1675_),
    .C1(net437),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _3049_ (.A0(\device.rxBuffer.buffer[3][0] ),
    .A1(\device.rxBuffer.buffer[2][0] ),
    .S(net521),
    .X(_1676_));
 sky130_fd_sc_hd__o221a_1 _3050_ (.A1(\device.rxBuffer.buffer[0][0] ),
    .A2(_1498_),
    .B1(net499),
    .B2(\device.rxBuffer.buffer[1][0] ),
    .C1(net475),
    .X(_1677_));
 sky130_fd_sc_hd__o21ai_1 _3051_ (.A1(net481),
    .A2(_1676_),
    .B1(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(\device.rxBuffer.buffer[7][0] ),
    .A1(\device.rxBuffer.buffer[6][0] ),
    .S(net522),
    .X(_1679_));
 sky130_fd_sc_hd__o221a_1 _3053_ (.A1(net514),
    .A2(\device.rxBuffer.buffer[4][0] ),
    .B1(net499),
    .B2(\device.rxBuffer.buffer[5][0] ),
    .C1(net477),
    .X(_1680_));
 sky130_fd_sc_hd__o21ai_1 _3054_ (.A1(net481),
    .A2(_1679_),
    .B1(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(\device.rxBuffer.buffer[19][0] ),
    .A1(\device.rxBuffer.buffer[18][0] ),
    .S(net522),
    .X(_1682_));
 sky130_fd_sc_hd__o221a_1 _3056_ (.A1(\device.rxBuffer.buffer[16][0] ),
    .A2(_1498_),
    .B1(net499),
    .B2(\device.rxBuffer.buffer[17][0] ),
    .C1(net475),
    .X(_1683_));
 sky130_fd_sc_hd__o21ai_1 _3057_ (.A1(net481),
    .A2(_1682_),
    .B1(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__mux2_1 _3058_ (.A0(\device.rxBuffer.buffer[23][0] ),
    .A1(\device.rxBuffer.buffer[22][0] ),
    .S(net522),
    .X(_1685_));
 sky130_fd_sc_hd__o221a_1 _3059_ (.A1(\device.rxBuffer.buffer[20][0] ),
    .A2(net513),
    .B1(net499),
    .B2(\device.rxBuffer.buffer[21][0] ),
    .C1(net477),
    .X(_1686_));
 sky130_fd_sc_hd__o21ai_1 _3060_ (.A1(net481),
    .A2(_1685_),
    .B1(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__a31o_1 _3061_ (.A1(_1517_),
    .A2(_1684_),
    .A3(_1687_),
    .B1(net456),
    .X(_1688_));
 sky130_fd_sc_hd__a31o_1 _3062_ (.A1(_1516_),
    .A2(_1678_),
    .A3(_1681_),
    .B1(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(\device.rxBuffer.buffer[15][0] ),
    .A1(\device.rxBuffer.buffer[14][0] ),
    .S(net522),
    .X(_1690_));
 sky130_fd_sc_hd__o221a_1 _3064_ (.A1(net514),
    .A2(\device.rxBuffer.buffer[12][0] ),
    .B1(net499),
    .B2(\device.rxBuffer.buffer[13][0] ),
    .C1(net477),
    .X(_1691_));
 sky130_fd_sc_hd__o21ai_2 _3065_ (.A1(net481),
    .A2(_1690_),
    .B1(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__mux2_1 _3066_ (.A0(\device.rxBuffer.buffer[11][0] ),
    .A1(\device.rxBuffer.buffer[10][0] ),
    .S(net521),
    .X(_1693_));
 sky130_fd_sc_hd__o221a_1 _3067_ (.A1(\device.rxBuffer.buffer[8][0] ),
    .A2(_1498_),
    .B1(net499),
    .B2(\device.rxBuffer.buffer[9][0] ),
    .C1(net473),
    .X(_1694_));
 sky130_fd_sc_hd__o21ai_1 _3068_ (.A1(net481),
    .A2(_1693_),
    .B1(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__mux2_1 _3069_ (.A0(\device.rxBuffer.buffer[27][0] ),
    .A1(\device.rxBuffer.buffer[26][0] ),
    .S(net527),
    .X(_1696_));
 sky130_fd_sc_hd__o221a_1 _3070_ (.A1(\device.rxBuffer.buffer[24][0] ),
    .A2(_1367_),
    .B1(net500),
    .B2(\device.rxBuffer.buffer[25][0] ),
    .C1(net475),
    .X(_1697_));
 sky130_fd_sc_hd__o21ai_1 _3071_ (.A1(net483),
    .A2(_1696_),
    .B1(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(\device.rxBuffer.buffer[31][0] ),
    .A1(\device.rxBuffer.buffer[30][0] ),
    .S(net525),
    .X(_1699_));
 sky130_fd_sc_hd__o221a_1 _3073_ (.A1(net514),
    .A2(\device.rxBuffer.buffer[28][0] ),
    .B1(\device.rxBuffer.buffer[29][0] ),
    .B2(net500),
    .C1(net478),
    .X(_1700_));
 sky130_fd_sc_hd__o21ai_1 _3074_ (.A1(net483),
    .A2(_1699_),
    .B1(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__a31o_2 _3075_ (.A1(_1517_),
    .A2(_1698_),
    .A3(_1701_),
    .B1(net455),
    .X(_1702_));
 sky130_fd_sc_hd__a31o_1 _3076_ (.A1(_1516_),
    .A2(_1692_),
    .A3(_1695_),
    .B1(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__nand2_1 _3077_ (.A(_1689_),
    .B(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__a221o_1 _3078_ (.A1(_1377_),
    .A2(\device.rxBuffer.dataOut[0] ),
    .B1(net435),
    .B2(_1704_),
    .C1(_1528_),
    .X(_1705_));
 sky130_fd_sc_hd__o211a_1 _3079_ (.A1(net622),
    .A2(_1529_),
    .B1(_1705_),
    .C1(net437),
    .X(_0573_));
 sky130_fd_sc_hd__o211a_1 _3080_ (.A1(\device.rxBuffer.lastWriteLostData ),
    .A2(\device.rxBuffer.we_buffered ),
    .B1(net437),
    .C1(_1459_),
    .X(_0572_));
 sky130_fd_sc_hd__nor2_1 _3081_ (.A(_1450_),
    .B(_1459_),
    .Y(_1706_));
 sky130_fd_sc_hd__and2_1 _3082_ (.A(net511),
    .B(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__or2_1 _3083_ (.A(\device.rxBuffer.endPointer[4] ),
    .B(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__nand3_4 _3084_ (.A(\device.rxBuffer.endPointer[4] ),
    .B(net511),
    .C(net512),
    .Y(_1709_));
 sky130_fd_sc_hd__o311a_1 _3085_ (.A1(_1449_),
    .A2(_1459_),
    .A3(_1709_),
    .B1(_1708_),
    .C1(net438),
    .X(_0571_));
 sky130_fd_sc_hd__o21ai_1 _3086_ (.A1(net511),
    .A2(_1706_),
    .B1(net438),
    .Y(_1710_));
 sky130_fd_sc_hd__nor2_1 _3087_ (.A(_1707_),
    .B(_1710_),
    .Y(_0570_));
 sky130_fd_sc_hd__o21ai_1 _3088_ (.A1(net512),
    .A2(_1483_),
    .B1(net438),
    .Y(_1711_));
 sky130_fd_sc_hd__nor2_1 _3089_ (.A(_1706_),
    .B(_1711_),
    .Y(_0569_));
 sky130_fd_sc_hd__o21ai_1 _3090_ (.A1(\device.rxBuffer.endPointer[1] ),
    .A2(_1482_),
    .B1(net438),
    .Y(_1712_));
 sky130_fd_sc_hd__nor2_1 _3091_ (.A(_1483_),
    .B(_1712_),
    .Y(_0568_));
 sky130_fd_sc_hd__o21ai_1 _3092_ (.A1(\device.rxBuffer.endPointer[0] ),
    .A2(_1458_),
    .B1(net438),
    .Y(_1713_));
 sky130_fd_sc_hd__nor2_1 _3093_ (.A(_1482_),
    .B(_1713_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _3094_ (.A(net435),
    .B(_1516_),
    .Y(_1714_));
 sky130_fd_sc_hd__o211a_1 _3095_ (.A1(\device.rxBuffer.startPointer[4] ),
    .A2(net436),
    .B1(_1714_),
    .C1(net439),
    .X(_0566_));
 sky130_fd_sc_hd__o211a_1 _3096_ (.A1(\device.rxBuffer.startPointer[3] ),
    .A2(net435),
    .B1(_1551_),
    .C1(net439),
    .X(_0565_));
 sky130_fd_sc_hd__nand2_1 _3097_ (.A(net436),
    .B(net475),
    .Y(_1715_));
 sky130_fd_sc_hd__o211a_1 _3098_ (.A1(net513),
    .A2(net436),
    .B1(_1715_),
    .C1(net439),
    .X(_0564_));
 sky130_fd_sc_hd__nand2_1 _3099_ (.A(net436),
    .B(net481),
    .Y(_1716_));
 sky130_fd_sc_hd__o211a_1 _3100_ (.A1(net517),
    .A2(net436),
    .B1(_1716_),
    .C1(net438),
    .X(_0563_));
 sky130_fd_sc_hd__o21ai_1 _3101_ (.A1(net521),
    .A2(net436),
    .B1(net438),
    .Y(_1717_));
 sky130_fd_sc_hd__a21oi_1 _3102_ (.A1(net521),
    .A2(net436),
    .B1(_1717_),
    .Y(_0562_));
 sky130_fd_sc_hd__nor2_8 _3103_ (.A(_1461_),
    .B(_1709_),
    .Y(_1718_));
 sky130_fd_sc_hd__mux2_1 _3104_ (.A0(\device.rxBuffer.buffer[28][7] ),
    .A1(net594),
    .S(_1718_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _3105_ (.A0(\device.rxBuffer.buffer[28][6] ),
    .A1(net599),
    .S(_1718_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(\device.rxBuffer.buffer[28][5] ),
    .A1(net605),
    .S(_1718_),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(\device.rxBuffer.buffer[28][4] ),
    .A1(net609),
    .S(_1718_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _3108_ (.A0(\device.rxBuffer.buffer[28][3] ),
    .A1(net612),
    .S(_1718_),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _3109_ (.A0(\device.rxBuffer.buffer[28][2] ),
    .A1(net616),
    .S(_1718_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(\device.rxBuffer.buffer[28][1] ),
    .A1(net620),
    .S(_1718_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _3111_ (.A0(\device.rxBuffer.buffer[28][0] ),
    .A1(net625),
    .S(_1718_),
    .X(_0553_));
 sky130_fd_sc_hd__or3_4 _3112_ (.A(\device.rxBuffer.endPointer[4] ),
    .B(net511),
    .C(net512),
    .X(_1719_));
 sky130_fd_sc_hd__or2_4 _3113_ (.A(_1467_),
    .B(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__mux2_1 _3114_ (.A0(net592),
    .A1(\device.rxBuffer.buffer[2][7] ),
    .S(_1720_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _3115_ (.A0(net597),
    .A1(\device.rxBuffer.buffer[2][6] ),
    .S(_1720_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(net602),
    .A1(\device.rxBuffer.buffer[2][5] ),
    .S(_1720_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _3117_ (.A0(net608),
    .A1(\device.rxBuffer.buffer[2][4] ),
    .S(_1720_),
    .X(_1339_));
 sky130_fd_sc_hd__mux2_1 _3118_ (.A0(net610),
    .A1(\device.rxBuffer.buffer[2][3] ),
    .S(_1720_),
    .X(_1338_));
 sky130_fd_sc_hd__mux2_1 _3119_ (.A0(net614),
    .A1(\device.rxBuffer.buffer[2][2] ),
    .S(_1720_),
    .X(_1337_));
 sky130_fd_sc_hd__mux2_1 _3120_ (.A0(net618),
    .A1(\device.rxBuffer.buffer[2][1] ),
    .S(_1720_),
    .X(_1336_));
 sky130_fd_sc_hd__mux2_1 _3121_ (.A0(net622),
    .A1(\device.rxBuffer.buffer[2][0] ),
    .S(_1720_),
    .X(_1335_));
 sky130_fd_sc_hd__and3_1 _3122_ (.A(_1380_),
    .B(_1381_),
    .C(_1383_),
    .X(_1721_));
 sky130_fd_sc_hd__or4b_2 _3123_ (.A(_1379_),
    .B(_1386_),
    .C(_1388_),
    .D_N(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__clkinv_2 _3124_ (.A(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__nor2_1 _3125_ (.A(_1376_),
    .B(net418),
    .Y(_1724_));
 sky130_fd_sc_hd__nand2_1 _3126_ (.A(net537),
    .B(net546),
    .Y(_1725_));
 sky130_fd_sc_hd__or2_1 _3127_ (.A(net536),
    .B(net546),
    .X(_1726_));
 sky130_fd_sc_hd__nand2_1 _3128_ (.A(_1725_),
    .B(net495),
    .Y(_1727_));
 sky130_fd_sc_hd__a21oi_4 _3129_ (.A1(net534),
    .A2(net541),
    .B1(net530),
    .Y(_1728_));
 sky130_fd_sc_hd__and3_2 _3130_ (.A(\device.txBuffer.startPointer[2] ),
    .B(net534),
    .C(net541),
    .X(_1729_));
 sky130_fd_sc_hd__nor2_4 _3131_ (.A(_1728_),
    .B(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__or2_1 _3132_ (.A(_1728_),
    .B(_1729_),
    .X(_1731_));
 sky130_fd_sc_hd__mux4_1 _3133_ (.A0(\device.txBuffer.buffer[5][7] ),
    .A1(\device.txBuffer.buffer[6][7] ),
    .A2(\device.txBuffer.buffer[7][7] ),
    .A3(\device.txBuffer.buffer[4][7] ),
    .S0(net541),
    .S1(net534),
    .X(_1732_));
 sky130_fd_sc_hd__and2_4 _3134_ (.A(\device.txBuffer.startPointer[3] ),
    .B(_1729_),
    .X(_1733_));
 sky130_fd_sc_hd__xnor2_4 _3135_ (.A(\device.txBuffer.startPointer[4] ),
    .B(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__xor2_4 _3136_ (.A(\device.txBuffer.startPointer[4] ),
    .B(_1733_),
    .X(_1735_));
 sky130_fd_sc_hd__mux4_2 _3137_ (.A0(\device.txBuffer.buffer[1][7] ),
    .A1(\device.txBuffer.buffer[3][7] ),
    .A2(\device.txBuffer.buffer[2][7] ),
    .A3(\device.txBuffer.buffer[0][7] ),
    .S0(net532),
    .S1(net538),
    .X(_1736_));
 sky130_fd_sc_hd__nor2_1 _3138_ (.A(\device.txBuffer.startPointer[3] ),
    .B(_1729_),
    .Y(_1737_));
 sky130_fd_sc_hd__nor2_2 _3139_ (.A(_1733_),
    .B(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__or2_2 _3140_ (.A(_1733_),
    .B(_1737_),
    .X(_1739_));
 sky130_fd_sc_hd__mux4_1 _3141_ (.A0(\device.txBuffer.buffer[17][7] ),
    .A1(\device.txBuffer.buffer[18][7] ),
    .A2(\device.txBuffer.buffer[19][7] ),
    .A3(\device.txBuffer.buffer[16][7] ),
    .S0(net543),
    .S1(net534),
    .X(_1740_));
 sky130_fd_sc_hd__mux4_2 _3142_ (.A0(\device.txBuffer.buffer[21][7] ),
    .A1(\device.txBuffer.buffer[22][7] ),
    .A2(\device.txBuffer.buffer[23][7] ),
    .A3(\device.txBuffer.buffer[20][7] ),
    .S0(net543),
    .S1(net535),
    .X(_1741_));
 sky130_fd_sc_hd__mux4_1 _3143_ (.A0(\device.txBuffer.buffer[13][7] ),
    .A1(\device.txBuffer.buffer[14][7] ),
    .A2(\device.txBuffer.buffer[15][7] ),
    .A3(\device.txBuffer.buffer[12][7] ),
    .S0(net540),
    .S1(net533),
    .X(_1742_));
 sky130_fd_sc_hd__mux4_2 _3144_ (.A0(\device.txBuffer.buffer[9][7] ),
    .A1(\device.txBuffer.buffer[10][7] ),
    .A2(\device.txBuffer.buffer[11][7] ),
    .A3(\device.txBuffer.buffer[8][7] ),
    .S0(net539),
    .S1(net533),
    .X(_1743_));
 sky130_fd_sc_hd__and2_1 _3145_ (.A(net461),
    .B(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__mux4_1 _3146_ (.A0(\device.txBuffer.buffer[29][7] ),
    .A1(\device.txBuffer.buffer[30][7] ),
    .A2(\device.txBuffer.buffer[31][7] ),
    .A3(\device.txBuffer.buffer[28][7] ),
    .S0(net545),
    .S1(net536),
    .X(_1745_));
 sky130_fd_sc_hd__mux4_2 _3147_ (.A0(\device.txBuffer.buffer[25][7] ),
    .A1(\device.txBuffer.buffer[26][7] ),
    .A2(\device.txBuffer.buffer[27][7] ),
    .A3(\device.txBuffer.buffer[24][7] ),
    .S0(net545),
    .S1(net536),
    .X(_1746_));
 sky130_fd_sc_hd__a21o_1 _3148_ (.A1(net465),
    .A2(_1742_),
    .B1(net450),
    .X(_1747_));
 sky130_fd_sc_hd__mux2_1 _3149_ (.A0(_1732_),
    .A1(_1736_),
    .S(net461),
    .X(_1748_));
 sky130_fd_sc_hd__o221a_2 _3150_ (.A1(_1744_),
    .A2(_1747_),
    .B1(_1748_),
    .B2(net452),
    .C1(_1734_),
    .X(_1749_));
 sky130_fd_sc_hd__a21o_1 _3151_ (.A1(net462),
    .A2(_1740_),
    .B1(net452),
    .X(_1750_));
 sky130_fd_sc_hd__a21o_1 _3152_ (.A1(net467),
    .A2(_1741_),
    .B1(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__a21o_1 _3153_ (.A1(net467),
    .A2(_1745_),
    .B1(net451),
    .X(_1752_));
 sky130_fd_sc_hd__a21o_1 _3154_ (.A1(net463),
    .A2(_1746_),
    .B1(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__a31o_1 _3155_ (.A1(_1735_),
    .A2(_1751_),
    .A3(_1753_),
    .B1(_1749_),
    .X(_1754_));
 sky130_fd_sc_hd__and2_4 _3156_ (.A(\device.txBuffer.we_buffered ),
    .B(net418),
    .X(_1755_));
 sky130_fd_sc_hd__nand2_4 _3157_ (.A(\device.txBuffer.we_buffered ),
    .B(net418),
    .Y(_1756_));
 sky130_fd_sc_hd__a22o_1 _3158_ (.A1(\device.txBuffer.dataOut[7] ),
    .A2(_1376_),
    .B1(net413),
    .B2(_1754_),
    .X(_1757_));
 sky130_fd_sc_hd__or2_1 _3159_ (.A(net562),
    .B(_1756_),
    .X(_1758_));
 sky130_fd_sc_hd__o211a_1 _3160_ (.A1(_1755_),
    .A2(_1757_),
    .B1(_1758_),
    .C1(net440),
    .X(_1332_));
 sky130_fd_sc_hd__mux4_1 _3161_ (.A0(\device.txBuffer.buffer[29][6] ),
    .A1(\device.txBuffer.buffer[30][6] ),
    .A2(\device.txBuffer.buffer[31][6] ),
    .A3(\device.txBuffer.buffer[28][6] ),
    .S0(net545),
    .S1(net536),
    .X(_1759_));
 sky130_fd_sc_hd__mux4_2 _3162_ (.A0(\device.txBuffer.buffer[25][6] ),
    .A1(\device.txBuffer.buffer[26][6] ),
    .A2(\device.txBuffer.buffer[27][6] ),
    .A3(\device.txBuffer.buffer[24][6] ),
    .S0(net545),
    .S1(net536),
    .X(_1760_));
 sky130_fd_sc_hd__a21o_1 _3163_ (.A1(net462),
    .A2(_1760_),
    .B1(net450),
    .X(_1761_));
 sky130_fd_sc_hd__a21o_1 _3164_ (.A1(net468),
    .A2(_1759_),
    .B1(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__mux4_2 _3165_ (.A0(\device.txBuffer.buffer[21][6] ),
    .A1(\device.txBuffer.buffer[22][6] ),
    .A2(\device.txBuffer.buffer[23][6] ),
    .A3(\device.txBuffer.buffer[20][6] ),
    .S0(net543),
    .S1(net535),
    .X(_1763_));
 sky130_fd_sc_hd__mux4_2 _3166_ (.A0(\device.txBuffer.buffer[17][6] ),
    .A1(\device.txBuffer.buffer[18][6] ),
    .A2(\device.txBuffer.buffer[19][6] ),
    .A3(\device.txBuffer.buffer[16][6] ),
    .S0(net543),
    .S1(net535),
    .X(_1764_));
 sky130_fd_sc_hd__a21o_1 _3167_ (.A1(net462),
    .A2(_1764_),
    .B1(net452),
    .X(_1765_));
 sky130_fd_sc_hd__a21o_1 _3168_ (.A1(net467),
    .A2(_1763_),
    .B1(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__nand2_1 _3169_ (.A(net412),
    .B(_1734_),
    .Y(_1767_));
 sky130_fd_sc_hd__mux4_1 _3170_ (.A0(\device.txBuffer.buffer[9][6] ),
    .A1(\device.txBuffer.buffer[10][6] ),
    .A2(\device.txBuffer.buffer[11][6] ),
    .A3(\device.txBuffer.buffer[8][6] ),
    .S0(net538),
    .S1(net532),
    .X(_1768_));
 sky130_fd_sc_hd__and2_1 _3171_ (.A(net461),
    .B(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__mux4_2 _3172_ (.A0(\device.txBuffer.buffer[13][6] ),
    .A1(\device.txBuffer.buffer[14][6] ),
    .A2(\device.txBuffer.buffer[15][6] ),
    .A3(\device.txBuffer.buffer[12][6] ),
    .S0(net540),
    .S1(net533),
    .X(_1770_));
 sky130_fd_sc_hd__a21o_1 _3173_ (.A1(net465),
    .A2(_1770_),
    .B1(net450),
    .X(_1771_));
 sky130_fd_sc_hd__mux4_2 _3174_ (.A0(\device.txBuffer.buffer[1][6] ),
    .A1(\device.txBuffer.buffer[3][6] ),
    .A2(\device.txBuffer.buffer[2][6] ),
    .A3(\device.txBuffer.buffer[0][6] ),
    .S0(net532),
    .S1(net539),
    .X(_1772_));
 sky130_fd_sc_hd__mux4_1 _3175_ (.A0(\device.txBuffer.buffer[5][6] ),
    .A1(\device.txBuffer.buffer[6][6] ),
    .A2(\device.txBuffer.buffer[7][6] ),
    .A3(\device.txBuffer.buffer[4][6] ),
    .S0(net540),
    .S1(net532),
    .X(_1773_));
 sky130_fd_sc_hd__mux2_1 _3176_ (.A0(_1772_),
    .A1(_1773_),
    .S(net465),
    .X(_1774_));
 sky130_fd_sc_hd__o221a_2 _3177_ (.A1(_1769_),
    .A2(_1771_),
    .B1(_1774_),
    .B2(net452),
    .C1(_1734_),
    .X(_1775_));
 sky130_fd_sc_hd__a31o_1 _3178_ (.A1(_1735_),
    .A2(_1762_),
    .A3(_1766_),
    .B1(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__a221o_1 _3179_ (.A1(\device.txBuffer.dataOut[6] ),
    .A2(_1376_),
    .B1(net413),
    .B2(_1776_),
    .C1(_1755_),
    .X(_1777_));
 sky130_fd_sc_hd__o211a_1 _3180_ (.A1(net566),
    .A2(_1756_),
    .B1(_1777_),
    .C1(net441),
    .X(_1331_));
 sky130_fd_sc_hd__mux4_2 _3181_ (.A0(\device.txBuffer.buffer[1][5] ),
    .A1(\device.txBuffer.buffer[3][5] ),
    .A2(\device.txBuffer.buffer[2][5] ),
    .A3(\device.txBuffer.buffer[0][5] ),
    .S0(net532),
    .S1(net538),
    .X(_1778_));
 sky130_fd_sc_hd__mux4_2 _3182_ (.A0(\device.txBuffer.buffer[5][5] ),
    .A1(\device.txBuffer.buffer[6][5] ),
    .A2(\device.txBuffer.buffer[7][5] ),
    .A3(\device.txBuffer.buffer[4][5] ),
    .S0(net541),
    .S1(net534),
    .X(_1779_));
 sky130_fd_sc_hd__mux2_1 _3183_ (.A0(_1778_),
    .A1(_1779_),
    .S(net465),
    .X(_1780_));
 sky130_fd_sc_hd__mux4_2 _3184_ (.A0(\device.txBuffer.buffer[9][5] ),
    .A1(\device.txBuffer.buffer[10][5] ),
    .A2(\device.txBuffer.buffer[11][5] ),
    .A3(\device.txBuffer.buffer[8][5] ),
    .S0(net539),
    .S1(net533),
    .X(_1781_));
 sky130_fd_sc_hd__and2_1 _3185_ (.A(net464),
    .B(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__mux4_1 _3186_ (.A0(\device.txBuffer.buffer[13][5] ),
    .A1(\device.txBuffer.buffer[14][5] ),
    .A2(\device.txBuffer.buffer[15][5] ),
    .A3(\device.txBuffer.buffer[12][5] ),
    .S0(net540),
    .S1(net532),
    .X(_1783_));
 sky130_fd_sc_hd__a21o_1 _3187_ (.A1(net465),
    .A2(_1783_),
    .B1(net450),
    .X(_1784_));
 sky130_fd_sc_hd__mux4_2 _3188_ (.A0(\device.txBuffer.buffer[21][5] ),
    .A1(\device.txBuffer.buffer[22][5] ),
    .A2(\device.txBuffer.buffer[23][5] ),
    .A3(\device.txBuffer.buffer[20][5] ),
    .S0(net544),
    .S1(net534),
    .X(_1785_));
 sky130_fd_sc_hd__mux4_2 _3189_ (.A0(\device.txBuffer.buffer[17][5] ),
    .A1(\device.txBuffer.buffer[18][5] ),
    .A2(\device.txBuffer.buffer[19][5] ),
    .A3(\device.txBuffer.buffer[16][5] ),
    .S0(net543),
    .S1(net535),
    .X(_1786_));
 sky130_fd_sc_hd__a21o_1 _3190_ (.A1(net462),
    .A2(_1786_),
    .B1(net453),
    .X(_1787_));
 sky130_fd_sc_hd__a21o_1 _3191_ (.A1(net467),
    .A2(_1785_),
    .B1(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__mux4_1 _3192_ (.A0(\device.txBuffer.buffer[29][5] ),
    .A1(\device.txBuffer.buffer[30][5] ),
    .A2(\device.txBuffer.buffer[31][5] ),
    .A3(\device.txBuffer.buffer[28][5] ),
    .S0(net542),
    .S1(net536),
    .X(_1789_));
 sky130_fd_sc_hd__mux4_2 _3193_ (.A0(\device.txBuffer.buffer[25][5] ),
    .A1(\device.txBuffer.buffer[26][5] ),
    .A2(\device.txBuffer.buffer[27][5] ),
    .A3(\device.txBuffer.buffer[24][5] ),
    .S0(net546),
    .S1(net536),
    .X(_1790_));
 sky130_fd_sc_hd__a21o_1 _3194_ (.A1(net462),
    .A2(_1790_),
    .B1(net450),
    .X(_1791_));
 sky130_fd_sc_hd__a21o_1 _3195_ (.A1(net468),
    .A2(_1789_),
    .B1(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__o221a_2 _3196_ (.A1(net452),
    .A2(_1780_),
    .B1(_1782_),
    .B2(_1784_),
    .C1(_1734_),
    .X(_1793_));
 sky130_fd_sc_hd__a31o_1 _3197_ (.A1(_1735_),
    .A2(_1788_),
    .A3(_1792_),
    .B1(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__a221o_1 _3198_ (.A1(\device.txBuffer.dataOut[5] ),
    .A2(_1376_),
    .B1(net413),
    .B2(_1794_),
    .C1(_1755_),
    .X(_1795_));
 sky130_fd_sc_hd__o211a_1 _3199_ (.A1(net570),
    .A2(_1756_),
    .B1(_1795_),
    .C1(net441),
    .X(_1330_));
 sky130_fd_sc_hd__mux4_2 _3200_ (.A0(\device.txBuffer.buffer[21][4] ),
    .A1(\device.txBuffer.buffer[22][4] ),
    .A2(\device.txBuffer.buffer[23][4] ),
    .A3(\device.txBuffer.buffer[20][4] ),
    .S0(net541),
    .S1(net534),
    .X(_1796_));
 sky130_fd_sc_hd__mux4_1 _3201_ (.A0(\device.txBuffer.buffer[17][4] ),
    .A1(\device.txBuffer.buffer[18][4] ),
    .A2(\device.txBuffer.buffer[19][4] ),
    .A3(\device.txBuffer.buffer[16][4] ),
    .S0(net543),
    .S1(net535),
    .X(_1797_));
 sky130_fd_sc_hd__a21o_1 _3202_ (.A1(net462),
    .A2(_1797_),
    .B1(net453),
    .X(_1798_));
 sky130_fd_sc_hd__a21o_1 _3203_ (.A1(net467),
    .A2(_1796_),
    .B1(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__mux4_1 _3204_ (.A0(\device.txBuffer.buffer[29][4] ),
    .A1(\device.txBuffer.buffer[30][4] ),
    .A2(\device.txBuffer.buffer[31][4] ),
    .A3(\device.txBuffer.buffer[28][4] ),
    .S0(net545),
    .S1(net536),
    .X(_1800_));
 sky130_fd_sc_hd__mux4_1 _3205_ (.A0(\device.txBuffer.buffer[25][4] ),
    .A1(\device.txBuffer.buffer[26][4] ),
    .A2(\device.txBuffer.buffer[27][4] ),
    .A3(\device.txBuffer.buffer[24][4] ),
    .S0(net546),
    .S1(net536),
    .X(_1801_));
 sky130_fd_sc_hd__a21o_1 _3206_ (.A1(net463),
    .A2(_1801_),
    .B1(net451),
    .X(_1802_));
 sky130_fd_sc_hd__a21o_1 _3207_ (.A1(net468),
    .A2(_1800_),
    .B1(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__mux4_2 _3208_ (.A0(\device.txBuffer.buffer[1][4] ),
    .A1(\device.txBuffer.buffer[3][4] ),
    .A2(\device.txBuffer.buffer[2][4] ),
    .A3(\device.txBuffer.buffer[0][4] ),
    .S0(net532),
    .S1(net538),
    .X(_1804_));
 sky130_fd_sc_hd__mux4_2 _3209_ (.A0(\device.txBuffer.buffer[5][4] ),
    .A1(\device.txBuffer.buffer[6][4] ),
    .A2(\device.txBuffer.buffer[7][4] ),
    .A3(\device.txBuffer.buffer[4][4] ),
    .S0(net541),
    .S1(net534),
    .X(_1805_));
 sky130_fd_sc_hd__mux2_1 _3210_ (.A0(_1804_),
    .A1(_1805_),
    .S(net465),
    .X(_1806_));
 sky130_fd_sc_hd__mux4_2 _3211_ (.A0(\device.txBuffer.buffer[13][4] ),
    .A1(\device.txBuffer.buffer[14][4] ),
    .A2(\device.txBuffer.buffer[15][4] ),
    .A3(\device.txBuffer.buffer[12][4] ),
    .S0(net540),
    .S1(net532),
    .X(_1807_));
 sky130_fd_sc_hd__mux4_2 _3212_ (.A0(\device.txBuffer.buffer[9][4] ),
    .A1(\device.txBuffer.buffer[10][4] ),
    .A2(\device.txBuffer.buffer[11][4] ),
    .A3(\device.txBuffer.buffer[8][4] ),
    .S0(net538),
    .S1(net532),
    .X(_1808_));
 sky130_fd_sc_hd__and2_1 _3213_ (.A(net464),
    .B(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__a21o_1 _3214_ (.A1(net466),
    .A2(_1807_),
    .B1(net450),
    .X(_1810_));
 sky130_fd_sc_hd__o221a_2 _3215_ (.A1(net452),
    .A2(_1806_),
    .B1(_1809_),
    .B2(_1810_),
    .C1(_1734_),
    .X(_1811_));
 sky130_fd_sc_hd__a31o_1 _3216_ (.A1(_1735_),
    .A2(_1799_),
    .A3(_1803_),
    .B1(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__a221o_1 _3217_ (.A1(\device.txBuffer.dataOut[4] ),
    .A2(_1376_),
    .B1(net413),
    .B2(_1812_),
    .C1(_1755_),
    .X(_1813_));
 sky130_fd_sc_hd__o211a_1 _3218_ (.A1(net575),
    .A2(_1756_),
    .B1(_1813_),
    .C1(net441),
    .X(_1329_));
 sky130_fd_sc_hd__mux4_2 _3219_ (.A0(\device.txBuffer.buffer[1][3] ),
    .A1(\device.txBuffer.buffer[3][3] ),
    .A2(\device.txBuffer.buffer[2][3] ),
    .A3(\device.txBuffer.buffer[0][3] ),
    .S0(net532),
    .S1(net538),
    .X(_1814_));
 sky130_fd_sc_hd__mux4_2 _3220_ (.A0(\device.txBuffer.buffer[5][3] ),
    .A1(\device.txBuffer.buffer[6][3] ),
    .A2(\device.txBuffer.buffer[7][3] ),
    .A3(\device.txBuffer.buffer[4][3] ),
    .S0(net542),
    .S1(net534),
    .X(_1815_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(\device.txBuffer.buffer[19][3] ),
    .A1(\device.txBuffer.buffer[18][3] ),
    .S(net543),
    .X(_1816_));
 sky130_fd_sc_hd__o22a_1 _3222_ (.A1(\device.txBuffer.buffer[16][3] ),
    .A2(_1728_),
    .B1(_1816_),
    .B2(net470),
    .X(_1817_));
 sky130_fd_sc_hd__o211a_1 _3223_ (.A1(\device.txBuffer.buffer[17][3] ),
    .A2(net494),
    .B1(net462),
    .C1(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__mux2_1 _3224_ (.A0(\device.txBuffer.buffer[23][3] ),
    .A1(\device.txBuffer.buffer[22][3] ),
    .S(net544),
    .X(_1819_));
 sky130_fd_sc_hd__o221a_1 _3225_ (.A1(\device.txBuffer.buffer[20][3] ),
    .A2(net530),
    .B1(net495),
    .B2(\device.txBuffer.buffer[21][3] ),
    .C1(net467),
    .X(_1820_));
 sky130_fd_sc_hd__o21a_1 _3226_ (.A1(net471),
    .A2(_1819_),
    .B1(_1820_),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(\device.txBuffer.buffer[31][3] ),
    .A1(\device.txBuffer.buffer[30][3] ),
    .S(net545),
    .X(_1822_));
 sky130_fd_sc_hd__o221a_1 _3228_ (.A1(net530),
    .A2(\device.txBuffer.buffer[28][3] ),
    .B1(\device.txBuffer.buffer[29][3] ),
    .B2(net495),
    .C1(net468),
    .X(_1823_));
 sky130_fd_sc_hd__o21a_1 _3229_ (.A1(net471),
    .A2(_1822_),
    .B1(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__mux2_1 _3230_ (.A0(\device.txBuffer.buffer[27][3] ),
    .A1(\device.txBuffer.buffer[26][3] ),
    .S(net546),
    .X(_1825_));
 sky130_fd_sc_hd__o22a_1 _3231_ (.A1(\device.txBuffer.buffer[24][3] ),
    .A2(_1728_),
    .B1(_1825_),
    .B2(net470),
    .X(_1826_));
 sky130_fd_sc_hd__o211a_1 _3232_ (.A1(\device.txBuffer.buffer[25][3] ),
    .A2(net494),
    .B1(net463),
    .C1(_1826_),
    .X(_1827_));
 sky130_fd_sc_hd__mux2_1 _3233_ (.A0(\device.txBuffer.buffer[15][3] ),
    .A1(\device.txBuffer.buffer[14][3] ),
    .S(net540),
    .X(_1828_));
 sky130_fd_sc_hd__o221a_1 _3234_ (.A1(\device.txBuffer.buffer[12][3] ),
    .A2(net531),
    .B1(net493),
    .B2(\device.txBuffer.buffer[13][3] ),
    .C1(net465),
    .X(_1829_));
 sky130_fd_sc_hd__o21a_1 _3235_ (.A1(net469),
    .A2(_1828_),
    .B1(_1829_),
    .X(_1830_));
 sky130_fd_sc_hd__mux2_2 _3236_ (.A0(\device.txBuffer.buffer[11][3] ),
    .A1(\device.txBuffer.buffer[10][3] ),
    .S(net538),
    .X(_1831_));
 sky130_fd_sc_hd__or2_1 _3237_ (.A(\device.txBuffer.buffer[9][3] ),
    .B(net493),
    .X(_1832_));
 sky130_fd_sc_hd__o221a_1 _3238_ (.A1(\device.txBuffer.buffer[8][3] ),
    .A2(net510),
    .B1(net469),
    .B2(_1831_),
    .C1(_1832_),
    .X(_1833_));
 sky130_fd_sc_hd__a211o_1 _3239_ (.A1(net461),
    .A2(_1833_),
    .B1(_1830_),
    .C1(net450),
    .X(_1834_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(_1814_),
    .A1(_1815_),
    .S(net465),
    .X(_1835_));
 sky130_fd_sc_hd__o211a_1 _3241_ (.A1(net452),
    .A2(_1835_),
    .B1(_1834_),
    .C1(_1734_),
    .X(_1836_));
 sky130_fd_sc_hd__or3_1 _3242_ (.A(net451),
    .B(_1824_),
    .C(_1827_),
    .X(_1837_));
 sky130_fd_sc_hd__o311a_1 _3243_ (.A1(net453),
    .A2(_1818_),
    .A3(_1821_),
    .B1(_1837_),
    .C1(_1735_),
    .X(_1838_));
 sky130_fd_sc_hd__o21a_1 _3244_ (.A1(_1836_),
    .A2(_1838_),
    .B1(net412),
    .X(_1839_));
 sky130_fd_sc_hd__a211o_1 _3245_ (.A1(\device.txBuffer.dataOut[3] ),
    .A2(_1376_),
    .B1(_1755_),
    .C1(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__o211a_1 _3246_ (.A1(net578),
    .A2(_1756_),
    .B1(_1840_),
    .C1(net441),
    .X(_1328_));
 sky130_fd_sc_hd__mux2_1 _3247_ (.A0(\device.txBuffer.buffer[7][2] ),
    .A1(\device.txBuffer.buffer[6][2] ),
    .S(net541),
    .X(_1841_));
 sky130_fd_sc_hd__o221a_1 _3248_ (.A1(\device.txBuffer.buffer[4][2] ),
    .A2(net531),
    .B1(net496),
    .B2(\device.txBuffer.buffer[5][2] ),
    .C1(net466),
    .X(_1842_));
 sky130_fd_sc_hd__o21a_1 _3249_ (.A1(net472),
    .A2(_1841_),
    .B1(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__mux2_1 _3250_ (.A0(\device.txBuffer.buffer[3][2] ),
    .A1(\device.txBuffer.buffer[2][2] ),
    .S(net539),
    .X(_1844_));
 sky130_fd_sc_hd__o22a_1 _3251_ (.A1(\device.txBuffer.buffer[0][2] ),
    .A2(_1728_),
    .B1(_1844_),
    .B2(net469),
    .X(_1845_));
 sky130_fd_sc_hd__o211a_1 _3252_ (.A1(\device.txBuffer.buffer[1][2] ),
    .A2(net493),
    .B1(net461),
    .C1(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(\device.txBuffer.buffer[19][2] ),
    .A1(\device.txBuffer.buffer[18][2] ),
    .S(net543),
    .X(_1847_));
 sky130_fd_sc_hd__o22a_1 _3254_ (.A1(\device.txBuffer.buffer[16][2] ),
    .A2(net510),
    .B1(net495),
    .B2(\device.txBuffer.buffer[17][2] ),
    .X(_1848_));
 sky130_fd_sc_hd__o211a_1 _3255_ (.A1(net470),
    .A2(_1847_),
    .B1(_1848_),
    .C1(net462),
    .X(_1849_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(\device.txBuffer.buffer[23][2] ),
    .A1(\device.txBuffer.buffer[22][2] ),
    .S(net543),
    .X(_1850_));
 sky130_fd_sc_hd__o221a_1 _3257_ (.A1(\device.txBuffer.buffer[20][2] ),
    .A2(net530),
    .B1(net495),
    .B2(\device.txBuffer.buffer[21][2] ),
    .C1(net467),
    .X(_1851_));
 sky130_fd_sc_hd__o21a_1 _3258_ (.A1(net470),
    .A2(_1850_),
    .B1(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__mux2_1 _3259_ (.A0(\device.txBuffer.buffer[27][2] ),
    .A1(\device.txBuffer.buffer[26][2] ),
    .S(net546),
    .X(_1853_));
 sky130_fd_sc_hd__o22a_1 _3260_ (.A1(\device.txBuffer.buffer[24][2] ),
    .A2(net510),
    .B1(net494),
    .B2(\device.txBuffer.buffer[25][2] ),
    .X(_1854_));
 sky130_fd_sc_hd__o211a_1 _3261_ (.A1(net471),
    .A2(_1853_),
    .B1(_1854_),
    .C1(net463),
    .X(_1855_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(\device.txBuffer.buffer[31][2] ),
    .A1(\device.txBuffer.buffer[30][2] ),
    .S(net545),
    .X(_1856_));
 sky130_fd_sc_hd__or2_1 _3263_ (.A(net471),
    .B(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__o221a_1 _3264_ (.A1(net530),
    .A2(\device.txBuffer.buffer[28][2] ),
    .B1(\device.txBuffer.buffer[29][2] ),
    .B2(net495),
    .C1(net468),
    .X(_1858_));
 sky130_fd_sc_hd__mux2_1 _3265_ (.A0(\device.txBuffer.buffer[15][2] ),
    .A1(\device.txBuffer.buffer[14][2] ),
    .S(net540),
    .X(_1859_));
 sky130_fd_sc_hd__or2_1 _3266_ (.A(net469),
    .B(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__o221a_1 _3267_ (.A1(\device.txBuffer.buffer[12][2] ),
    .A2(net531),
    .B1(net493),
    .B2(\device.txBuffer.buffer[13][2] ),
    .C1(net466),
    .X(_1861_));
 sky130_fd_sc_hd__mux2_1 _3268_ (.A0(\device.txBuffer.buffer[11][2] ),
    .A1(\device.txBuffer.buffer[10][2] ),
    .S(net539),
    .X(_1862_));
 sky130_fd_sc_hd__o22a_1 _3269_ (.A1(\device.txBuffer.buffer[8][2] ),
    .A2(net510),
    .B1(net493),
    .B2(\device.txBuffer.buffer[9][2] ),
    .X(_1863_));
 sky130_fd_sc_hd__o211a_1 _3270_ (.A1(net469),
    .A2(_1862_),
    .B1(_1863_),
    .C1(net461),
    .X(_1864_));
 sky130_fd_sc_hd__a211o_1 _3271_ (.A1(_1860_),
    .A2(_1861_),
    .B1(_1864_),
    .C1(net450),
    .X(_1865_));
 sky130_fd_sc_hd__o311a_1 _3272_ (.A1(net452),
    .A2(_1843_),
    .A3(_1846_),
    .B1(_1865_),
    .C1(_1734_),
    .X(_1866_));
 sky130_fd_sc_hd__a211o_1 _3273_ (.A1(_1857_),
    .A2(_1858_),
    .B1(net451),
    .C1(_1855_),
    .X(_1867_));
 sky130_fd_sc_hd__o311a_1 _3274_ (.A1(net453),
    .A2(_1849_),
    .A3(_1852_),
    .B1(_1867_),
    .C1(_1735_),
    .X(_1868_));
 sky130_fd_sc_hd__o21a_1 _3275_ (.A1(_1866_),
    .A2(_1868_),
    .B1(net412),
    .X(_1869_));
 sky130_fd_sc_hd__a211o_1 _3276_ (.A1(\device.txBuffer.dataOut[2] ),
    .A2(_1376_),
    .B1(_1755_),
    .C1(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__o211a_1 _3277_ (.A1(net583),
    .A2(_1756_),
    .B1(_1870_),
    .C1(net441),
    .X(_1327_));
 sky130_fd_sc_hd__mux2_2 _3278_ (.A0(\device.txBuffer.buffer[3][1] ),
    .A1(\device.txBuffer.buffer[2][1] ),
    .S(net538),
    .X(_1871_));
 sky130_fd_sc_hd__o221a_1 _3279_ (.A1(\device.txBuffer.buffer[0][1] ),
    .A2(net510),
    .B1(net493),
    .B2(\device.txBuffer.buffer[1][1] ),
    .C1(net461),
    .X(_1872_));
 sky130_fd_sc_hd__o21a_2 _3280_ (.A1(net469),
    .A2(_1871_),
    .B1(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__mux2_1 _3281_ (.A0(\device.txBuffer.buffer[7][1] ),
    .A1(\device.txBuffer.buffer[6][1] ),
    .S(net541),
    .X(_1874_));
 sky130_fd_sc_hd__o221a_1 _3282_ (.A1(\device.txBuffer.buffer[4][1] ),
    .A2(net531),
    .B1(net496),
    .B2(\device.txBuffer.buffer[5][1] ),
    .C1(net466),
    .X(_1875_));
 sky130_fd_sc_hd__o21a_1 _3283_ (.A1(net472),
    .A2(_1874_),
    .B1(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__mux2_1 _3284_ (.A0(\device.txBuffer.buffer[19][1] ),
    .A1(\device.txBuffer.buffer[18][1] ),
    .S(net543),
    .X(_1877_));
 sky130_fd_sc_hd__o22a_1 _3285_ (.A1(\device.txBuffer.buffer[16][1] ),
    .A2(net510),
    .B1(net494),
    .B2(\device.txBuffer.buffer[17][1] ),
    .X(_1878_));
 sky130_fd_sc_hd__o211a_1 _3286_ (.A1(net470),
    .A2(_1877_),
    .B1(_1878_),
    .C1(net462),
    .X(_1879_));
 sky130_fd_sc_hd__mux2_1 _3287_ (.A0(\device.txBuffer.buffer[23][1] ),
    .A1(\device.txBuffer.buffer[22][1] ),
    .S(net544),
    .X(_1880_));
 sky130_fd_sc_hd__o221a_1 _3288_ (.A1(\device.txBuffer.buffer[20][1] ),
    .A2(net530),
    .B1(net494),
    .B2(\device.txBuffer.buffer[21][1] ),
    .C1(net467),
    .X(_1881_));
 sky130_fd_sc_hd__o21a_1 _3289_ (.A1(net470),
    .A2(_1880_),
    .B1(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(\device.txBuffer.buffer[27][1] ),
    .A1(\device.txBuffer.buffer[26][1] ),
    .S(net546),
    .X(_1883_));
 sky130_fd_sc_hd__o22a_1 _3291_ (.A1(\device.txBuffer.buffer[24][1] ),
    .A2(net510),
    .B1(net494),
    .B2(\device.txBuffer.buffer[25][1] ),
    .X(_1884_));
 sky130_fd_sc_hd__o211a_1 _3292_ (.A1(net471),
    .A2(_1883_),
    .B1(_1884_),
    .C1(net463),
    .X(_1885_));
 sky130_fd_sc_hd__mux2_1 _3293_ (.A0(\device.txBuffer.buffer[31][1] ),
    .A1(\device.txBuffer.buffer[30][1] ),
    .S(net545),
    .X(_1886_));
 sky130_fd_sc_hd__or2_1 _3294_ (.A(net470),
    .B(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__o221a_1 _3295_ (.A1(net531),
    .A2(\device.txBuffer.buffer[28][1] ),
    .B1(\device.txBuffer.buffer[29][1] ),
    .B2(net494),
    .C1(net468),
    .X(_1888_));
 sky130_fd_sc_hd__mux2_1 _3296_ (.A0(\device.txBuffer.buffer[15][1] ),
    .A1(\device.txBuffer.buffer[14][1] ),
    .S(net540),
    .X(_1889_));
 sky130_fd_sc_hd__or2_1 _3297_ (.A(net469),
    .B(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__o221a_1 _3298_ (.A1(\device.txBuffer.buffer[12][1] ),
    .A2(net531),
    .B1(net496),
    .B2(\device.txBuffer.buffer[13][1] ),
    .C1(net465),
    .X(_1891_));
 sky130_fd_sc_hd__mux2_2 _3299_ (.A0(\device.txBuffer.buffer[11][1] ),
    .A1(\device.txBuffer.buffer[10][1] ),
    .S(net539),
    .X(_1892_));
 sky130_fd_sc_hd__o22a_1 _3300_ (.A1(\device.txBuffer.buffer[8][1] ),
    .A2(net510),
    .B1(net493),
    .B2(\device.txBuffer.buffer[9][1] ),
    .X(_1893_));
 sky130_fd_sc_hd__o211a_1 _3301_ (.A1(net472),
    .A2(_1892_),
    .B1(_1893_),
    .C1(net461),
    .X(_1894_));
 sky130_fd_sc_hd__a211o_1 _3302_ (.A1(_1890_),
    .A2(_1891_),
    .B1(_1894_),
    .C1(net450),
    .X(_1895_));
 sky130_fd_sc_hd__o311a_1 _3303_ (.A1(net452),
    .A2(_1873_),
    .A3(_1876_),
    .B1(_1895_),
    .C1(_1734_),
    .X(_1896_));
 sky130_fd_sc_hd__a211o_1 _3304_ (.A1(_1887_),
    .A2(_1888_),
    .B1(net451),
    .C1(_1885_),
    .X(_1897_));
 sky130_fd_sc_hd__o311a_1 _3305_ (.A1(net453),
    .A2(_1879_),
    .A3(_1882_),
    .B1(_1897_),
    .C1(_1735_),
    .X(_1898_));
 sky130_fd_sc_hd__o21a_1 _3306_ (.A1(_1896_),
    .A2(_1898_),
    .B1(net412),
    .X(_1899_));
 sky130_fd_sc_hd__a211o_1 _3307_ (.A1(\device.txBuffer.dataOut[1] ),
    .A2(_1376_),
    .B1(_1755_),
    .C1(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__o211a_1 _3308_ (.A1(net587),
    .A2(_1756_),
    .B1(_1900_),
    .C1(net440),
    .X(_1326_));
 sky130_fd_sc_hd__mux2_2 _3309_ (.A0(\device.txBuffer.buffer[3][0] ),
    .A1(\device.txBuffer.buffer[2][0] ),
    .S(net538),
    .X(_1901_));
 sky130_fd_sc_hd__o22a_1 _3310_ (.A1(\device.txBuffer.buffer[0][0] ),
    .A2(net510),
    .B1(net493),
    .B2(\device.txBuffer.buffer[1][0] ),
    .X(_1902_));
 sky130_fd_sc_hd__o211a_1 _3311_ (.A1(net469),
    .A2(_1901_),
    .B1(_1902_),
    .C1(net461),
    .X(_1903_));
 sky130_fd_sc_hd__mux2_1 _3312_ (.A0(\device.txBuffer.buffer[7][0] ),
    .A1(\device.txBuffer.buffer[6][0] ),
    .S(net542),
    .X(_1904_));
 sky130_fd_sc_hd__o221a_1 _3313_ (.A1(\device.txBuffer.buffer[4][0] ),
    .A2(net530),
    .B1(net495),
    .B2(\device.txBuffer.buffer[5][0] ),
    .C1(net467),
    .X(_1905_));
 sky130_fd_sc_hd__o21a_1 _3314_ (.A1(net471),
    .A2(_1904_),
    .B1(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(\device.txBuffer.buffer[23][0] ),
    .A1(\device.txBuffer.buffer[22][0] ),
    .S(net544),
    .X(_1907_));
 sky130_fd_sc_hd__o221a_1 _3316_ (.A1(\device.txBuffer.buffer[20][0] ),
    .A2(net530),
    .B1(net495),
    .B2(\device.txBuffer.buffer[21][0] ),
    .C1(net467),
    .X(_1908_));
 sky130_fd_sc_hd__o21a_1 _3317_ (.A1(net470),
    .A2(_1907_),
    .B1(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__mux2_1 _3318_ (.A0(\device.txBuffer.buffer[19][0] ),
    .A1(\device.txBuffer.buffer[18][0] ),
    .S(net544),
    .X(_1910_));
 sky130_fd_sc_hd__o22a_1 _3319_ (.A1(\device.txBuffer.buffer[16][0] ),
    .A2(_1371_),
    .B1(net494),
    .B2(\device.txBuffer.buffer[17][0] ),
    .X(_1911_));
 sky130_fd_sc_hd__o211a_1 _3320_ (.A1(net470),
    .A2(_1910_),
    .B1(_1911_),
    .C1(net462),
    .X(_1912_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(\device.txBuffer.buffer[27][0] ),
    .A1(\device.txBuffer.buffer[26][0] ),
    .S(net545),
    .X(_1913_));
 sky130_fd_sc_hd__o22a_1 _3322_ (.A1(\device.txBuffer.buffer[24][0] ),
    .A2(_1371_),
    .B1(net494),
    .B2(\device.txBuffer.buffer[25][0] ),
    .X(_1914_));
 sky130_fd_sc_hd__o211a_1 _3323_ (.A1(net471),
    .A2(_1913_),
    .B1(_1914_),
    .C1(net463),
    .X(_1915_));
 sky130_fd_sc_hd__mux2_1 _3324_ (.A0(\device.txBuffer.buffer[31][0] ),
    .A1(\device.txBuffer.buffer[30][0] ),
    .S(net545),
    .X(_1916_));
 sky130_fd_sc_hd__or2_1 _3325_ (.A(net470),
    .B(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__o221a_1 _3326_ (.A1(net531),
    .A2(\device.txBuffer.buffer[28][0] ),
    .B1(\device.txBuffer.buffer[29][0] ),
    .B2(net494),
    .C1(net468),
    .X(_1918_));
 sky130_fd_sc_hd__mux2_1 _3327_ (.A0(\device.txBuffer.buffer[15][0] ),
    .A1(\device.txBuffer.buffer[14][0] ),
    .S(net540),
    .X(_1919_));
 sky130_fd_sc_hd__or2_1 _3328_ (.A(net469),
    .B(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__o221a_1 _3329_ (.A1(\device.txBuffer.buffer[12][0] ),
    .A2(net531),
    .B1(net493),
    .B2(\device.txBuffer.buffer[13][0] ),
    .C1(net465),
    .X(_1921_));
 sky130_fd_sc_hd__mux2_2 _3330_ (.A0(\device.txBuffer.buffer[11][0] ),
    .A1(\device.txBuffer.buffer[10][0] ),
    .S(net538),
    .X(_1922_));
 sky130_fd_sc_hd__o22a_1 _3331_ (.A1(\device.txBuffer.buffer[8][0] ),
    .A2(net510),
    .B1(net493),
    .B2(\device.txBuffer.buffer[9][0] ),
    .X(_1923_));
 sky130_fd_sc_hd__o211a_1 _3332_ (.A1(net469),
    .A2(_1922_),
    .B1(_1923_),
    .C1(net461),
    .X(_1924_));
 sky130_fd_sc_hd__a211o_1 _3333_ (.A1(_1920_),
    .A2(_1921_),
    .B1(_1924_),
    .C1(net450),
    .X(_1925_));
 sky130_fd_sc_hd__o311a_2 _3334_ (.A1(net452),
    .A2(_1903_),
    .A3(_1906_),
    .B1(_1925_),
    .C1(_1734_),
    .X(_1926_));
 sky130_fd_sc_hd__a211o_1 _3335_ (.A1(_1917_),
    .A2(_1918_),
    .B1(net451),
    .C1(_1915_),
    .X(_1927_));
 sky130_fd_sc_hd__o311a_1 _3336_ (.A1(net453),
    .A2(_1909_),
    .A3(_1912_),
    .B1(_1927_),
    .C1(_1735_),
    .X(_1928_));
 sky130_fd_sc_hd__o21a_1 _3337_ (.A1(_1926_),
    .A2(_1928_),
    .B1(net412),
    .X(_1929_));
 sky130_fd_sc_hd__a211o_1 _3338_ (.A1(\device.txBuffer.dataOut[0] ),
    .A2(_1376_),
    .B1(_1755_),
    .C1(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__o211a_1 _3339_ (.A1(net591),
    .A2(_1756_),
    .B1(_1930_),
    .C1(net440),
    .X(_1325_));
 sky130_fd_sc_hd__o211a_1 _3340_ (.A1(\device.txBuffer.lastWriteLostData ),
    .A2(\device.txBuffer.we_buffered ),
    .B1(_1394_),
    .C1(_1419_),
    .X(_1324_));
 sky130_fd_sc_hd__nand2_1 _3341_ (.A(net529),
    .B(_1427_),
    .Y(_1931_));
 sky130_fd_sc_hd__a31o_1 _3342_ (.A1(\device.txBuffer.endPointer[3] ),
    .A2(\device.txBuffer.endPointer[2] ),
    .A3(_1427_),
    .B1(\device.txBuffer.endPointer[4] ),
    .X(_1932_));
 sky130_fd_sc_hd__o311a_1 _3343_ (.A1(_1384_),
    .A2(_1394_),
    .A3(_1471_),
    .B1(_1932_),
    .C1(net440),
    .X(_1323_));
 sky130_fd_sc_hd__nand2_1 _3344_ (.A(_1368_),
    .B(_1931_),
    .Y(_1933_));
 sky130_fd_sc_hd__o211a_1 _3345_ (.A1(_1368_),
    .A2(_1931_),
    .B1(_1933_),
    .C1(net1284),
    .X(_1322_));
 sky130_fd_sc_hd__or2_1 _3346_ (.A(net529),
    .B(_1427_),
    .X(_1934_));
 sky130_fd_sc_hd__and3_1 _3347_ (.A(net1284),
    .B(_1931_),
    .C(_1934_),
    .X(_1321_));
 sky130_fd_sc_hd__o21ai_1 _3348_ (.A1(\device.txBuffer.endPointer[1] ),
    .A2(_1395_),
    .B1(net1284),
    .Y(_1935_));
 sky130_fd_sc_hd__nor2_1 _3349_ (.A(_1427_),
    .B(_1935_),
    .Y(_1320_));
 sky130_fd_sc_hd__nand2_1 _3350_ (.A(_1369_),
    .B(_1394_),
    .Y(_1936_));
 sky130_fd_sc_hd__and3b_1 _3351_ (.A_N(_1395_),
    .B(net1284),
    .C(_1936_),
    .X(_1319_));
 sky130_fd_sc_hd__o211a_1 _3352_ (.A1(\device.txBuffer.startPointer[4] ),
    .A2(net412),
    .B1(_1767_),
    .C1(net440),
    .X(_1318_));
 sky130_fd_sc_hd__nand2_1 _3353_ (.A(net413),
    .B(net451),
    .Y(_1937_));
 sky130_fd_sc_hd__o211a_1 _3354_ (.A1(\device.txBuffer.startPointer[3] ),
    .A2(net413),
    .B1(_1937_),
    .C1(net440),
    .X(_1317_));
 sky130_fd_sc_hd__nand2_1 _3355_ (.A(net412),
    .B(net464),
    .Y(_1938_));
 sky130_fd_sc_hd__o211a_1 _3356_ (.A1(net530),
    .A2(net412),
    .B1(_1938_),
    .C1(net440),
    .X(_1316_));
 sky130_fd_sc_hd__nand2_1 _3357_ (.A(net412),
    .B(net471),
    .Y(_1939_));
 sky130_fd_sc_hd__o211a_1 _3358_ (.A1(net534),
    .A2(net412),
    .B1(_1939_),
    .C1(net440),
    .X(_1315_));
 sky130_fd_sc_hd__o21ai_1 _3359_ (.A1(net541),
    .A2(net413),
    .B1(net440),
    .Y(_1940_));
 sky130_fd_sc_hd__a21oi_1 _3360_ (.A1(net541),
    .A2(net413),
    .B1(_1940_),
    .Y(_1314_));
 sky130_fd_sc_hd__or2_4 _3361_ (.A(_1467_),
    .B(_1709_),
    .X(_1941_));
 sky130_fd_sc_hd__mux2_1 _3362_ (.A0(net595),
    .A1(\device.rxBuffer.buffer[30][7] ),
    .S(_1941_),
    .X(_1305_));
 sky130_fd_sc_hd__mux2_1 _3363_ (.A0(net600),
    .A1(\device.rxBuffer.buffer[30][6] ),
    .S(_1941_),
    .X(_1304_));
 sky130_fd_sc_hd__mux2_1 _3364_ (.A0(net605),
    .A1(\device.rxBuffer.buffer[30][5] ),
    .S(_1941_),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_1 _3365_ (.A0(net609),
    .A1(\device.rxBuffer.buffer[30][4] ),
    .S(_1941_),
    .X(_1302_));
 sky130_fd_sc_hd__mux2_1 _3366_ (.A0(net612),
    .A1(\device.rxBuffer.buffer[30][3] ),
    .S(_1941_),
    .X(_1301_));
 sky130_fd_sc_hd__mux2_1 _3367_ (.A0(net616),
    .A1(\device.rxBuffer.buffer[30][2] ),
    .S(_1941_),
    .X(_1300_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(net620),
    .A1(\device.rxBuffer.buffer[30][1] ),
    .S(_1941_),
    .X(_1299_));
 sky130_fd_sc_hd__mux2_1 _3369_ (.A0(net625),
    .A1(\device.rxBuffer.buffer[30][0] ),
    .S(_1941_),
    .X(_1298_));
 sky130_fd_sc_hd__or2_4 _3370_ (.A(_1424_),
    .B(_1471_),
    .X(_1942_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(net563),
    .A1(\device.txBuffer.buffer[28][7] ),
    .S(_1942_),
    .X(_1296_));
 sky130_fd_sc_hd__mux2_1 _3372_ (.A0(net567),
    .A1(\device.txBuffer.buffer[28][6] ),
    .S(_1942_),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_1 _3373_ (.A0(net570),
    .A1(\device.txBuffer.buffer[28][5] ),
    .S(_1942_),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_1 _3374_ (.A0(net573),
    .A1(\device.txBuffer.buffer[28][4] ),
    .S(_1942_),
    .X(_1293_));
 sky130_fd_sc_hd__mux2_1 _3375_ (.A0(net578),
    .A1(\device.txBuffer.buffer[28][3] ),
    .S(_1942_),
    .X(_1292_));
 sky130_fd_sc_hd__mux2_1 _3376_ (.A0(net582),
    .A1(\device.txBuffer.buffer[28][2] ),
    .S(_1942_),
    .X(_1291_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(net585),
    .A1(\device.txBuffer.buffer[28][1] ),
    .S(_1942_),
    .X(_1290_));
 sky130_fd_sc_hd__mux2_1 _3378_ (.A0(net589),
    .A1(\device.txBuffer.buffer[28][0] ),
    .S(_1942_),
    .X(_1289_));
 sky130_fd_sc_hd__nor2_8 _3379_ (.A(_1378_),
    .B(_1433_),
    .Y(_1943_));
 sky130_fd_sc_hd__mux2_1 _3380_ (.A0(\device.txBuffer.buffer[26][7] ),
    .A1(net563),
    .S(_1943_),
    .X(_1288_));
 sky130_fd_sc_hd__mux2_1 _3381_ (.A0(\device.txBuffer.buffer[26][6] ),
    .A1(net567),
    .S(_1943_),
    .X(_1287_));
 sky130_fd_sc_hd__mux2_1 _3382_ (.A0(\device.txBuffer.buffer[26][5] ),
    .A1(net570),
    .S(_1943_),
    .X(_1286_));
 sky130_fd_sc_hd__mux2_1 _3383_ (.A0(\device.txBuffer.buffer[26][4] ),
    .A1(net574),
    .S(_1943_),
    .X(_1285_));
 sky130_fd_sc_hd__mux2_1 _3384_ (.A0(\device.txBuffer.buffer[26][3] ),
    .A1(net577),
    .S(_1943_),
    .X(_1284_));
 sky130_fd_sc_hd__mux2_1 _3385_ (.A0(\device.txBuffer.buffer[26][2] ),
    .A1(net582),
    .S(_1943_),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_1 _3386_ (.A0(\device.txBuffer.buffer[26][1] ),
    .A1(net586),
    .S(_1943_),
    .X(_1282_));
 sky130_fd_sc_hd__mux2_1 _3387_ (.A0(\device.txBuffer.buffer[26][0] ),
    .A1(net590),
    .S(_1943_),
    .X(_1281_));
 sky130_fd_sc_hd__or2_4 _3388_ (.A(_1433_),
    .B(_1435_),
    .X(_1944_));
 sky130_fd_sc_hd__mux2_4 _3389_ (.A0(net560),
    .A1(\device.txBuffer.buffer[2][7] ),
    .S(_1944_),
    .X(_1277_));
 sky130_fd_sc_hd__mux2_4 _3390_ (.A0(net564),
    .A1(\device.txBuffer.buffer[2][6] ),
    .S(_1944_),
    .X(_1276_));
 sky130_fd_sc_hd__mux2_4 _3391_ (.A0(net568),
    .A1(\device.txBuffer.buffer[2][5] ),
    .S(_1944_),
    .X(_1275_));
 sky130_fd_sc_hd__mux2_1 _3392_ (.A0(net572),
    .A1(\device.txBuffer.buffer[2][4] ),
    .S(_1944_),
    .X(_1274_));
 sky130_fd_sc_hd__mux2_1 _3393_ (.A0(net576),
    .A1(\device.txBuffer.buffer[2][3] ),
    .S(_1944_),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_1 _3394_ (.A0(net580),
    .A1(\device.txBuffer.buffer[2][2] ),
    .S(_1944_),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_1 _3395_ (.A0(net584),
    .A1(\device.txBuffer.buffer[2][1] ),
    .S(_1944_),
    .X(_1271_));
 sky130_fd_sc_hd__mux2_1 _3396_ (.A0(net588),
    .A1(\device.txBuffer.buffer[2][0] ),
    .S(_1944_),
    .X(_1270_));
 sky130_fd_sc_hd__nor2_8 _3397_ (.A(_1433_),
    .B(_1471_),
    .Y(_1945_));
 sky130_fd_sc_hd__mux2_1 _3398_ (.A0(\device.txBuffer.buffer[30][7] ),
    .A1(net563),
    .S(_1945_),
    .X(_1269_));
 sky130_fd_sc_hd__mux2_1 _3399_ (.A0(\device.txBuffer.buffer[30][6] ),
    .A1(net567),
    .S(_1945_),
    .X(_1268_));
 sky130_fd_sc_hd__mux2_1 _3400_ (.A0(\device.txBuffer.buffer[30][5] ),
    .A1(net570),
    .S(_1945_),
    .X(_1267_));
 sky130_fd_sc_hd__mux2_1 _3401_ (.A0(\device.txBuffer.buffer[30][4] ),
    .A1(net573),
    .S(_1945_),
    .X(_1266_));
 sky130_fd_sc_hd__mux2_1 _3402_ (.A0(\device.txBuffer.buffer[30][3] ),
    .A1(net579),
    .S(_1945_),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_1 _3403_ (.A0(\device.txBuffer.buffer[30][2] ),
    .A1(net581),
    .S(_1945_),
    .X(_1264_));
 sky130_fd_sc_hd__mux2_1 _3404_ (.A0(\device.txBuffer.buffer[30][1] ),
    .A1(net585),
    .S(_1945_),
    .X(_1263_));
 sky130_fd_sc_hd__mux2_1 _3405_ (.A0(\device.txBuffer.buffer[30][0] ),
    .A1(net589),
    .S(_1945_),
    .X(_1262_));
 sky130_fd_sc_hd__nor2_8 _3406_ (.A(_1378_),
    .B(_1428_),
    .Y(_1946_));
 sky130_fd_sc_hd__mux2_1 _3407_ (.A0(\device.txBuffer.buffer[27][7] ),
    .A1(net563),
    .S(_1946_),
    .X(_1261_));
 sky130_fd_sc_hd__mux2_1 _3408_ (.A0(\device.txBuffer.buffer[27][6] ),
    .A1(net567),
    .S(_1946_),
    .X(_1260_));
 sky130_fd_sc_hd__mux2_1 _3409_ (.A0(\device.txBuffer.buffer[27][5] ),
    .A1(net571),
    .S(_1946_),
    .X(_1259_));
 sky130_fd_sc_hd__mux2_1 _3410_ (.A0(\device.txBuffer.buffer[27][4] ),
    .A1(net574),
    .S(_1946_),
    .X(_1258_));
 sky130_fd_sc_hd__mux2_1 _3411_ (.A0(\device.txBuffer.buffer[27][3] ),
    .A1(net577),
    .S(_1946_),
    .X(_1257_));
 sky130_fd_sc_hd__mux2_1 _3412_ (.A0(\device.txBuffer.buffer[27][2] ),
    .A1(net582),
    .S(_1946_),
    .X(_1256_));
 sky130_fd_sc_hd__mux2_1 _3413_ (.A0(\device.txBuffer.buffer[27][1] ),
    .A1(net586),
    .S(_1946_),
    .X(_1255_));
 sky130_fd_sc_hd__mux2_1 _3414_ (.A0(\device.txBuffer.buffer[27][0] ),
    .A1(net589),
    .S(_1946_),
    .X(_1254_));
 sky130_fd_sc_hd__or3b_4 _3415_ (.A(\device.rxBuffer.endPointer[4] ),
    .B(net512),
    .C_N(net511),
    .X(_1947_));
 sky130_fd_sc_hd__or2_4 _3416_ (.A(_1467_),
    .B(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(net592),
    .A1(\device.rxBuffer.buffer[10][7] ),
    .S(_1948_),
    .X(_1229_));
 sky130_fd_sc_hd__mux2_1 _3418_ (.A0(net597),
    .A1(\device.rxBuffer.buffer[10][6] ),
    .S(_1948_),
    .X(_1228_));
 sky130_fd_sc_hd__mux2_1 _3419_ (.A0(net602),
    .A1(\device.rxBuffer.buffer[10][5] ),
    .S(_1948_),
    .X(_1227_));
 sky130_fd_sc_hd__mux2_1 _3420_ (.A0(net608),
    .A1(\device.rxBuffer.buffer[10][4] ),
    .S(_1948_),
    .X(_1226_));
 sky130_fd_sc_hd__mux2_1 _3421_ (.A0(net610),
    .A1(\device.rxBuffer.buffer[10][3] ),
    .S(_1948_),
    .X(_1225_));
 sky130_fd_sc_hd__mux2_1 _3422_ (.A0(net614),
    .A1(\device.rxBuffer.buffer[10][2] ),
    .S(_1948_),
    .X(_1224_));
 sky130_fd_sc_hd__mux2_1 _3423_ (.A0(net618),
    .A1(\device.rxBuffer.buffer[10][1] ),
    .S(_1948_),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_1 _3424_ (.A0(net622),
    .A1(\device.rxBuffer.buffer[10][0] ),
    .S(_1948_),
    .X(_1222_));
 sky130_fd_sc_hd__nor2_8 _3425_ (.A(net405),
    .B(_1719_),
    .Y(_1949_));
 sky130_fd_sc_hd__mux2_1 _3426_ (.A0(\device.rxBuffer.buffer[0][7] ),
    .A1(net593),
    .S(_1949_),
    .X(_1221_));
 sky130_fd_sc_hd__mux2_1 _3427_ (.A0(\device.rxBuffer.buffer[0][6] ),
    .A1(net597),
    .S(_1949_),
    .X(_1220_));
 sky130_fd_sc_hd__mux2_1 _3428_ (.A0(\device.rxBuffer.buffer[0][5] ),
    .A1(net602),
    .S(_1949_),
    .X(_1219_));
 sky130_fd_sc_hd__mux2_1 _3429_ (.A0(\device.rxBuffer.buffer[0][4] ),
    .A1(net608),
    .S(_1949_),
    .X(_1218_));
 sky130_fd_sc_hd__mux2_1 _3430_ (.A0(\device.rxBuffer.buffer[0][3] ),
    .A1(net610),
    .S(_1949_),
    .X(_1217_));
 sky130_fd_sc_hd__mux2_1 _3431_ (.A0(\device.rxBuffer.buffer[0][2] ),
    .A1(net614),
    .S(_1949_),
    .X(_1216_));
 sky130_fd_sc_hd__mux2_1 _3432_ (.A0(\device.rxBuffer.buffer[0][1] ),
    .A1(net618),
    .S(_1949_),
    .X(_1215_));
 sky130_fd_sc_hd__mux2_1 _3433_ (.A0(\device.rxBuffer.buffer[0][0] ),
    .A1(net622),
    .S(_1949_),
    .X(_1214_));
 sky130_fd_sc_hd__nor2_8 _3434_ (.A(net405),
    .B(_1947_),
    .Y(_1950_));
 sky130_fd_sc_hd__mux2_1 _3435_ (.A0(\device.rxBuffer.buffer[8][7] ),
    .A1(net592),
    .S(_1950_),
    .X(_1213_));
 sky130_fd_sc_hd__mux2_1 _3436_ (.A0(\device.rxBuffer.buffer[8][6] ),
    .A1(net597),
    .S(_1950_),
    .X(_1212_));
 sky130_fd_sc_hd__mux2_1 _3437_ (.A0(\device.rxBuffer.buffer[8][5] ),
    .A1(net602),
    .S(_1950_),
    .X(_1211_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(\device.rxBuffer.buffer[8][4] ),
    .A1(net608),
    .S(_1950_),
    .X(_1210_));
 sky130_fd_sc_hd__mux2_1 _3439_ (.A0(\device.rxBuffer.buffer[8][3] ),
    .A1(net610),
    .S(_1950_),
    .X(_1209_));
 sky130_fd_sc_hd__mux2_1 _3440_ (.A0(\device.rxBuffer.buffer[8][2] ),
    .A1(net614),
    .S(_1950_),
    .X(_1208_));
 sky130_fd_sc_hd__mux2_1 _3441_ (.A0(\device.rxBuffer.buffer[8][1] ),
    .A1(net618),
    .S(_1950_),
    .X(_1207_));
 sky130_fd_sc_hd__mux2_1 _3442_ (.A0(\device.rxBuffer.buffer[8][0] ),
    .A1(net622),
    .S(_1950_),
    .X(_1206_));
 sky130_fd_sc_hd__or3b_4 _3443_ (.A(\device.rxBuffer.endPointer[4] ),
    .B(net511),
    .C_N(net512),
    .X(_1951_));
 sky130_fd_sc_hd__or2_4 _3444_ (.A(_1484_),
    .B(_1951_),
    .X(_1952_));
 sky130_fd_sc_hd__mux2_1 _3445_ (.A0(net592),
    .A1(\device.rxBuffer.buffer[7][7] ),
    .S(_1952_),
    .X(_1205_));
 sky130_fd_sc_hd__mux2_1 _3446_ (.A0(net597),
    .A1(\device.rxBuffer.buffer[7][6] ),
    .S(_1952_),
    .X(_1204_));
 sky130_fd_sc_hd__mux2_1 _3447_ (.A0(net602),
    .A1(\device.rxBuffer.buffer[7][5] ),
    .S(_1952_),
    .X(_1203_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(net606),
    .A1(\device.rxBuffer.buffer[7][4] ),
    .S(_1952_),
    .X(_1202_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(net611),
    .A1(\device.rxBuffer.buffer[7][3] ),
    .S(_1952_),
    .X(_1201_));
 sky130_fd_sc_hd__mux2_1 _3450_ (.A0(net615),
    .A1(\device.rxBuffer.buffer[7][2] ),
    .S(_1952_),
    .X(_1200_));
 sky130_fd_sc_hd__mux2_1 _3451_ (.A0(net619),
    .A1(\device.rxBuffer.buffer[7][1] ),
    .S(_1952_),
    .X(_1199_));
 sky130_fd_sc_hd__mux2_1 _3452_ (.A0(net623),
    .A1(\device.rxBuffer.buffer[7][0] ),
    .S(_1952_),
    .X(_1198_));
 sky130_fd_sc_hd__nand3b_4 _3453_ (.A_N(\device.rxBuffer.endPointer[4] ),
    .B(\device.rxBuffer.endPointer[3] ),
    .C(net512),
    .Y(_1953_));
 sky130_fd_sc_hd__or2_4 _3454_ (.A(_1464_),
    .B(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__mux2_1 _3455_ (.A0(net593),
    .A1(\device.rxBuffer.buffer[13][7] ),
    .S(_1954_),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_1 _3456_ (.A0(net598),
    .A1(\device.rxBuffer.buffer[13][6] ),
    .S(_1954_),
    .X(_1188_));
 sky130_fd_sc_hd__mux2_1 _3457_ (.A0(net603),
    .A1(\device.rxBuffer.buffer[13][5] ),
    .S(_1954_),
    .X(_1187_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(net606),
    .A1(\device.rxBuffer.buffer[13][4] ),
    .S(_1954_),
    .X(_1186_));
 sky130_fd_sc_hd__mux2_1 _3459_ (.A0(net611),
    .A1(\device.rxBuffer.buffer[13][3] ),
    .S(_1954_),
    .X(_1185_));
 sky130_fd_sc_hd__mux2_1 _3460_ (.A0(net615),
    .A1(\device.rxBuffer.buffer[13][2] ),
    .S(_1954_),
    .X(_1184_));
 sky130_fd_sc_hd__mux2_1 _3461_ (.A0(net619),
    .A1(\device.rxBuffer.buffer[13][1] ),
    .S(_1954_),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(net623),
    .A1(\device.rxBuffer.buffer[13][0] ),
    .S(_1954_),
    .X(_1182_));
 sky130_fd_sc_hd__nor2_8 _3463_ (.A(net405),
    .B(_1953_),
    .Y(_1955_));
 sky130_fd_sc_hd__mux2_1 _3464_ (.A0(\device.rxBuffer.buffer[12][7] ),
    .A1(net593),
    .S(_1955_),
    .X(_1181_));
 sky130_fd_sc_hd__mux2_1 _3465_ (.A0(\device.rxBuffer.buffer[12][6] ),
    .A1(net598),
    .S(_1955_),
    .X(_1180_));
 sky130_fd_sc_hd__mux2_1 _3466_ (.A0(\device.rxBuffer.buffer[12][5] ),
    .A1(net603),
    .S(_1955_),
    .X(_1179_));
 sky130_fd_sc_hd__mux2_1 _3467_ (.A0(\device.rxBuffer.buffer[12][4] ),
    .A1(net606),
    .S(_1955_),
    .X(_1178_));
 sky130_fd_sc_hd__mux2_1 _3468_ (.A0(\device.rxBuffer.buffer[12][3] ),
    .A1(net611),
    .S(_1955_),
    .X(_1177_));
 sky130_fd_sc_hd__mux2_1 _3469_ (.A0(\device.rxBuffer.buffer[12][2] ),
    .A1(net615),
    .S(_1955_),
    .X(_1176_));
 sky130_fd_sc_hd__mux2_1 _3470_ (.A0(\device.rxBuffer.buffer[12][1] ),
    .A1(net619),
    .S(_1955_),
    .X(_1175_));
 sky130_fd_sc_hd__mux2_1 _3471_ (.A0(\device.rxBuffer.buffer[12][0] ),
    .A1(net623),
    .S(_1955_),
    .X(_1174_));
 sky130_fd_sc_hd__or2_4 _3472_ (.A(_1467_),
    .B(_1953_),
    .X(_1956_));
 sky130_fd_sc_hd__mux2_1 _3473_ (.A0(net593),
    .A1(\device.rxBuffer.buffer[14][7] ),
    .S(_1956_),
    .X(_1173_));
 sky130_fd_sc_hd__mux2_1 _3474_ (.A0(net598),
    .A1(\device.rxBuffer.buffer[14][6] ),
    .S(_1956_),
    .X(_1172_));
 sky130_fd_sc_hd__mux2_1 _3475_ (.A0(net603),
    .A1(\device.rxBuffer.buffer[14][5] ),
    .S(_1956_),
    .X(_1171_));
 sky130_fd_sc_hd__mux2_1 _3476_ (.A0(net606),
    .A1(\device.rxBuffer.buffer[14][4] ),
    .S(_1956_),
    .X(_1170_));
 sky130_fd_sc_hd__mux2_1 _3477_ (.A0(net611),
    .A1(\device.rxBuffer.buffer[14][3] ),
    .S(_1956_),
    .X(_1169_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(net615),
    .A1(\device.rxBuffer.buffer[14][2] ),
    .S(_1956_),
    .X(_1168_));
 sky130_fd_sc_hd__mux2_1 _3479_ (.A0(net619),
    .A1(\device.rxBuffer.buffer[14][1] ),
    .S(_1956_),
    .X(_1167_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(net623),
    .A1(\device.rxBuffer.buffer[14][0] ),
    .S(_1956_),
    .X(_1166_));
 sky130_fd_sc_hd__or2_4 _3481_ (.A(_1484_),
    .B(_1947_),
    .X(_1957_));
 sky130_fd_sc_hd__mux2_1 _3482_ (.A0(net592),
    .A1(\device.rxBuffer.buffer[11][7] ),
    .S(_1957_),
    .X(_1165_));
 sky130_fd_sc_hd__mux2_1 _3483_ (.A0(net597),
    .A1(\device.rxBuffer.buffer[11][6] ),
    .S(_1957_),
    .X(_1164_));
 sky130_fd_sc_hd__mux2_1 _3484_ (.A0(net602),
    .A1(\device.rxBuffer.buffer[11][5] ),
    .S(_1957_),
    .X(_1163_));
 sky130_fd_sc_hd__mux2_1 _3485_ (.A0(net608),
    .A1(\device.rxBuffer.buffer[11][4] ),
    .S(_1957_),
    .X(_1162_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(net610),
    .A1(\device.rxBuffer.buffer[11][3] ),
    .S(_1957_),
    .X(_1161_));
 sky130_fd_sc_hd__mux2_1 _3487_ (.A0(net614),
    .A1(\device.rxBuffer.buffer[11][2] ),
    .S(_1957_),
    .X(_1160_));
 sky130_fd_sc_hd__mux2_1 _3488_ (.A0(net618),
    .A1(\device.rxBuffer.buffer[11][1] ),
    .S(_1957_),
    .X(_1159_));
 sky130_fd_sc_hd__mux2_1 _3489_ (.A0(net622),
    .A1(\device.rxBuffer.buffer[11][0] ),
    .S(_1957_),
    .X(_1158_));
 sky130_fd_sc_hd__or2_4 _3490_ (.A(_1484_),
    .B(_1719_),
    .X(_1958_));
 sky130_fd_sc_hd__mux2_1 _3491_ (.A0(net592),
    .A1(\device.rxBuffer.buffer[3][7] ),
    .S(_1958_),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_1 _3492_ (.A0(net597),
    .A1(\device.rxBuffer.buffer[3][6] ),
    .S(_1958_),
    .X(_1156_));
 sky130_fd_sc_hd__mux2_1 _3493_ (.A0(net602),
    .A1(\device.rxBuffer.buffer[3][5] ),
    .S(_1958_),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(net608),
    .A1(\device.rxBuffer.buffer[3][4] ),
    .S(_1958_),
    .X(_1154_));
 sky130_fd_sc_hd__mux2_1 _3495_ (.A0(net610),
    .A1(\device.rxBuffer.buffer[3][3] ),
    .S(_1958_),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(net614),
    .A1(\device.rxBuffer.buffer[3][2] ),
    .S(_1958_),
    .X(_1152_));
 sky130_fd_sc_hd__mux2_1 _3497_ (.A0(net618),
    .A1(\device.rxBuffer.buffer[3][1] ),
    .S(_1958_),
    .X(_1151_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(net622),
    .A1(\device.rxBuffer.buffer[3][0] ),
    .S(_1958_),
    .X(_1150_));
 sky130_fd_sc_hd__nor2_8 _3499_ (.A(_1484_),
    .B(_1709_),
    .Y(_1959_));
 sky130_fd_sc_hd__mux2_1 _3500_ (.A0(\device.rxBuffer.buffer[31][7] ),
    .A1(net594),
    .S(_1959_),
    .X(_1149_));
 sky130_fd_sc_hd__mux2_1 _3501_ (.A0(\device.rxBuffer.buffer[31][6] ),
    .A1(net600),
    .S(_1959_),
    .X(_1148_));
 sky130_fd_sc_hd__mux2_1 _3502_ (.A0(\device.rxBuffer.buffer[31][5] ),
    .A1(net605),
    .S(_1959_),
    .X(_1147_));
 sky130_fd_sc_hd__mux2_1 _3503_ (.A0(\device.rxBuffer.buffer[31][4] ),
    .A1(net609),
    .S(_1959_),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(\device.rxBuffer.buffer[31][3] ),
    .A1(net612),
    .S(_1959_),
    .X(_1145_));
 sky130_fd_sc_hd__mux2_1 _3505_ (.A0(\device.rxBuffer.buffer[31][2] ),
    .A1(net616),
    .S(_1959_),
    .X(_1144_));
 sky130_fd_sc_hd__mux2_1 _3506_ (.A0(\device.rxBuffer.buffer[31][1] ),
    .A1(net620),
    .S(_1959_),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_1 _3507_ (.A0(\device.rxBuffer.buffer[31][0] ),
    .A1(net625),
    .S(_1959_),
    .X(_1142_));
 sky130_fd_sc_hd__or2_4 _3508_ (.A(_1467_),
    .B(_1951_),
    .X(_1960_));
 sky130_fd_sc_hd__mux2_1 _3509_ (.A0(net592),
    .A1(\device.rxBuffer.buffer[6][7] ),
    .S(_1960_),
    .X(_1141_));
 sky130_fd_sc_hd__mux2_1 _3510_ (.A0(net597),
    .A1(\device.rxBuffer.buffer[6][6] ),
    .S(_1960_),
    .X(_1140_));
 sky130_fd_sc_hd__mux2_1 _3511_ (.A0(net603),
    .A1(\device.rxBuffer.buffer[6][5] ),
    .S(_1960_),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_1 _3512_ (.A0(net606),
    .A1(\device.rxBuffer.buffer[6][4] ),
    .S(_1960_),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_1 _3513_ (.A0(net610),
    .A1(\device.rxBuffer.buffer[6][3] ),
    .S(_1960_),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_1 _3514_ (.A0(net614),
    .A1(\device.rxBuffer.buffer[6][2] ),
    .S(_1960_),
    .X(_1136_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(net618),
    .A1(\device.rxBuffer.buffer[6][1] ),
    .S(_1960_),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _3516_ (.A0(net623),
    .A1(\device.rxBuffer.buffer[6][0] ),
    .S(_1960_),
    .X(_1134_));
 sky130_fd_sc_hd__nor2_8 _3517_ (.A(_1464_),
    .B(_1951_),
    .Y(_1961_));
 sky130_fd_sc_hd__mux2_1 _3518_ (.A0(\device.rxBuffer.buffer[5][7] ),
    .A1(net592),
    .S(_1961_),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _3519_ (.A0(\device.rxBuffer.buffer[5][6] ),
    .A1(net598),
    .S(_1961_),
    .X(_1132_));
 sky130_fd_sc_hd__mux2_1 _3520_ (.A0(\device.rxBuffer.buffer[5][5] ),
    .A1(net603),
    .S(_1961_),
    .X(_1131_));
 sky130_fd_sc_hd__mux2_1 _3521_ (.A0(\device.rxBuffer.buffer[5][4] ),
    .A1(net606),
    .S(_1961_),
    .X(_1130_));
 sky130_fd_sc_hd__mux2_1 _3522_ (.A0(\device.rxBuffer.buffer[5][3] ),
    .A1(net611),
    .S(_1961_),
    .X(_1129_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(\device.rxBuffer.buffer[5][2] ),
    .A1(net615),
    .S(_1961_),
    .X(_1128_));
 sky130_fd_sc_hd__mux2_1 _3524_ (.A0(\device.rxBuffer.buffer[5][1] ),
    .A1(net619),
    .S(_1961_),
    .X(_1127_));
 sky130_fd_sc_hd__mux2_1 _3525_ (.A0(\device.rxBuffer.buffer[5][0] ),
    .A1(net623),
    .S(_1961_),
    .X(_1126_));
 sky130_fd_sc_hd__nor2_8 _3526_ (.A(net405),
    .B(_1951_),
    .Y(_1962_));
 sky130_fd_sc_hd__mux2_1 _3527_ (.A0(\device.rxBuffer.buffer[4][7] ),
    .A1(net592),
    .S(_1962_),
    .X(_1125_));
 sky130_fd_sc_hd__mux2_1 _3528_ (.A0(\device.rxBuffer.buffer[4][6] ),
    .A1(net598),
    .S(_1962_),
    .X(_1124_));
 sky130_fd_sc_hd__mux2_1 _3529_ (.A0(\device.rxBuffer.buffer[4][5] ),
    .A1(net603),
    .S(_1962_),
    .X(_1123_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(\device.rxBuffer.buffer[4][4] ),
    .A1(net606),
    .S(_1962_),
    .X(_1122_));
 sky130_fd_sc_hd__mux2_1 _3531_ (.A0(\device.rxBuffer.buffer[4][3] ),
    .A1(net611),
    .S(_1962_),
    .X(_1121_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(\device.rxBuffer.buffer[4][2] ),
    .A1(net615),
    .S(_1962_),
    .X(_1120_));
 sky130_fd_sc_hd__mux2_1 _3533_ (.A0(\device.rxBuffer.buffer[4][1] ),
    .A1(net619),
    .S(_1962_),
    .X(_1119_));
 sky130_fd_sc_hd__mux2_1 _3534_ (.A0(\device.rxBuffer.buffer[4][0] ),
    .A1(net623),
    .S(_1962_),
    .X(_1118_));
 sky130_fd_sc_hd__or2_4 _3535_ (.A(_1464_),
    .B(_1709_),
    .X(_1963_));
 sky130_fd_sc_hd__mux2_1 _3536_ (.A0(net595),
    .A1(\device.rxBuffer.buffer[29][7] ),
    .S(_1963_),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_1 _3537_ (.A0(net599),
    .A1(\device.rxBuffer.buffer[29][6] ),
    .S(_1963_),
    .X(_1116_));
 sky130_fd_sc_hd__mux2_1 _3538_ (.A0(net605),
    .A1(\device.rxBuffer.buffer[29][5] ),
    .S(_1963_),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_1 _3539_ (.A0(net609),
    .A1(\device.rxBuffer.buffer[29][4] ),
    .S(_1963_),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_1 _3540_ (.A0(net612),
    .A1(\device.rxBuffer.buffer[29][3] ),
    .S(_1963_),
    .X(_1113_));
 sky130_fd_sc_hd__mux2_1 _3541_ (.A0(net616),
    .A1(\device.rxBuffer.buffer[29][2] ),
    .S(_1963_),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _3542_ (.A0(net620),
    .A1(\device.rxBuffer.buffer[29][1] ),
    .S(_1963_),
    .X(_1111_));
 sky130_fd_sc_hd__mux2_1 _3543_ (.A0(net625),
    .A1(\device.rxBuffer.buffer[29][0] ),
    .S(_1963_),
    .X(_1110_));
 sky130_fd_sc_hd__nor2_8 _3544_ (.A(_1464_),
    .B(_1719_),
    .Y(_1964_));
 sky130_fd_sc_hd__mux2_1 _3545_ (.A0(\device.rxBuffer.buffer[1][7] ),
    .A1(net593),
    .S(_1964_),
    .X(_1109_));
 sky130_fd_sc_hd__mux2_1 _3546_ (.A0(\device.rxBuffer.buffer[1][6] ),
    .A1(net597),
    .S(_1964_),
    .X(_1108_));
 sky130_fd_sc_hd__mux2_1 _3547_ (.A0(\device.rxBuffer.buffer[1][5] ),
    .A1(net602),
    .S(_1964_),
    .X(_1107_));
 sky130_fd_sc_hd__mux2_1 _3548_ (.A0(\device.rxBuffer.buffer[1][4] ),
    .A1(net608),
    .S(_1964_),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_1 _3549_ (.A0(\device.rxBuffer.buffer[1][3] ),
    .A1(net610),
    .S(_1964_),
    .X(_1105_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(\device.rxBuffer.buffer[1][2] ),
    .A1(net614),
    .S(_1964_),
    .X(_1104_));
 sky130_fd_sc_hd__mux2_1 _3551_ (.A0(\device.rxBuffer.buffer[1][1] ),
    .A1(net618),
    .S(_1964_),
    .X(_1103_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(\device.rxBuffer.buffer[1][0] ),
    .A1(net623),
    .S(_1964_),
    .X(_1102_));
 sky130_fd_sc_hd__nor2_8 _3553_ (.A(_1464_),
    .B(_1469_),
    .Y(_1965_));
 sky130_fd_sc_hd__mux2_1 _3554_ (.A0(\device.rxBuffer.buffer[17][7] ),
    .A1(net594),
    .S(_1965_),
    .X(_1053_));
 sky130_fd_sc_hd__mux2_1 _3555_ (.A0(\device.rxBuffer.buffer[17][6] ),
    .A1(net599),
    .S(_1965_),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _3556_ (.A0(\device.rxBuffer.buffer[17][5] ),
    .A1(net604),
    .S(_1965_),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _3557_ (.A0(\device.rxBuffer.buffer[17][4] ),
    .A1(net606),
    .S(_1965_),
    .X(_1050_));
 sky130_fd_sc_hd__mux2_1 _3558_ (.A0(\device.rxBuffer.buffer[17][3] ),
    .A1(net612),
    .S(_1965_),
    .X(_1049_));
 sky130_fd_sc_hd__mux2_1 _3559_ (.A0(\device.rxBuffer.buffer[17][2] ),
    .A1(net616),
    .S(_1965_),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_1 _3560_ (.A0(\device.rxBuffer.buffer[17][1] ),
    .A1(net620),
    .S(_1965_),
    .X(_1047_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(\device.rxBuffer.buffer[17][0] ),
    .A1(net624),
    .S(_1965_),
    .X(_1046_));
 sky130_fd_sc_hd__nor2_8 _3562_ (.A(_1420_),
    .B(_1471_),
    .Y(_1966_));
 sky130_fd_sc_hd__mux2_1 _3563_ (.A0(\device.txBuffer.buffer[29][7] ),
    .A1(net563),
    .S(_1966_),
    .X(_1045_));
 sky130_fd_sc_hd__mux2_1 _3564_ (.A0(\device.txBuffer.buffer[29][6] ),
    .A1(net567),
    .S(_1966_),
    .X(_1044_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(\device.txBuffer.buffer[29][5] ),
    .A1(net570),
    .S(_1966_),
    .X(_1043_));
 sky130_fd_sc_hd__mux2_1 _3566_ (.A0(\device.txBuffer.buffer[29][4] ),
    .A1(net574),
    .S(_1966_),
    .X(_1042_));
 sky130_fd_sc_hd__mux2_1 _3567_ (.A0(\device.txBuffer.buffer[29][3] ),
    .A1(net578),
    .S(_1966_),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_1 _3568_ (.A0(\device.txBuffer.buffer[29][2] ),
    .A1(net582),
    .S(_1966_),
    .X(_1040_));
 sky130_fd_sc_hd__mux2_1 _3569_ (.A0(\device.txBuffer.buffer[29][1] ),
    .A1(net585),
    .S(_1966_),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _3570_ (.A0(\device.txBuffer.buffer[29][0] ),
    .A1(net589),
    .S(_1966_),
    .X(_1038_));
 sky130_fd_sc_hd__or2_4 _3571_ (.A(_1428_),
    .B(_1430_),
    .X(_1967_));
 sky130_fd_sc_hd__mux2_1 _3572_ (.A0(net563),
    .A1(\device.txBuffer.buffer[19][7] ),
    .S(_1967_),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _3573_ (.A0(net566),
    .A1(\device.txBuffer.buffer[19][6] ),
    .S(_1967_),
    .X(_1036_));
 sky130_fd_sc_hd__mux2_1 _3574_ (.A0(net570),
    .A1(\device.txBuffer.buffer[19][5] ),
    .S(_1967_),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _3575_ (.A0(net573),
    .A1(\device.txBuffer.buffer[19][4] ),
    .S(_1967_),
    .X(_1034_));
 sky130_fd_sc_hd__mux2_1 _3576_ (.A0(net577),
    .A1(\device.txBuffer.buffer[19][3] ),
    .S(_1967_),
    .X(_1033_));
 sky130_fd_sc_hd__mux2_1 _3577_ (.A0(net581),
    .A1(\device.txBuffer.buffer[19][2] ),
    .S(_1967_),
    .X(_1032_));
 sky130_fd_sc_hd__mux2_1 _3578_ (.A0(net586),
    .A1(\device.txBuffer.buffer[19][1] ),
    .S(_1967_),
    .X(_1031_));
 sky130_fd_sc_hd__mux2_1 _3579_ (.A0(net589),
    .A1(\device.txBuffer.buffer[19][0] ),
    .S(_1967_),
    .X(_1030_));
 sky130_fd_sc_hd__or2_4 _3580_ (.A(_1469_),
    .B(_1484_),
    .X(_1968_));
 sky130_fd_sc_hd__mux2_1 _3581_ (.A0(net594),
    .A1(\device.rxBuffer.buffer[19][7] ),
    .S(_1968_),
    .X(_1029_));
 sky130_fd_sc_hd__mux2_1 _3582_ (.A0(net599),
    .A1(\device.rxBuffer.buffer[19][6] ),
    .S(_1968_),
    .X(_1028_));
 sky130_fd_sc_hd__mux2_1 _3583_ (.A0(net604),
    .A1(\device.rxBuffer.buffer[19][5] ),
    .S(_1968_),
    .X(_1027_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(net609),
    .A1(\device.rxBuffer.buffer[19][4] ),
    .S(_1968_),
    .X(_1026_));
 sky130_fd_sc_hd__mux2_1 _3585_ (.A0(net612),
    .A1(\device.rxBuffer.buffer[19][3] ),
    .S(_1968_),
    .X(_1025_));
 sky130_fd_sc_hd__mux2_1 _3586_ (.A0(net616),
    .A1(\device.rxBuffer.buffer[19][2] ),
    .S(_1968_),
    .X(_1024_));
 sky130_fd_sc_hd__mux2_1 _3587_ (.A0(net620),
    .A1(\device.rxBuffer.buffer[19][1] ),
    .S(_1968_),
    .X(_1023_));
 sky130_fd_sc_hd__mux2_1 _3588_ (.A0(net622),
    .A1(\device.rxBuffer.buffer[19][0] ),
    .S(_1968_),
    .X(_1022_));
 sky130_fd_sc_hd__nor2_8 _3589_ (.A(_1464_),
    .B(_1947_),
    .Y(_1969_));
 sky130_fd_sc_hd__mux2_1 _3590_ (.A0(\device.rxBuffer.buffer[9][7] ),
    .A1(net592),
    .S(_1969_),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_1 _3591_ (.A0(\device.rxBuffer.buffer[9][6] ),
    .A1(net597),
    .S(_1969_),
    .X(_1020_));
 sky130_fd_sc_hd__mux2_1 _3592_ (.A0(\device.rxBuffer.buffer[9][5] ),
    .A1(net602),
    .S(_1969_),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_1 _3593_ (.A0(\device.rxBuffer.buffer[9][4] ),
    .A1(net608),
    .S(_1969_),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_1 _3594_ (.A0(\device.rxBuffer.buffer[9][3] ),
    .A1(net610),
    .S(_1969_),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_1 _3595_ (.A0(\device.rxBuffer.buffer[9][2] ),
    .A1(net614),
    .S(_1969_),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_1 _3596_ (.A0(\device.rxBuffer.buffer[9][1] ),
    .A1(net618),
    .S(_1969_),
    .X(_1015_));
 sky130_fd_sc_hd__mux2_1 _3597_ (.A0(\device.rxBuffer.buffer[9][0] ),
    .A1(net622),
    .S(_1969_),
    .X(_1014_));
 sky130_fd_sc_hd__nor2_8 _3598_ (.A(_1461_),
    .B(_1469_),
    .Y(_1970_));
 sky130_fd_sc_hd__mux2_1 _3599_ (.A0(\device.rxBuffer.buffer[16][7] ),
    .A1(net594),
    .S(_1970_),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_1 _3600_ (.A0(\device.rxBuffer.buffer[16][6] ),
    .A1(net599),
    .S(_1970_),
    .X(_0969_));
 sky130_fd_sc_hd__mux2_1 _3601_ (.A0(\device.rxBuffer.buffer[16][5] ),
    .A1(net604),
    .S(_1970_),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_1 _3602_ (.A0(\device.rxBuffer.buffer[16][4] ),
    .A1(net607),
    .S(_1970_),
    .X(_0967_));
 sky130_fd_sc_hd__mux2_1 _3603_ (.A0(\device.rxBuffer.buffer[16][3] ),
    .A1(net612),
    .S(_1970_),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_1 _3604_ (.A0(\device.rxBuffer.buffer[16][2] ),
    .A1(net616),
    .S(_1970_),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_1 _3605_ (.A0(\device.rxBuffer.buffer[16][1] ),
    .A1(net620),
    .S(_1970_),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _3606_ (.A0(\device.rxBuffer.buffer[16][0] ),
    .A1(net624),
    .S(_1970_),
    .X(_0963_));
 sky130_fd_sc_hd__nor2_8 _3607_ (.A(_1484_),
    .B(_1953_),
    .Y(_1971_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(\device.rxBuffer.buffer[15][7] ),
    .A1(net593),
    .S(_1971_),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_1 _3609_ (.A0(\device.rxBuffer.buffer[15][6] ),
    .A1(net598),
    .S(_1971_),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _3610_ (.A0(\device.rxBuffer.buffer[15][5] ),
    .A1(net603),
    .S(_1971_),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _3611_ (.A0(\device.rxBuffer.buffer[15][4] ),
    .A1(net606),
    .S(_1971_),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _3612_ (.A0(\device.rxBuffer.buffer[15][3] ),
    .A1(net611),
    .S(_1971_),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _3613_ (.A0(\device.rxBuffer.buffer[15][2] ),
    .A1(net615),
    .S(_1971_),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _3614_ (.A0(\device.rxBuffer.buffer[15][1] ),
    .A1(net619),
    .S(_1971_),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _3615_ (.A0(\device.rxBuffer.buffer[15][0] ),
    .A1(net623),
    .S(_1971_),
    .X(_0955_));
 sky130_fd_sc_hd__and4bb_4 _3616_ (.A_N(\wbAddressExtension.currentAddress[30] ),
    .B_N(\wbAddressExtension.currentAddress[31] ),
    .C(\wbAddressExtension.currentAddress[28] ),
    .D(\wbAddressExtension.currentAddress[29] ),
    .X(_1972_));
 sky130_fd_sc_hd__nand2_1 _3617_ (.A(net487),
    .B(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__and4_4 _3618_ (.A(\wbAddressExtension.currentAddress[24] ),
    .B(\wbAddressExtension.currentAddress[25] ),
    .C(\wbAddressExtension.currentAddress[26] ),
    .D(\wbAddressExtension.currentAddress[27] ),
    .X(_1974_));
 sky130_fd_sc_hd__a31oi_4 _3619_ (.A1(net487),
    .A2(_1972_),
    .A3(_1974_),
    .B1(hostConfigLatch),
    .Y(_1975_));
 sky130_fd_sc_hd__a31o_4 _3620_ (.A1(net487),
    .A2(_1972_),
    .A3(_1974_),
    .B1(hostConfigLatch),
    .X(_1976_));
 sky130_fd_sc_hd__or2_4 _3621_ (.A(_1973_),
    .B(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__inv_2 _3622_ (.A(net433),
    .Y(net235));
 sky130_fd_sc_hd__and2_1 _3623_ (.A(net204),
    .B(net414),
    .X(net272));
 sky130_fd_sc_hd__and2_1 _3624_ (.A(net205),
    .B(net414),
    .X(net273));
 sky130_fd_sc_hd__and2_1 _3625_ (.A(net200),
    .B(net414),
    .X(net268));
 sky130_fd_sc_hd__and2_1 _3626_ (.A(net201),
    .B(net414),
    .X(net269));
 sky130_fd_sc_hd__and2_1 _3627_ (.A(net202),
    .B(net414),
    .X(net270));
 sky130_fd_sc_hd__and2_1 _3628_ (.A(net203),
    .B(net414),
    .X(net271));
 sky130_fd_sc_hd__or2_1 _3629_ (.A(net168),
    .B(net431),
    .X(net236));
 sky130_fd_sc_hd__or2_1 _3630_ (.A(net179),
    .B(net431),
    .X(net247));
 sky130_fd_sc_hd__or2_1 _3631_ (.A(net190),
    .B(net431),
    .X(net258));
 sky130_fd_sc_hd__or2_1 _3632_ (.A(net193),
    .B(net431),
    .X(net261));
 sky130_fd_sc_hd__or2_1 _3633_ (.A(net194),
    .B(net431),
    .X(net262));
 sky130_fd_sc_hd__or2_1 _3634_ (.A(net195),
    .B(net431),
    .X(net263));
 sky130_fd_sc_hd__or2_1 _3635_ (.A(net196),
    .B(net431),
    .X(net264));
 sky130_fd_sc_hd__or2_1 _3636_ (.A(net197),
    .B(net432),
    .X(net265));
 sky130_fd_sc_hd__or2_1 _3637_ (.A(net198),
    .B(net431),
    .X(net266));
 sky130_fd_sc_hd__or2_1 _3638_ (.A(net199),
    .B(net431),
    .X(net267));
 sky130_fd_sc_hd__or2_1 _3639_ (.A(net169),
    .B(net432),
    .X(net237));
 sky130_fd_sc_hd__or2_1 _3640_ (.A(net170),
    .B(net432),
    .X(net238));
 sky130_fd_sc_hd__or2_1 _3641_ (.A(net171),
    .B(net432),
    .X(net239));
 sky130_fd_sc_hd__or2_1 _3642_ (.A(net172),
    .B(net432),
    .X(net240));
 sky130_fd_sc_hd__or2_1 _3643_ (.A(net173),
    .B(net434),
    .X(net241));
 sky130_fd_sc_hd__or2_1 _3644_ (.A(net174),
    .B(net434),
    .X(net242));
 sky130_fd_sc_hd__or2_1 _3645_ (.A(net175),
    .B(net434),
    .X(net243));
 sky130_fd_sc_hd__or2_1 _3646_ (.A(net176),
    .B(net434),
    .X(net244));
 sky130_fd_sc_hd__or2_1 _3647_ (.A(net177),
    .B(net434),
    .X(net245));
 sky130_fd_sc_hd__or2_1 _3648_ (.A(net178),
    .B(net434),
    .X(net246));
 sky130_fd_sc_hd__or2_1 _3649_ (.A(net180),
    .B(net434),
    .X(net248));
 sky130_fd_sc_hd__or2_1 _3650_ (.A(net181),
    .B(net434),
    .X(net249));
 sky130_fd_sc_hd__or2_1 _3651_ (.A(net182),
    .B(net433),
    .X(net250));
 sky130_fd_sc_hd__or2_1 _3652_ (.A(net183),
    .B(net433),
    .X(net251));
 sky130_fd_sc_hd__or2_1 _3653_ (.A(net184),
    .B(net433),
    .X(net252));
 sky130_fd_sc_hd__or2_1 _3654_ (.A(net185),
    .B(net433),
    .X(net253));
 sky130_fd_sc_hd__or2_1 _3655_ (.A(net186),
    .B(net433),
    .X(net254));
 sky130_fd_sc_hd__or2_1 _3656_ (.A(net187),
    .B(net433),
    .X(net255));
 sky130_fd_sc_hd__or2_1 _3657_ (.A(net188),
    .B(net433),
    .X(net256));
 sky130_fd_sc_hd__or2_1 _3658_ (.A(net189),
    .B(net433),
    .X(net257));
 sky130_fd_sc_hd__or2_1 _3659_ (.A(net191),
    .B(net433),
    .X(net259));
 sky130_fd_sc_hd__or2_1 _3660_ (.A(net192),
    .B(net434),
    .X(net260));
 sky130_fd_sc_hd__and2_1 _3661_ (.A(net135),
    .B(net414),
    .X(net207));
 sky130_fd_sc_hd__and2_1 _3662_ (.A(net146),
    .B(net414),
    .X(net218));
 sky130_fd_sc_hd__and2_1 _3663_ (.A(net157),
    .B(net414),
    .X(net227));
 sky130_fd_sc_hd__and2_1 _3664_ (.A(net160),
    .B(net415),
    .X(net228));
 sky130_fd_sc_hd__and2_1 _3665_ (.A(net161),
    .B(net415),
    .X(net229));
 sky130_fd_sc_hd__and2_1 _3666_ (.A(net162),
    .B(net415),
    .X(net230));
 sky130_fd_sc_hd__and2_1 _3667_ (.A(net163),
    .B(net415),
    .X(net231));
 sky130_fd_sc_hd__and2_1 _3668_ (.A(net164),
    .B(net415),
    .X(net232));
 sky130_fd_sc_hd__and2_1 _3669_ (.A(net165),
    .B(net415),
    .X(net233));
 sky130_fd_sc_hd__and2_1 _3670_ (.A(net166),
    .B(net415),
    .X(net234));
 sky130_fd_sc_hd__and2_1 _3671_ (.A(net136),
    .B(net415),
    .X(net208));
 sky130_fd_sc_hd__and2_1 _3672_ (.A(net137),
    .B(net415),
    .X(net209));
 sky130_fd_sc_hd__and2_1 _3673_ (.A(net138),
    .B(net416),
    .X(net210));
 sky130_fd_sc_hd__and2_1 _3674_ (.A(net139),
    .B(net416),
    .X(net211));
 sky130_fd_sc_hd__and2_1 _3675_ (.A(net140),
    .B(net416),
    .X(net212));
 sky130_fd_sc_hd__and2_1 _3676_ (.A(\wbAddressExtension.currentAddress[15] ),
    .B(net416),
    .X(net213));
 sky130_fd_sc_hd__and2_1 _3677_ (.A(\wbAddressExtension.currentAddress[16] ),
    .B(net416),
    .X(net214));
 sky130_fd_sc_hd__and2_1 _3678_ (.A(\wbAddressExtension.currentAddress[17] ),
    .B(net416),
    .X(net215));
 sky130_fd_sc_hd__and2_1 _3679_ (.A(\wbAddressExtension.currentAddress[18] ),
    .B(net416),
    .X(net216));
 sky130_fd_sc_hd__and2_1 _3680_ (.A(\wbAddressExtension.currentAddress[19] ),
    .B(net416),
    .X(net217));
 sky130_fd_sc_hd__and2_1 _3681_ (.A(\wbAddressExtension.currentAddress[20] ),
    .B(net416),
    .X(net219));
 sky130_fd_sc_hd__and2_1 _3682_ (.A(\wbAddressExtension.currentAddress[21] ),
    .B(net416),
    .X(net220));
 sky130_fd_sc_hd__and2_1 _3683_ (.A(\wbAddressExtension.currentAddress[22] ),
    .B(net417),
    .X(net221));
 sky130_fd_sc_hd__and2_1 _3684_ (.A(\wbAddressExtension.currentAddress[23] ),
    .B(net417),
    .X(net222));
 sky130_fd_sc_hd__and2_1 _3685_ (.A(\wbAddressExtension.currentAddress[24] ),
    .B(net417),
    .X(net223));
 sky130_fd_sc_hd__and2_1 _3686_ (.A(\wbAddressExtension.currentAddress[25] ),
    .B(net417),
    .X(net224));
 sky130_fd_sc_hd__and2_1 _3687_ (.A(\wbAddressExtension.currentAddress[26] ),
    .B(net417),
    .X(net225));
 sky130_fd_sc_hd__and2_1 _3688_ (.A(\wbAddressExtension.currentAddress[27] ),
    .B(net417),
    .X(net226));
 sky130_fd_sc_hd__mux2_4 _3689_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[0] ),
    .A1(net3),
    .S(net446),
    .X(_1978_));
 sky130_fd_sc_hd__or2_1 _3690_ (.A(\wbAddressExtension.dataRead_buffered[0] ),
    .B(net638),
    .X(_1979_));
 sky130_fd_sc_hd__o211a_1 _3691_ (.A1(net635),
    .A2(_1978_),
    .B1(_1979_),
    .C1(net1285),
    .X(net373));
 sky130_fd_sc_hd__mux2_4 _3692_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[1] ),
    .A1(net14),
    .S(net446),
    .X(_1980_));
 sky130_fd_sc_hd__or2_1 _3693_ (.A(\wbAddressExtension.dataRead_buffered[1] ),
    .B(net638),
    .X(_1981_));
 sky130_fd_sc_hd__o211a_1 _3694_ (.A1(net635),
    .A2(_1980_),
    .B1(_1981_),
    .C1(net1285),
    .X(net384));
 sky130_fd_sc_hd__mux2_1 _3695_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[2] ),
    .A1(net25),
    .S(net446),
    .X(_1982_));
 sky130_fd_sc_hd__or2_1 _3696_ (.A(\wbAddressExtension.dataRead_buffered[2] ),
    .B(net638),
    .X(_1983_));
 sky130_fd_sc_hd__o211a_2 _3697_ (.A1(net635),
    .A2(_1982_),
    .B1(_1983_),
    .C1(net1283),
    .X(net395));
 sky130_fd_sc_hd__mux2_4 _3698_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[3] ),
    .A1(net28),
    .S(net446),
    .X(_1984_));
 sky130_fd_sc_hd__or2_1 _3699_ (.A(\wbAddressExtension.dataRead_buffered[3] ),
    .B(net638),
    .X(_1985_));
 sky130_fd_sc_hd__o211a_1 _3700_ (.A1(net635),
    .A2(_1984_),
    .B1(_1985_),
    .C1(net1285),
    .X(net398));
 sky130_fd_sc_hd__mux2_4 _3701_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[4] ),
    .A1(net29),
    .S(net446),
    .X(_1986_));
 sky130_fd_sc_hd__or2_1 _3702_ (.A(\wbAddressExtension.dataRead_buffered[4] ),
    .B(net638),
    .X(_1987_));
 sky130_fd_sc_hd__o211a_1 _3703_ (.A1(net635),
    .A2(_1986_),
    .B1(_1987_),
    .C1(net1285),
    .X(net399));
 sky130_fd_sc_hd__mux2_4 _3704_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[5] ),
    .A1(net30),
    .S(net446),
    .X(_1988_));
 sky130_fd_sc_hd__or2_1 _3705_ (.A(\wbAddressExtension.dataRead_buffered[5] ),
    .B(net638),
    .X(_1989_));
 sky130_fd_sc_hd__o211a_1 _3706_ (.A1(net635),
    .A2(_1988_),
    .B1(_1989_),
    .C1(net1285),
    .X(net400));
 sky130_fd_sc_hd__mux2_4 _3707_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[6] ),
    .A1(net31),
    .S(net446),
    .X(_1990_));
 sky130_fd_sc_hd__or2_1 _3708_ (.A(\wbAddressExtension.dataRead_buffered[6] ),
    .B(net638),
    .X(_1991_));
 sky130_fd_sc_hd__o211a_1 _3709_ (.A1(net635),
    .A2(_1990_),
    .B1(_1991_),
    .C1(net502),
    .X(net401));
 sky130_fd_sc_hd__mux2_4 _3710_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[7] ),
    .A1(net32),
    .S(net447),
    .X(_1992_));
 sky130_fd_sc_hd__or2_1 _3711_ (.A(\wbAddressExtension.dataRead_buffered[7] ),
    .B(net638),
    .X(_1993_));
 sky130_fd_sc_hd__o211a_1 _3712_ (.A1(net635),
    .A2(_1992_),
    .B1(_1993_),
    .C1(net1283),
    .X(net402));
 sky130_fd_sc_hd__mux2_4 _3713_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[8] ),
    .A1(net33),
    .S(net446),
    .X(_1994_));
 sky130_fd_sc_hd__or2_1 _3714_ (.A(\wbAddressExtension.dataRead_buffered[8] ),
    .B(net639),
    .X(_1995_));
 sky130_fd_sc_hd__o211a_1 _3715_ (.A1(net635),
    .A2(_1994_),
    .B1(_1995_),
    .C1(net1283),
    .X(net403));
 sky130_fd_sc_hd__mux2_4 _3716_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[9] ),
    .A1(net34),
    .S(net447),
    .X(_1996_));
 sky130_fd_sc_hd__or2_1 _3717_ (.A(\wbAddressExtension.dataRead_buffered[9] ),
    .B(net639),
    .X(_1997_));
 sky130_fd_sc_hd__o211a_1 _3718_ (.A1(net635),
    .A2(_1996_),
    .B1(_1997_),
    .C1(net1283),
    .X(net404));
 sky130_fd_sc_hd__mux2_4 _3719_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[10] ),
    .A1(net4),
    .S(net447),
    .X(_1998_));
 sky130_fd_sc_hd__or2_1 _3720_ (.A(\wbAddressExtension.dataRead_buffered[10] ),
    .B(net639),
    .X(_1999_));
 sky130_fd_sc_hd__o211a_1 _3721_ (.A1(net636),
    .A2(_1998_),
    .B1(_1999_),
    .C1(net503),
    .X(net374));
 sky130_fd_sc_hd__mux2_4 _3722_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[11] ),
    .A1(net5),
    .S(net447),
    .X(_2000_));
 sky130_fd_sc_hd__or2_1 _3723_ (.A(\wbAddressExtension.dataRead_buffered[11] ),
    .B(net639),
    .X(_2001_));
 sky130_fd_sc_hd__o211a_1 _3724_ (.A1(net636),
    .A2(_2000_),
    .B1(_2001_),
    .C1(net503),
    .X(net375));
 sky130_fd_sc_hd__mux2_4 _3725_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[12] ),
    .A1(net6),
    .S(net447),
    .X(_2002_));
 sky130_fd_sc_hd__or2_1 _3726_ (.A(\wbAddressExtension.dataRead_buffered[12] ),
    .B(net639),
    .X(_2003_));
 sky130_fd_sc_hd__o211a_1 _3727_ (.A1(net636),
    .A2(_2002_),
    .B1(_2003_),
    .C1(net503),
    .X(net376));
 sky130_fd_sc_hd__mux2_1 _3728_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[13] ),
    .A1(net7),
    .S(net447),
    .X(_2004_));
 sky130_fd_sc_hd__or2_1 _3729_ (.A(\wbAddressExtension.dataRead_buffered[13] ),
    .B(net639),
    .X(_2005_));
 sky130_fd_sc_hd__o211a_1 _3730_ (.A1(net636),
    .A2(_2004_),
    .B1(_2005_),
    .C1(net503),
    .X(net377));
 sky130_fd_sc_hd__mux2_2 _3731_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[14] ),
    .A1(net8),
    .S(net448),
    .X(_2006_));
 sky130_fd_sc_hd__or2_1 _3732_ (.A(\wbAddressExtension.dataRead_buffered[14] ),
    .B(net141),
    .X(_2007_));
 sky130_fd_sc_hd__o211a_1 _3733_ (.A1(net636),
    .A2(_2006_),
    .B1(_2007_),
    .C1(net506),
    .X(net378));
 sky130_fd_sc_hd__mux2_1 _3734_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[15] ),
    .A1(net9),
    .S(net448),
    .X(_2008_));
 sky130_fd_sc_hd__or2_1 _3735_ (.A(\wbAddressExtension.dataRead_buffered[15] ),
    .B(net640),
    .X(_2009_));
 sky130_fd_sc_hd__o211a_4 _3736_ (.A1(net637),
    .A2(_2008_),
    .B1(_2009_),
    .C1(net504),
    .X(net379));
 sky130_fd_sc_hd__mux2_1 _3737_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[16] ),
    .A1(net10),
    .S(net448),
    .X(_2010_));
 sky130_fd_sc_hd__or2_1 _3738_ (.A(\wbAddressExtension.dataRead_buffered[16] ),
    .B(net640),
    .X(_2011_));
 sky130_fd_sc_hd__o211a_4 _3739_ (.A1(net637),
    .A2(_2010_),
    .B1(_2011_),
    .C1(net504),
    .X(net380));
 sky130_fd_sc_hd__mux2_1 _3740_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[17] ),
    .A1(net11),
    .S(net448),
    .X(_2012_));
 sky130_fd_sc_hd__or2_1 _3741_ (.A(\wbAddressExtension.dataRead_buffered[17] ),
    .B(net640),
    .X(_2013_));
 sky130_fd_sc_hd__o211a_4 _3742_ (.A1(net637),
    .A2(_2012_),
    .B1(_2013_),
    .C1(net504),
    .X(net381));
 sky130_fd_sc_hd__mux2_1 _3743_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[18] ),
    .A1(net12),
    .S(net448),
    .X(_2014_));
 sky130_fd_sc_hd__or2_1 _3744_ (.A(\wbAddressExtension.dataRead_buffered[18] ),
    .B(net640),
    .X(_2015_));
 sky130_fd_sc_hd__o211a_4 _3745_ (.A1(net637),
    .A2(_2014_),
    .B1(_2015_),
    .C1(net504),
    .X(net382));
 sky130_fd_sc_hd__mux2_1 _3746_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[19] ),
    .A1(net13),
    .S(net448),
    .X(_2016_));
 sky130_fd_sc_hd__or2_1 _3747_ (.A(\wbAddressExtension.dataRead_buffered[19] ),
    .B(net640),
    .X(_2017_));
 sky130_fd_sc_hd__o211a_4 _3748_ (.A1(net637),
    .A2(_2016_),
    .B1(_2017_),
    .C1(net504),
    .X(net383));
 sky130_fd_sc_hd__mux2_1 _3749_ (.A0(\wbPeripheralBusInterface.dataRead_buffered[20] ),
    .A1(net15),
    .S(net448),
    .X(_2018_));
 sky130_fd_sc_hd__or2_2 _3750_ (.A(\wbAddressExtension.dataRead_buffered[20] ),
    .B(net640),
    .X(_2019_));
 sky130_fd_sc_hd__o211a_4 _3751_ (.A1(net637),
    .A2(_2018_),
    .B1(_2019_),
    .C1(net504),
    .X(net385));
 sky130_fd_sc_hd__and2_1 _3752_ (.A(net16),
    .B(net448),
    .X(_2020_));
 sky130_fd_sc_hd__a21bo_4 _3753_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[21] ),
    .A2(_1976_),
    .B1_N(net488),
    .X(_2021_));
 sky130_fd_sc_hd__o221a_4 _3754_ (.A1(\wbAddressExtension.dataRead_buffered[21] ),
    .A2(net640),
    .B1(_2020_),
    .B2(net430),
    .C1(net504),
    .X(net386));
 sky130_fd_sc_hd__and2_1 _3755_ (.A(net17),
    .B(net449),
    .X(_2022_));
 sky130_fd_sc_hd__o221a_4 _3756_ (.A1(\wbAddressExtension.dataRead_buffered[22] ),
    .A2(net640),
    .B1(net430),
    .B2(_2022_),
    .C1(net505),
    .X(net387));
 sky130_fd_sc_hd__and2_1 _3757_ (.A(net18),
    .B(net449),
    .X(_2023_));
 sky130_fd_sc_hd__o221a_4 _3758_ (.A1(\wbAddressExtension.dataRead_buffered[23] ),
    .A2(net640),
    .B1(net430),
    .B2(_2023_),
    .C1(net505),
    .X(net388));
 sky130_fd_sc_hd__and2_1 _3759_ (.A(net19),
    .B(net449),
    .X(_2024_));
 sky130_fd_sc_hd__o221a_4 _3760_ (.A1(\wbAddressExtension.dataRead_buffered[24] ),
    .A2(net640),
    .B1(net430),
    .B2(_2024_),
    .C1(net505),
    .X(net389));
 sky130_fd_sc_hd__and2_1 _3761_ (.A(net20),
    .B(net448),
    .X(_2025_));
 sky130_fd_sc_hd__o221a_4 _3762_ (.A1(\wbAddressExtension.dataRead_buffered[25] ),
    .A2(net641),
    .B1(_2021_),
    .B2(_2025_),
    .C1(net504),
    .X(net390));
 sky130_fd_sc_hd__and2_1 _3763_ (.A(net21),
    .B(net448),
    .X(_2026_));
 sky130_fd_sc_hd__o221a_4 _3764_ (.A1(\wbAddressExtension.dataRead_buffered[26] ),
    .A2(net641),
    .B1(net430),
    .B2(_2026_),
    .C1(net504),
    .X(net391));
 sky130_fd_sc_hd__and2_1 _3765_ (.A(net22),
    .B(net449),
    .X(_2027_));
 sky130_fd_sc_hd__o221a_4 _3766_ (.A1(\wbAddressExtension.dataRead_buffered[27] ),
    .A2(net641),
    .B1(net430),
    .B2(_2027_),
    .C1(net504),
    .X(net392));
 sky130_fd_sc_hd__and2_1 _3767_ (.A(net23),
    .B(net449),
    .X(_2028_));
 sky130_fd_sc_hd__o221a_4 _3768_ (.A1(\wbAddressExtension.dataRead_buffered[28] ),
    .A2(net641),
    .B1(net430),
    .B2(_2028_),
    .C1(net505),
    .X(net393));
 sky130_fd_sc_hd__and2_1 _3769_ (.A(net24),
    .B(net449),
    .X(_2029_));
 sky130_fd_sc_hd__o221a_4 _3770_ (.A1(\wbAddressExtension.dataRead_buffered[29] ),
    .A2(net641),
    .B1(net430),
    .B2(_2029_),
    .C1(net505),
    .X(net394));
 sky130_fd_sc_hd__and2_1 _3771_ (.A(net26),
    .B(net449),
    .X(_2030_));
 sky130_fd_sc_hd__o221a_4 _3772_ (.A1(\wbAddressExtension.dataRead_buffered[30] ),
    .A2(net641),
    .B1(net430),
    .B2(_2030_),
    .C1(net505),
    .X(net396));
 sky130_fd_sc_hd__and2_1 _3773_ (.A(net27),
    .B(net449),
    .X(_2031_));
 sky130_fd_sc_hd__o221a_4 _3774_ (.A1(\wbAddressExtension.dataRead_buffered[31] ),
    .A2(net641),
    .B1(net430),
    .B2(_2031_),
    .C1(net505),
    .X(net397));
 sky130_fd_sc_hd__or2_1 _3775_ (.A(\wbPeripheralBusInterface.acknowledge ),
    .B(net446),
    .X(_2032_));
 sky130_fd_sc_hd__o311a_2 _3776_ (.A1(net35),
    .A2(net2),
    .A3(net431),
    .B1(_2032_),
    .C1(net486),
    .X(_2033_));
 sky130_fd_sc_hd__a31o_4 _3777_ (.A1(net637),
    .A2(\wbAddressExtension.acknowledge ),
    .A3(net506),
    .B1(_2033_),
    .X(net372));
 sky130_fd_sc_hd__and3_1 _3778_ (.A(net634),
    .B(net488),
    .C(_1976_),
    .X(_0954_));
 sky130_fd_sc_hd__nand2b_1 _3779_ (.A_N(\wbAddressExtension.state[0] ),
    .B(\wbAddressExtension.state[1] ),
    .Y(_2034_));
 sky130_fd_sc_hd__nand2b_4 _3780_ (.A_N(\wbAddressExtension.state[1] ),
    .B(\wbAddressExtension.state[0] ),
    .Y(_2035_));
 sky130_fd_sc_hd__nor2_8 _3781_ (.A(net642),
    .B(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__or2_4 _3782_ (.A(net642),
    .B(_2035_),
    .X(_2037_));
 sky130_fd_sc_hd__o32a_1 _3783_ (.A1(net3993),
    .A2(\wbAddressExtension.currentAddress[0] ),
    .A3(net553),
    .B1(net489),
    .B2(\wbAddressExtension.dataRead_buffered[0] ),
    .X(_0971_));
 sky130_fd_sc_hd__o32a_1 _3784_ (.A1(net3993),
    .A2(\wbAddressExtension.currentAddress[1] ),
    .A3(net553),
    .B1(net489),
    .B2(\wbAddressExtension.dataRead_buffered[1] ),
    .X(_0972_));
 sky130_fd_sc_hd__o32a_1 _3785_ (.A1(net2731),
    .A2(\wbAddressExtension.currentAddress[2] ),
    .A3(net553),
    .B1(net489),
    .B2(\wbAddressExtension.dataRead_buffered[2] ),
    .X(_0973_));
 sky130_fd_sc_hd__o32a_1 _3786_ (.A1(net3993),
    .A2(\wbAddressExtension.currentAddress[3] ),
    .A3(net553),
    .B1(net489),
    .B2(\wbAddressExtension.dataRead_buffered[3] ),
    .X(_0974_));
 sky130_fd_sc_hd__o32a_1 _3787_ (.A1(net3993),
    .A2(\wbAddressExtension.currentAddress[4] ),
    .A3(net553),
    .B1(net489),
    .B2(\wbAddressExtension.dataRead_buffered[4] ),
    .X(_0975_));
 sky130_fd_sc_hd__o32a_1 _3788_ (.A1(net3993),
    .A2(\wbAddressExtension.currentAddress[5] ),
    .A3(net553),
    .B1(net489),
    .B2(\wbAddressExtension.dataRead_buffered[5] ),
    .X(_0976_));
 sky130_fd_sc_hd__o32a_1 _3789_ (.A1(net3993),
    .A2(\wbAddressExtension.currentAddress[6] ),
    .A3(net553),
    .B1(net489),
    .B2(\wbAddressExtension.dataRead_buffered[6] ),
    .X(_0977_));
 sky130_fd_sc_hd__o32a_1 _3790_ (.A1(net1418),
    .A2(\wbAddressExtension.currentAddress[7] ),
    .A3(net553),
    .B1(net489),
    .B2(\wbAddressExtension.dataRead_buffered[7] ),
    .X(_0978_));
 sky130_fd_sc_hd__o32a_1 _3791_ (.A1(net1418),
    .A2(\wbAddressExtension.currentAddress[8] ),
    .A3(net554),
    .B1(net490),
    .B2(\wbAddressExtension.dataRead_buffered[8] ),
    .X(_0979_));
 sky130_fd_sc_hd__o32a_1 _3792_ (.A1(net1418),
    .A2(\wbAddressExtension.currentAddress[9] ),
    .A3(net554),
    .B1(net490),
    .B2(\wbAddressExtension.dataRead_buffered[9] ),
    .X(_0980_));
 sky130_fd_sc_hd__o32a_1 _3793_ (.A1(net1418),
    .A2(\wbAddressExtension.currentAddress[10] ),
    .A3(net554),
    .B1(net489),
    .B2(\wbAddressExtension.dataRead_buffered[10] ),
    .X(_0981_));
 sky130_fd_sc_hd__o32a_1 _3794_ (.A1(net1418),
    .A2(\wbAddressExtension.currentAddress[11] ),
    .A3(net554),
    .B1(net490),
    .B2(\wbAddressExtension.dataRead_buffered[11] ),
    .X(_0982_));
 sky130_fd_sc_hd__o32a_1 _3795_ (.A1(net1418),
    .A2(\wbAddressExtension.currentAddress[12] ),
    .A3(net554),
    .B1(net490),
    .B2(\wbAddressExtension.dataRead_buffered[12] ),
    .X(_0983_));
 sky130_fd_sc_hd__o32a_1 _3796_ (.A1(net1418),
    .A2(\wbAddressExtension.currentAddress[13] ),
    .A3(net554),
    .B1(net489),
    .B2(\wbAddressExtension.dataRead_buffered[13] ),
    .X(_0984_));
 sky130_fd_sc_hd__o32a_1 _3797_ (.A1(net1466),
    .A2(\wbAddressExtension.currentAddress[14] ),
    .A3(net557),
    .B1(net1645),
    .B2(\wbAddressExtension.dataRead_buffered[14] ),
    .X(_0985_));
 sky130_fd_sc_hd__o32a_1 _3798_ (.A1(net1558),
    .A2(\wbAddressExtension.currentAddress[15] ),
    .A3(net555),
    .B1(net1630),
    .B2(\wbAddressExtension.dataRead_buffered[15] ),
    .X(_0986_));
 sky130_fd_sc_hd__o32a_1 _3799_ (.A1(net1558),
    .A2(\wbAddressExtension.currentAddress[16] ),
    .A3(net555),
    .B1(net1630),
    .B2(\wbAddressExtension.dataRead_buffered[16] ),
    .X(_0987_));
 sky130_fd_sc_hd__o32a_1 _3800_ (.A1(net1558),
    .A2(\wbAddressExtension.currentAddress[17] ),
    .A3(net555),
    .B1(net1630),
    .B2(\wbAddressExtension.dataRead_buffered[17] ),
    .X(_0988_));
 sky130_fd_sc_hd__o32a_1 _3801_ (.A1(net1558),
    .A2(\wbAddressExtension.currentAddress[18] ),
    .A3(net555),
    .B1(net1630),
    .B2(\wbAddressExtension.dataRead_buffered[18] ),
    .X(_0989_));
 sky130_fd_sc_hd__o32a_1 _3802_ (.A1(net1558),
    .A2(\wbAddressExtension.currentAddress[19] ),
    .A3(net555),
    .B1(net1630),
    .B2(\wbAddressExtension.dataRead_buffered[19] ),
    .X(_0990_));
 sky130_fd_sc_hd__o32a_1 _3803_ (.A1(net1558),
    .A2(\wbAddressExtension.currentAddress[20] ),
    .A3(net555),
    .B1(net1630),
    .B2(\wbAddressExtension.dataRead_buffered[20] ),
    .X(_0991_));
 sky130_fd_sc_hd__o32a_1 _3804_ (.A1(net1558),
    .A2(\wbAddressExtension.currentAddress[21] ),
    .A3(net555),
    .B1(net1630),
    .B2(\wbAddressExtension.dataRead_buffered[21] ),
    .X(_0992_));
 sky130_fd_sc_hd__o32a_1 _3805_ (.A1(net1558),
    .A2(\wbAddressExtension.currentAddress[22] ),
    .A3(net556),
    .B1(net492),
    .B2(\wbAddressExtension.dataRead_buffered[22] ),
    .X(_0993_));
 sky130_fd_sc_hd__o32a_1 _3806_ (.A1(net1558),
    .A2(\wbAddressExtension.currentAddress[23] ),
    .A3(net556),
    .B1(net492),
    .B2(\wbAddressExtension.dataRead_buffered[23] ),
    .X(_0994_));
 sky130_fd_sc_hd__o32a_1 _3807_ (.A1(\wbAddressExtension.currentAddress[24] ),
    .A2(net1558),
    .A3(net556),
    .B1(net492),
    .B2(\wbAddressExtension.dataRead_buffered[24] ),
    .X(_0995_));
 sky130_fd_sc_hd__o32a_1 _3808_ (.A1(\wbAddressExtension.currentAddress[25] ),
    .A2(net1639),
    .A3(net555),
    .B1(net1630),
    .B2(\wbAddressExtension.dataRead_buffered[25] ),
    .X(_0996_));
 sky130_fd_sc_hd__o32a_1 _3809_ (.A1(\wbAddressExtension.currentAddress[26] ),
    .A2(net1639),
    .A3(net555),
    .B1(net1630),
    .B2(\wbAddressExtension.dataRead_buffered[26] ),
    .X(_0997_));
 sky130_fd_sc_hd__o32a_1 _3810_ (.A1(\wbAddressExtension.currentAddress[27] ),
    .A2(net1639),
    .A3(net555),
    .B1(net1630),
    .B2(\wbAddressExtension.dataRead_buffered[27] ),
    .X(_0998_));
 sky130_fd_sc_hd__o32a_1 _3811_ (.A1(\wbAddressExtension.currentAddress[28] ),
    .A2(net1639),
    .A3(net556),
    .B1(net492),
    .B2(\wbAddressExtension.dataRead_buffered[28] ),
    .X(_0999_));
 sky130_fd_sc_hd__o32a_1 _3812_ (.A1(\wbAddressExtension.currentAddress[29] ),
    .A2(net1639),
    .A3(net556),
    .B1(net492),
    .B2(\wbAddressExtension.dataRead_buffered[29] ),
    .X(_1000_));
 sky130_fd_sc_hd__o32a_1 _3813_ (.A1(\wbAddressExtension.currentAddress[30] ),
    .A2(net1639),
    .A3(net556),
    .B1(net492),
    .B2(\wbAddressExtension.dataRead_buffered[30] ),
    .X(_1001_));
 sky130_fd_sc_hd__o32a_1 _3814_ (.A1(\wbAddressExtension.currentAddress[31] ),
    .A2(net1639),
    .A3(net556),
    .B1(net492),
    .B2(\wbAddressExtension.dataRead_buffered[31] ),
    .X(_1002_));
 sky130_fd_sc_hd__nand2_8 _3815_ (.A(net1350),
    .B(net1357),
    .Y(_2038_));
 sky130_fd_sc_hd__mux2_1 _3816_ (.A0(net168),
    .A1(\wbAddressExtension.currentAddress[0] ),
    .S(net1361),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _3817_ (.A0(net179),
    .A1(\wbAddressExtension.currentAddress[1] ),
    .S(net1361),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _3818_ (.A0(net190),
    .A1(\wbAddressExtension.currentAddress[2] ),
    .S(net1361),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_1 _3819_ (.A0(net193),
    .A1(\wbAddressExtension.currentAddress[3] ),
    .S(net1361),
    .X(_1006_));
 sky130_fd_sc_hd__mux2_1 _3820_ (.A0(net194),
    .A1(\wbAddressExtension.currentAddress[4] ),
    .S(net1361),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_1 _3821_ (.A0(net195),
    .A1(\wbAddressExtension.currentAddress[5] ),
    .S(net1361),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_1 _3822_ (.A0(net196),
    .A1(\wbAddressExtension.currentAddress[6] ),
    .S(net1361),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _3823_ (.A0(net197),
    .A1(\wbAddressExtension.currentAddress[7] ),
    .S(net1361),
    .X(_1010_));
 sky130_fd_sc_hd__a31o_1 _3824_ (.A1(net637),
    .A2(net1580),
    .A3(net502),
    .B1(\wbAddressExtension.state[0] ),
    .X(_2039_));
 sky130_fd_sc_hd__o21a_1 _3825_ (.A1(\wbAddressExtension.state[1] ),
    .A2(net3112),
    .B1(net632),
    .X(_2040_));
 sky130_fd_sc_hd__nand2_1 _3826_ (.A(\wbAddressExtension.state[1] ),
    .B(\wbAddressExtension.state[0] ),
    .Y(_2041_));
 sky130_fd_sc_hd__or3_1 _3827_ (.A(\wbAddressExtension.state[1] ),
    .B(\wbAddressExtension.state[0] ),
    .C(net2329),
    .X(_2042_));
 sky130_fd_sc_hd__and3_1 _3828_ (.A(net3116),
    .B(_2041_),
    .C(net2331),
    .X(_1011_));
 sky130_fd_sc_hd__and3_1 _3829_ (.A(net553),
    .B(_2035_),
    .C(net2331),
    .X(_2043_));
 sky130_fd_sc_hd__and2b_1 _3830_ (.A_N(_2043_),
    .B(net3116),
    .X(_1012_));
 sky130_fd_sc_hd__a31oi_4 _3831_ (.A1(net179),
    .A2(net1971),
    .A3(net459),
    .B1(net3863),
    .Y(_2044_));
 sky130_fd_sc_hd__a31o_1 _3832_ (.A1(net179),
    .A2(net1971),
    .A3(net459),
    .B1(net3863),
    .X(_2045_));
 sky130_fd_sc_hd__mux4_1 _3833_ (.A0(\device.uartTx.savedData[0] ),
    .A1(\device.uartTx.savedData[1] ),
    .A2(\device.uartTx.savedData[2] ),
    .A3(\device.uartTx.savedData[3] ),
    .S0(\device.uartTx.bitCounter[0] ),
    .S1(\device.uartTx.bitCounter[1] ),
    .X(_2046_));
 sky130_fd_sc_hd__and2b_1 _3834_ (.A_N(\device.uartTx.bitCounter[2] ),
    .B(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__mux4_2 _3835_ (.A0(\device.uartTx.savedData[4] ),
    .A1(\device.uartTx.savedData[5] ),
    .A2(\device.uartTx.savedData[6] ),
    .A3(\device.uartTx.savedData[7] ),
    .S0(\device.uartTx.bitCounter[0] ),
    .S1(\device.uartTx.bitCounter[1] ),
    .X(_2048_));
 sky130_fd_sc_hd__or2_1 _3836_ (.A(_1364_),
    .B(\device.uartTx.state[0] ),
    .X(_2049_));
 sky130_fd_sc_hd__nor2_8 _3837_ (.A(\device.uartTx.state[1] ),
    .B(\device.uartTx.state[0] ),
    .Y(_2050_));
 sky130_fd_sc_hd__or2_4 _3838_ (.A(\device.uartTx.state[1] ),
    .B(\device.uartTx.state[0] ),
    .X(_2051_));
 sky130_fd_sc_hd__a211o_1 _3839_ (.A1(\device.uartTx.bitCounter[2] ),
    .A2(_2048_),
    .B1(_2047_),
    .C1(\device.uartTx.state[0] ),
    .X(_2052_));
 sky130_fd_sc_hd__a211o_4 _3840_ (.A1(\device.uartTx.state[1] ),
    .A2(_2052_),
    .B1(_2050_),
    .C1(net1984),
    .X(_1013_));
 sky130_fd_sc_hd__nor2_2 _3841_ (.A(_1372_),
    .B(net631),
    .Y(_2053_));
 sky130_fd_sc_hd__or3_2 _3842_ (.A(\wbPeripheralBusInterface.currentAddress[2] ),
    .B(\wbPeripheralBusInterface.currentAddress[10] ),
    .C(\wbPeripheralBusInterface.currentAddress[11] ),
    .X(_2054_));
 sky130_fd_sc_hd__or3_2 _3843_ (.A(\wbPeripheralBusInterface.currentAddress[3] ),
    .B(_1414_),
    .C(_2054_),
    .X(_2055_));
 sky130_fd_sc_hd__or3_4 _3844_ (.A(_1372_),
    .B(net631),
    .C(_2055_),
    .X(_2056_));
 sky130_fd_sc_hd__nor2_1 _3845_ (.A(_1410_),
    .B(_2056_),
    .Y(_2057_));
 sky130_fd_sc_hd__or2_4 _3846_ (.A(_1410_),
    .B(_2056_),
    .X(_2058_));
 sky130_fd_sc_hd__a31o_1 _3847_ (.A1(\device.configuration[0] ),
    .A2(net627),
    .A3(net558),
    .B1(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__o21a_1 _3848_ (.A1(\wbPeripheralBusInterface.currentAddress[3] ),
    .A2(_2054_),
    .B1(_1407_),
    .X(_2060_));
 sky130_fd_sc_hd__nand2_1 _3849_ (.A(\wbPeripheralBusInterface.currentAddress[3] ),
    .B(_2053_),
    .Y(_2061_));
 sky130_fd_sc_hd__or4_4 _3850_ (.A(_1410_),
    .B(_1414_),
    .C(_2054_),
    .D(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__or3b_4 _3851_ (.A(\wbPeripheralBusInterface.currentAddress[5] ),
    .B(_1409_),
    .C_N(\wbPeripheralBusInterface.currentAddress[4] ),
    .X(_2063_));
 sky130_fd_sc_hd__or2_1 _3852_ (.A(_1416_),
    .B(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__o31a_4 _3853_ (.A1(_1372_),
    .A2(net631),
    .A3(_2064_),
    .B1(_2062_),
    .X(_2065_));
 sky130_fd_sc_hd__nor2_1 _3854_ (.A(_2056_),
    .B(_2063_),
    .Y(_2066_));
 sky130_fd_sc_hd__or2_4 _3855_ (.A(_2056_),
    .B(_2063_),
    .X(_2067_));
 sky130_fd_sc_hd__a31o_1 _3856_ (.A1(net627),
    .A2(\device.rxRegister.baseReadData[0] ),
    .A3(net558),
    .B1(_2067_),
    .X(_2068_));
 sky130_fd_sc_hd__nor2_4 _3857_ (.A(_1408_),
    .B(_2062_),
    .Y(_2069_));
 sky130_fd_sc_hd__a221o_1 _3858_ (.A1(_2065_),
    .A2(_2068_),
    .B1(_2069_),
    .B2(\device.statusRegister.baseReadData[0] ),
    .C1(net426),
    .X(_2070_));
 sky130_fd_sc_hd__a31o_1 _3859_ (.A1(net507),
    .A2(_2059_),
    .A3(_2070_),
    .B1(net3863),
    .X(_2071_));
 sky130_fd_sc_hd__a21o_1 _3860_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[0] ),
    .A2(net509),
    .B1(net3436),
    .X(_1054_));
 sky130_fd_sc_hd__a31o_1 _3861_ (.A1(\device.configuration[1] ),
    .A2(net627),
    .A3(net558),
    .B1(_2058_),
    .X(_2072_));
 sky130_fd_sc_hd__a31o_1 _3862_ (.A1(net627),
    .A2(\device.rxRegister.baseReadData[1] ),
    .A3(net558),
    .B1(_2067_),
    .X(_2073_));
 sky130_fd_sc_hd__a221o_1 _3863_ (.A1(\device.statusRegister.baseReadData[1] ),
    .A2(_2069_),
    .B1(_2073_),
    .B2(_2065_),
    .C1(net426),
    .X(_2074_));
 sky130_fd_sc_hd__a31o_1 _3864_ (.A1(net507),
    .A2(_2072_),
    .A3(_2074_),
    .B1(net3863),
    .X(_2075_));
 sky130_fd_sc_hd__a21o_1 _3865_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[1] ),
    .A2(net509),
    .B1(net3409),
    .X(_1055_));
 sky130_fd_sc_hd__a31o_1 _3866_ (.A1(\device.configuration[2] ),
    .A2(net627),
    .A3(net558),
    .B1(_2058_),
    .X(_2076_));
 sky130_fd_sc_hd__a31o_1 _3867_ (.A1(net627),
    .A2(\device.rxRegister.baseReadData[2] ),
    .A3(net558),
    .B1(_2067_),
    .X(_2077_));
 sky130_fd_sc_hd__a221o_1 _3868_ (.A1(\device.statusRegister.baseReadData[2] ),
    .A2(_2069_),
    .B1(_2077_),
    .B2(_2065_),
    .C1(net426),
    .X(_2078_));
 sky130_fd_sc_hd__a31o_1 _3869_ (.A1(net507),
    .A2(_2076_),
    .A3(_2078_),
    .B1(net3863),
    .X(_2079_));
 sky130_fd_sc_hd__a21o_1 _3870_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[2] ),
    .A2(net509),
    .B1(net3400),
    .X(_1056_));
 sky130_fd_sc_hd__a31o_1 _3871_ (.A1(\device.configuration[3] ),
    .A2(net628),
    .A3(net559),
    .B1(_2058_),
    .X(_2080_));
 sky130_fd_sc_hd__a31o_1 _3872_ (.A1(net628),
    .A2(\device.rxRegister.baseReadData[3] ),
    .A3(net559),
    .B1(_2067_),
    .X(_2081_));
 sky130_fd_sc_hd__a221o_1 _3873_ (.A1(\device.statusRegister.baseReadData[3] ),
    .A2(_2069_),
    .B1(_2081_),
    .B2(_2065_),
    .C1(net426),
    .X(_2082_));
 sky130_fd_sc_hd__a31o_1 _3874_ (.A1(_1397_),
    .A2(_2080_),
    .A3(_2082_),
    .B1(net3863),
    .X(_2083_));
 sky130_fd_sc_hd__a21o_1 _3875_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[3] ),
    .A2(net509),
    .B1(net3418),
    .X(_1057_));
 sky130_fd_sc_hd__a31o_1 _3876_ (.A1(\device.configuration[4] ),
    .A2(net627),
    .A3(net558),
    .B1(_2058_),
    .X(_2084_));
 sky130_fd_sc_hd__a31o_1 _3877_ (.A1(net627),
    .A2(\device.rxRegister.baseReadData[4] ),
    .A3(net558),
    .B1(_2067_),
    .X(_2085_));
 sky130_fd_sc_hd__a221o_1 _3878_ (.A1(\device.statusRegister.baseReadData[4] ),
    .A2(_2069_),
    .B1(_2085_),
    .B2(_2065_),
    .C1(net426),
    .X(_2086_));
 sky130_fd_sc_hd__a31o_1 _3879_ (.A1(net507),
    .A2(_2084_),
    .A3(_2086_),
    .B1(net1835),
    .X(_2087_));
 sky130_fd_sc_hd__a21o_1 _3880_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[4] ),
    .A2(net509),
    .B1(net1807),
    .X(_1058_));
 sky130_fd_sc_hd__a31o_1 _3881_ (.A1(\device.configuration[5] ),
    .A2(net627),
    .A3(net558),
    .B1(_2058_),
    .X(_2088_));
 sky130_fd_sc_hd__a31o_1 _3882_ (.A1(net628),
    .A2(\device.rxRegister.baseReadData[5] ),
    .A3(net558),
    .B1(_2067_),
    .X(_2089_));
 sky130_fd_sc_hd__a221o_1 _3883_ (.A1(\device.statusRegister.baseReadData[5] ),
    .A2(_2069_),
    .B1(_2089_),
    .B2(_2065_),
    .C1(net426),
    .X(_2090_));
 sky130_fd_sc_hd__a31o_1 _3884_ (.A1(net507),
    .A2(_2088_),
    .A3(_2090_),
    .B1(net3863),
    .X(_2091_));
 sky130_fd_sc_hd__a21o_1 _3885_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[5] ),
    .A2(net509),
    .B1(net3427),
    .X(_1059_));
 sky130_fd_sc_hd__a31o_1 _3886_ (.A1(net628),
    .A2(\device.rxRegister.baseReadData[6] ),
    .A3(net559),
    .B1(_2067_),
    .X(_2092_));
 sky130_fd_sc_hd__and2_2 _3887_ (.A(_2058_),
    .B(_2065_),
    .X(_2093_));
 sky130_fd_sc_hd__nor3_1 _3888_ (.A(_1408_),
    .B(_1410_),
    .C(_2056_),
    .Y(_2094_));
 sky130_fd_sc_hd__a22o_1 _3889_ (.A1(_2092_),
    .A2(_2093_),
    .B1(_2094_),
    .B2(\device.configuration[6] ),
    .X(_2095_));
 sky130_fd_sc_hd__a31o_1 _3890_ (.A1(_1372_),
    .A2(net631),
    .A3(\wbPeripheralBusInterface.dataRead_buffered[6] ),
    .B1(net1835),
    .X(_2096_));
 sky130_fd_sc_hd__a21o_1 _3891_ (.A1(net507),
    .A2(_2095_),
    .B1(net1817),
    .X(_1060_));
 sky130_fd_sc_hd__a31o_1 _3892_ (.A1(net628),
    .A2(\device.rxRegister.baseReadData[7] ),
    .A3(net559),
    .B1(_2067_),
    .X(_2097_));
 sky130_fd_sc_hd__a22o_1 _3893_ (.A1(\device.configuration[7] ),
    .A2(_2094_),
    .B1(_2097_),
    .B2(_2093_),
    .X(_2098_));
 sky130_fd_sc_hd__a31o_1 _3894_ (.A1(_1372_),
    .A2(net631),
    .A3(\wbPeripheralBusInterface.dataRead_buffered[7] ),
    .B1(net1835),
    .X(_2099_));
 sky130_fd_sc_hd__a21o_1 _3895_ (.A1(net507),
    .A2(_2098_),
    .B1(net1836),
    .X(_1061_));
 sky130_fd_sc_hd__a31o_1 _3896_ (.A1(net626),
    .A2(\device.rxDataAvailableBuffered ),
    .A3(net559),
    .B1(_2067_),
    .X(_2100_));
 sky130_fd_sc_hd__and3_1 _3897_ (.A(\device.configuration[8] ),
    .B(net626),
    .C(net559),
    .X(_2101_));
 sky130_fd_sc_hd__a22o_1 _3898_ (.A1(_2093_),
    .A2(_2100_),
    .B1(_2101_),
    .B2(net426),
    .X(_2102_));
 sky130_fd_sc_hd__a31o_1 _3899_ (.A1(_1372_),
    .A2(net631),
    .A3(\wbPeripheralBusInterface.dataRead_buffered[8] ),
    .B1(net1835),
    .X(_2103_));
 sky130_fd_sc_hd__a21o_1 _3900_ (.A1(net507),
    .A2(_2102_),
    .B1(_2103_),
    .X(_1062_));
 sky130_fd_sc_hd__a31o_4 _3901_ (.A1(_1397_),
    .A2(_2067_),
    .A3(_2093_),
    .B1(net1835),
    .X(_2104_));
 sky130_fd_sc_hd__and3_1 _3902_ (.A(\device.configuration[9] ),
    .B(net629),
    .C(net626),
    .X(_2105_));
 sky130_fd_sc_hd__a221o_1 _3903_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[9] ),
    .A2(net508),
    .B1(net426),
    .B2(_2105_),
    .C1(net411),
    .X(_1063_));
 sky130_fd_sc_hd__and3_1 _3904_ (.A(\device.configuration[10] ),
    .B(net629),
    .C(net626),
    .X(_2106_));
 sky130_fd_sc_hd__a221o_1 _3905_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[10] ),
    .A2(net508),
    .B1(net425),
    .B2(_2106_),
    .C1(net411),
    .X(_1064_));
 sky130_fd_sc_hd__and3_1 _3906_ (.A(\device.configuration[11] ),
    .B(net629),
    .C(net626),
    .X(_2107_));
 sky130_fd_sc_hd__a221o_1 _3907_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[11] ),
    .A2(net508),
    .B1(net425),
    .B2(_2107_),
    .C1(net411),
    .X(_1065_));
 sky130_fd_sc_hd__and3_1 _3908_ (.A(\device.configuration[12] ),
    .B(net629),
    .C(net626),
    .X(_2108_));
 sky130_fd_sc_hd__a221o_1 _3909_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[12] ),
    .A2(net508),
    .B1(net425),
    .B2(_2108_),
    .C1(net411),
    .X(_1066_));
 sky130_fd_sc_hd__and3_1 _3910_ (.A(\device.configuration[13] ),
    .B(net629),
    .C(net626),
    .X(_2109_));
 sky130_fd_sc_hd__a221o_1 _3911_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[13] ),
    .A2(net508),
    .B1(net425),
    .B2(_2109_),
    .C1(net411),
    .X(_1067_));
 sky130_fd_sc_hd__and3_1 _3912_ (.A(\device.configuration[14] ),
    .B(net629),
    .C(net626),
    .X(_2110_));
 sky130_fd_sc_hd__a221o_1 _3913_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[14] ),
    .A2(_1396_),
    .B1(net425),
    .B2(_2110_),
    .C1(net411),
    .X(_1068_));
 sky130_fd_sc_hd__and3_1 _3914_ (.A(\device.configuration[15] ),
    .B(net629),
    .C(net626),
    .X(_2111_));
 sky130_fd_sc_hd__a221o_1 _3915_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[15] ),
    .A2(net508),
    .B1(net425),
    .B2(_2111_),
    .C1(net411),
    .X(_1069_));
 sky130_fd_sc_hd__and3_1 _3916_ (.A(\device.configuration[16] ),
    .B(net629),
    .C(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .X(_2112_));
 sky130_fd_sc_hd__a221o_1 _3917_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[16] ),
    .A2(net508),
    .B1(net425),
    .B2(_2112_),
    .C1(net411),
    .X(_1070_));
 sky130_fd_sc_hd__and3_1 _3918_ (.A(\device.configuration[17] ),
    .B(net630),
    .C(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .X(_2113_));
 sky130_fd_sc_hd__a221o_1 _3919_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[17] ),
    .A2(net508),
    .B1(net425),
    .B2(_2113_),
    .C1(net411),
    .X(_1071_));
 sky130_fd_sc_hd__and3_1 _3920_ (.A(\device.configuration[18] ),
    .B(net630),
    .C(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .X(_2114_));
 sky130_fd_sc_hd__a221o_1 _3921_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[18] ),
    .A2(net508),
    .B1(net425),
    .B2(_2114_),
    .C1(net411),
    .X(_1072_));
 sky130_fd_sc_hd__and3_1 _3922_ (.A(\device.configuration[19] ),
    .B(net629),
    .C(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .X(_2115_));
 sky130_fd_sc_hd__a221o_1 _3923_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[19] ),
    .A2(_1396_),
    .B1(net425),
    .B2(_2115_),
    .C1(_2104_),
    .X(_1073_));
 sky130_fd_sc_hd__and3_1 _3924_ (.A(\device.configuration[20] ),
    .B(net629),
    .C(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .X(_2116_));
 sky130_fd_sc_hd__a221o_1 _3925_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[20] ),
    .A2(_1396_),
    .B1(net426),
    .B2(_2116_),
    .C1(_2104_),
    .X(_1074_));
 sky130_fd_sc_hd__a21o_1 _3926_ (.A1(\wbPeripheralBusInterface.dataRead_buffered[21] ),
    .A2(net508),
    .B1(_2104_),
    .X(_1075_));
 sky130_fd_sc_hd__nor2_1 _3927_ (.A(net507),
    .B(_2064_),
    .Y(_2117_));
 sky130_fd_sc_hd__or4b_2 _3928_ (.A(_1342_),
    .B(_1343_),
    .C(_1393_),
    .D_N(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__o221a_1 _3929_ (.A1(net509),
    .A2(_2053_),
    .B1(_2118_),
    .B2(\wbPeripheralBusInterface.acknowledge ),
    .C1(net1954),
    .X(_1076_));
 sky130_fd_sc_hd__nand3_1 _3930_ (.A(net1580),
    .B(net486),
    .C(_1406_),
    .Y(_2119_));
 sky130_fd_sc_hd__or4b_2 _3931_ (.A(net645),
    .B(net446),
    .C(net1581),
    .D_N(net486),
    .X(_2120_));
 sky130_fd_sc_hd__mux2_1 _3932_ (.A0(net2848),
    .A1(\wbPeripheralBusInterface.currentAddress[2] ),
    .S(net422),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_1 _3933_ (.A0(net2860),
    .A1(\wbPeripheralBusInterface.currentAddress[3] ),
    .S(net422),
    .X(_1078_));
 sky130_fd_sc_hd__mux2_1 _3934_ (.A0(net2752),
    .A1(\wbPeripheralBusInterface.currentAddress[4] ),
    .S(net422),
    .X(_1079_));
 sky130_fd_sc_hd__mux2_1 _3935_ (.A0(net2764),
    .A1(\wbPeripheralBusInterface.currentAddress[5] ),
    .S(net422),
    .X(_1080_));
 sky130_fd_sc_hd__mux2_1 _3936_ (.A0(net2776),
    .A1(\wbPeripheralBusInterface.currentAddress[6] ),
    .S(net422),
    .X(_1081_));
 sky130_fd_sc_hd__mux2_1 _3937_ (.A0(net2788),
    .A1(\wbPeripheralBusInterface.currentAddress[7] ),
    .S(net422),
    .X(_1082_));
 sky130_fd_sc_hd__mux2_1 _3938_ (.A0(net2800),
    .A1(\wbPeripheralBusInterface.currentAddress[8] ),
    .S(net422),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _3939_ (.A0(net2812),
    .A1(\wbPeripheralBusInterface.currentAddress[9] ),
    .S(net422),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _3940_ (.A0(net2824),
    .A1(\wbPeripheralBusInterface.currentAddress[10] ),
    .S(net423),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_1 _3941_ (.A0(net2836),
    .A1(\wbPeripheralBusInterface.currentAddress[11] ),
    .S(net423),
    .X(_1086_));
 sky130_fd_sc_hd__mux2_1 _3942_ (.A0(net2872),
    .A1(\wbPeripheralBusInterface.currentAddress[12] ),
    .S(net423),
    .X(_1087_));
 sky130_fd_sc_hd__mux2_1 _3943_ (.A0(net2896),
    .A1(\wbPeripheralBusInterface.currentAddress[13] ),
    .S(net423),
    .X(_1088_));
 sky130_fd_sc_hd__mux2_1 _3944_ (.A0(net2884),
    .A1(\wbPeripheralBusInterface.currentAddress[14] ),
    .S(net423),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_1 _3945_ (.A0(\wbAddressExtension.currentAddress[15] ),
    .A1(\wbPeripheralBusInterface.currentAddress[15] ),
    .S(net423),
    .X(_1090_));
 sky130_fd_sc_hd__mux2_1 _3946_ (.A0(\wbAddressExtension.currentAddress[16] ),
    .A1(\wbPeripheralBusInterface.currentAddress[16] ),
    .S(net1602),
    .X(_1091_));
 sky130_fd_sc_hd__mux2_1 _3947_ (.A0(\wbAddressExtension.currentAddress[17] ),
    .A1(\wbPeripheralBusInterface.currentAddress[17] ),
    .S(net1602),
    .X(_1092_));
 sky130_fd_sc_hd__mux2_1 _3948_ (.A0(\wbAddressExtension.currentAddress[18] ),
    .A1(\wbPeripheralBusInterface.currentAddress[18] ),
    .S(net1602),
    .X(_1093_));
 sky130_fd_sc_hd__mux2_1 _3949_ (.A0(\wbAddressExtension.currentAddress[19] ),
    .A1(\wbPeripheralBusInterface.currentAddress[19] ),
    .S(net1602),
    .X(_1094_));
 sky130_fd_sc_hd__mux2_1 _3950_ (.A0(\wbAddressExtension.currentAddress[20] ),
    .A1(\wbPeripheralBusInterface.currentAddress[20] ),
    .S(net1602),
    .X(_1095_));
 sky130_fd_sc_hd__mux2_1 _3951_ (.A0(\wbAddressExtension.currentAddress[21] ),
    .A1(\wbPeripheralBusInterface.currentAddress[21] ),
    .S(net1602),
    .X(_1096_));
 sky130_fd_sc_hd__mux2_1 _3952_ (.A0(\wbAddressExtension.currentAddress[22] ),
    .A1(\wbPeripheralBusInterface.currentAddress[22] ),
    .S(net1602),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _3953_ (.A0(\wbAddressExtension.currentAddress[23] ),
    .A1(\wbPeripheralBusInterface.currentAddress[23] ),
    .S(net1602),
    .X(_1098_));
 sky130_fd_sc_hd__a21oi_1 _3954_ (.A1(net2329),
    .A2(net1282),
    .B1(net630),
    .Y(_2121_));
 sky130_fd_sc_hd__nor2_1 _3955_ (.A(net631),
    .B(net2403),
    .Y(_2122_));
 sky130_fd_sc_hd__a31o_1 _3956_ (.A1(net1580),
    .A2(net1282),
    .A3(_1976_),
    .B1(net559),
    .X(_2123_));
 sky130_fd_sc_hd__and2_1 _3957_ (.A(net632),
    .B(net3242),
    .X(_2124_));
 sky130_fd_sc_hd__o21a_1 _3958_ (.A1(net509),
    .A2(net2340),
    .B1(net3244),
    .X(_1099_));
 sky130_fd_sc_hd__or3_1 _3959_ (.A(net509),
    .B(_2053_),
    .C(net2403),
    .X(_2125_));
 sky130_fd_sc_hd__and3_1 _3960_ (.A(_2118_),
    .B(net3244),
    .C(net2405),
    .X(_1100_));
 sky130_fd_sc_hd__a21oi_1 _3961_ (.A1(net553),
    .A2(_2035_),
    .B1(net2731),
    .Y(_1101_));
 sky130_fd_sc_hd__nor2_4 _3962_ (.A(net1483),
    .B(_1496_),
    .Y(_0561_));
 sky130_fd_sc_hd__and2_1 _3963_ (.A(\device.rxBuffer.dataOut[0] ),
    .B(net1675),
    .X(_1190_));
 sky130_fd_sc_hd__and2_1 _3964_ (.A(\device.rxBuffer.dataOut[1] ),
    .B(net1675),
    .X(_1191_));
 sky130_fd_sc_hd__and2_1 _3965_ (.A(\device.rxBuffer.dataOut[2] ),
    .B(net1675),
    .X(_1192_));
 sky130_fd_sc_hd__and2_1 _3966_ (.A(\device.rxBuffer.dataOut[3] ),
    .B(net1675),
    .X(_1193_));
 sky130_fd_sc_hd__and2_1 _3967_ (.A(\device.rxBuffer.dataOut[4] ),
    .B(net1675),
    .X(_1194_));
 sky130_fd_sc_hd__and2_1 _3968_ (.A(\device.rxBuffer.dataOut[5] ),
    .B(net1675),
    .X(_1195_));
 sky130_fd_sc_hd__and2_1 _3969_ (.A(\device.rxBuffer.dataOut[6] ),
    .B(net1675),
    .X(_1196_));
 sky130_fd_sc_hd__and2_1 _3970_ (.A(\device.rxBuffer.dataOut[7] ),
    .B(net1675),
    .X(_1197_));
 sky130_fd_sc_hd__nand2_8 _3971_ (.A(net1440),
    .B(net1385),
    .Y(_2126_));
 sky130_fd_sc_hd__mux2_1 _3972_ (.A0(net198),
    .A1(\wbAddressExtension.currentAddress[8] ),
    .S(net1442),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _3973_ (.A0(net199),
    .A1(\wbAddressExtension.currentAddress[9] ),
    .S(net1442),
    .X(_1231_));
 sky130_fd_sc_hd__mux2_1 _3974_ (.A0(net169),
    .A1(\wbAddressExtension.currentAddress[10] ),
    .S(net1442),
    .X(_1232_));
 sky130_fd_sc_hd__mux2_1 _3975_ (.A0(net170),
    .A1(\wbAddressExtension.currentAddress[11] ),
    .S(net1442),
    .X(_1233_));
 sky130_fd_sc_hd__mux2_1 _3976_ (.A0(net171),
    .A1(\wbAddressExtension.currentAddress[12] ),
    .S(net1442),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_1 _3977_ (.A0(net172),
    .A1(\wbAddressExtension.currentAddress[13] ),
    .S(net1442),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_1 _3978_ (.A0(net173),
    .A1(\wbAddressExtension.currentAddress[14] ),
    .S(net1442),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_1 _3979_ (.A0(net174),
    .A1(\wbAddressExtension.currentAddress[15] ),
    .S(net1442),
    .X(_1237_));
 sky130_fd_sc_hd__nand2_8 _3980_ (.A(net1399),
    .B(net1385),
    .Y(_2127_));
 sky130_fd_sc_hd__mux2_1 _3981_ (.A0(net175),
    .A1(\wbAddressExtension.currentAddress[16] ),
    .S(net1401),
    .X(_1238_));
 sky130_fd_sc_hd__mux2_1 _3982_ (.A0(net176),
    .A1(\wbAddressExtension.currentAddress[17] ),
    .S(net1401),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_1 _3983_ (.A0(net177),
    .A1(\wbAddressExtension.currentAddress[18] ),
    .S(net1401),
    .X(_1240_));
 sky130_fd_sc_hd__mux2_1 _3984_ (.A0(net178),
    .A1(\wbAddressExtension.currentAddress[19] ),
    .S(net1401),
    .X(_1241_));
 sky130_fd_sc_hd__mux2_1 _3985_ (.A0(net180),
    .A1(\wbAddressExtension.currentAddress[20] ),
    .S(net1401),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _3986_ (.A0(net181),
    .A1(\wbAddressExtension.currentAddress[21] ),
    .S(net1401),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_1 _3987_ (.A0(net182),
    .A1(\wbAddressExtension.currentAddress[22] ),
    .S(net1401),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_1 _3988_ (.A0(net183),
    .A1(\wbAddressExtension.currentAddress[23] ),
    .S(net1401),
    .X(_1245_));
 sky130_fd_sc_hd__and2_4 _3989_ (.A(net1509),
    .B(net1385),
    .X(_2128_));
 sky130_fd_sc_hd__mux2_1 _3990_ (.A0(\wbAddressExtension.currentAddress[24] ),
    .A1(net184),
    .S(net1513),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_1 _3991_ (.A0(\wbAddressExtension.currentAddress[25] ),
    .A1(net185),
    .S(net1513),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _3992_ (.A0(\wbAddressExtension.currentAddress[26] ),
    .A1(net186),
    .S(net1513),
    .X(_1248_));
 sky130_fd_sc_hd__mux2_1 _3993_ (.A0(\wbAddressExtension.currentAddress[27] ),
    .A1(net187),
    .S(net1513),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_1 _3994_ (.A0(\wbAddressExtension.currentAddress[28] ),
    .A1(net188),
    .S(net1513),
    .X(_1250_));
 sky130_fd_sc_hd__mux2_1 _3995_ (.A0(\wbAddressExtension.currentAddress[29] ),
    .A1(net189),
    .S(net1513),
    .X(_1251_));
 sky130_fd_sc_hd__mux2_1 _3996_ (.A0(\wbAddressExtension.currentAddress[30] ),
    .A1(net191),
    .S(net1513),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_1 _3997_ (.A0(\wbAddressExtension.currentAddress[31] ),
    .A1(net192),
    .S(net1513),
    .X(_1253_));
 sky130_fd_sc_hd__mux2_1 _3998_ (.A0(net1378),
    .A1(net627),
    .S(net422),
    .X(_1278_));
 sky130_fd_sc_hd__mux2_1 _3999_ (.A0(net1440),
    .A1(net626),
    .S(net422),
    .X(_1279_));
 sky130_fd_sc_hd__mux2_1 _4000_ (.A0(net1399),
    .A1(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .S(net423),
    .X(_1280_));
 sky130_fd_sc_hd__a31oi_4 _4001_ (.A1(net168),
    .A2(net1282),
    .A3(net458),
    .B1(net1483),
    .Y(_2129_));
 sky130_fd_sc_hd__and2_2 _4002_ (.A(\device.uartRx.delayCounter[9] ),
    .B(\device.uartRx.delayCounter[8] ),
    .X(_2130_));
 sky130_fd_sc_hd__nand4_1 _4003_ (.A(\device.uartRx.delayCounter[11] ),
    .B(\device.uartRx.delayCounter[10] ),
    .C(\device.uartRx.delayCounter[9] ),
    .D(\device.uartRx.delayCounter[8] ),
    .Y(_2131_));
 sky130_fd_sc_hd__nand3_2 _4004_ (.A(\device.uartRx.delayCounter[2] ),
    .B(\device.uartRx.delayCounter[1] ),
    .C(\device.uartRx.delayCounter[0] ),
    .Y(_2132_));
 sky130_fd_sc_hd__and4_4 _4005_ (.A(\device.uartRx.delayCounter[3] ),
    .B(\device.uartRx.delayCounter[2] ),
    .C(\device.uartRx.delayCounter[1] ),
    .D(\device.uartRx.delayCounter[0] ),
    .X(_2133_));
 sky130_fd_sc_hd__nand4_4 _4006_ (.A(\device.uartRx.delayCounter[3] ),
    .B(\device.uartRx.delayCounter[2] ),
    .C(\device.uartRx.delayCounter[1] ),
    .D(\device.uartRx.delayCounter[0] ),
    .Y(_2134_));
 sky130_fd_sc_hd__and2_2 _4007_ (.A(\device.uartRx.delayCounter[5] ),
    .B(\device.uartRx.delayCounter[4] ),
    .X(_2135_));
 sky130_fd_sc_hd__nand2_2 _4008_ (.A(net552),
    .B(_2135_),
    .Y(_2136_));
 sky130_fd_sc_hd__and4_4 _4009_ (.A(\device.uartRx.delayCounter[7] ),
    .B(\device.uartRx.delayCounter[6] ),
    .C(\device.uartRx.delayCounter[5] ),
    .D(\device.uartRx.delayCounter[4] ),
    .X(_2137_));
 sky130_fd_sc_hd__nand2_1 _4010_ (.A(net552),
    .B(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__or3b_4 _4011_ (.A(_2131_),
    .B(_2134_),
    .C_N(_2137_),
    .X(_2139_));
 sky130_fd_sc_hd__and4bb_4 _4012_ (.A_N(_1348_),
    .B_N(_2131_),
    .C(net552),
    .D(_2137_),
    .X(_2140_));
 sky130_fd_sc_hd__or3b_4 _4013_ (.A(_1346_),
    .B(_1347_),
    .C_N(_2140_),
    .X(_2141_));
 sky130_fd_sc_hd__and4b_2 _4014_ (.A_N(\device.uartRx.delayCounter[15] ),
    .B(\device.uartRx.delayCounter[14] ),
    .C(\device.uartRx.delayCounter[13] ),
    .D(_2140_),
    .X(_2142_));
 sky130_fd_sc_hd__a21oi_4 _4015_ (.A1(\device.uartRx.delayCounter[15] ),
    .A2(_2141_),
    .B1(_2142_),
    .Y(_2143_));
 sky130_fd_sc_hd__xor2_2 _4016_ (.A(\device.configuration[15] ),
    .B(_2143_),
    .X(_2144_));
 sky130_fd_sc_hd__a21o_1 _4017_ (.A1(\device.uartRx.delayCounter[13] ),
    .A2(_2140_),
    .B1(\device.uartRx.delayCounter[14] ),
    .X(_2145_));
 sky130_fd_sc_hd__nand2_1 _4018_ (.A(_2141_),
    .B(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__a21oi_1 _4019_ (.A1(_2141_),
    .A2(_2145_),
    .B1(_1341_),
    .Y(_2147_));
 sky130_fd_sc_hd__and3_1 _4020_ (.A(_2130_),
    .B(net552),
    .C(_2137_),
    .X(_2148_));
 sky130_fd_sc_hd__nand4_4 _4021_ (.A(\device.uartRx.delayCounter[10] ),
    .B(_2130_),
    .C(_2133_),
    .D(_2137_),
    .Y(_2149_));
 sky130_fd_sc_hd__a21bo_2 _4022_ (.A1(_1349_),
    .A2(_2149_),
    .B1_N(_2139_),
    .X(_2150_));
 sky130_fd_sc_hd__xnor2_1 _4023_ (.A(\device.configuration[11] ),
    .B(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__and3_1 _4024_ (.A(_1341_),
    .B(_2141_),
    .C(_2145_),
    .X(_2152_));
 sky130_fd_sc_hd__or2_1 _4025_ (.A(_2147_),
    .B(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__or3_1 _4026_ (.A(_2147_),
    .B(_2151_),
    .C(_2152_),
    .X(_2154_));
 sky130_fd_sc_hd__xnor2_4 _4027_ (.A(_1348_),
    .B(_2139_),
    .Y(_2155_));
 sky130_fd_sc_hd__xor2_2 _4028_ (.A(\device.configuration[12] ),
    .B(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__and3_2 _4029_ (.A(\device.uartRx.delayCounter[8] ),
    .B(net552),
    .C(_2137_),
    .X(_2157_));
 sky130_fd_sc_hd__o21bai_4 _4030_ (.A1(\device.uartRx.delayCounter[9] ),
    .A2(_2157_),
    .B1_N(_2148_),
    .Y(_2158_));
 sky130_fd_sc_hd__xor2_4 _4031_ (.A(\device.configuration[9] ),
    .B(_2158_),
    .X(_2159_));
 sky130_fd_sc_hd__xnor2_4 _4032_ (.A(\device.uartRx.delayCounter[13] ),
    .B(_2140_),
    .Y(_2160_));
 sky130_fd_sc_hd__o211ai_4 _4033_ (.A1(\device.configuration[13] ),
    .A2(_2160_),
    .B1(_2159_),
    .C1(_2156_),
    .Y(_2161_));
 sky130_fd_sc_hd__or3b_2 _4034_ (.A(_1354_),
    .B(_2134_),
    .C_N(_2135_),
    .X(_2162_));
 sky130_fd_sc_hd__a31o_1 _4035_ (.A1(\device.uartRx.delayCounter[6] ),
    .A2(net552),
    .A3(_2135_),
    .B1(\device.uartRx.delayCounter[7] ),
    .X(_2163_));
 sky130_fd_sc_hd__nand2_1 _4036_ (.A(_2138_),
    .B(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__a21oi_1 _4037_ (.A1(_2138_),
    .A2(_2163_),
    .B1(_1340_),
    .Y(_2165_));
 sky130_fd_sc_hd__a21oi_1 _4038_ (.A1(net552),
    .A2(_2137_),
    .B1(\device.uartRx.delayCounter[8] ),
    .Y(_2166_));
 sky130_fd_sc_hd__or2_2 _4039_ (.A(_2157_),
    .B(_2166_),
    .X(_2167_));
 sky130_fd_sc_hd__o21a_1 _4040_ (.A1(_2157_),
    .A2(_2166_),
    .B1(\device.configuration[8] ),
    .X(_2168_));
 sky130_fd_sc_hd__nand3_1 _4041_ (.A(_1340_),
    .B(_2138_),
    .C(_2163_),
    .Y(_2169_));
 sky130_fd_sc_hd__or3b_1 _4042_ (.A(_2165_),
    .B(_2168_),
    .C_N(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__a21o_1 _4043_ (.A1(net552),
    .A2(_2135_),
    .B1(\device.uartRx.delayCounter[6] ),
    .X(_2171_));
 sky130_fd_sc_hd__nand2_1 _4044_ (.A(_2162_),
    .B(_2171_),
    .Y(_2172_));
 sky130_fd_sc_hd__a21bo_1 _4045_ (.A1(_2162_),
    .A2(_2171_),
    .B1_N(\device.configuration[6] ),
    .X(_2173_));
 sky130_fd_sc_hd__nand3b_1 _4046_ (.A_N(\device.configuration[6] ),
    .B(_2162_),
    .C(_2171_),
    .Y(_2174_));
 sky130_fd_sc_hd__a21o_2 _4047_ (.A1(\device.uartRx.delayCounter[4] ),
    .A2(net552),
    .B1(\device.uartRx.delayCounter[5] ),
    .X(_2175_));
 sky130_fd_sc_hd__nand2_1 _4048_ (.A(_2136_),
    .B(_2175_),
    .Y(_2176_));
 sky130_fd_sc_hd__a21oi_1 _4049_ (.A1(_2136_),
    .A2(_2175_),
    .B1(\device.configuration[5] ),
    .Y(_2177_));
 sky130_fd_sc_hd__and3_1 _4050_ (.A(\device.configuration[5] ),
    .B(_2136_),
    .C(_2175_),
    .X(_2178_));
 sky130_fd_sc_hd__o211a_1 _4051_ (.A1(_2177_),
    .A2(_2178_),
    .B1(_2173_),
    .C1(_2174_),
    .X(_2179_));
 sky130_fd_sc_hd__or3_1 _4052_ (.A(\device.configuration[8] ),
    .B(_2157_),
    .C(_2166_),
    .X(_2180_));
 sky130_fd_sc_hd__xnor2_1 _4053_ (.A(\device.configuration[1] ),
    .B(\device.uartRx.delayCounter[0] ),
    .Y(_2181_));
 sky130_fd_sc_hd__xnor2_4 _4054_ (.A(\device.uartRx.delayCounter[1] ),
    .B(\device.uartRx.delayCounter[0] ),
    .Y(_2182_));
 sky130_fd_sc_hd__xor2_1 _4055_ (.A(\device.configuration[1] ),
    .B(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__xor2_1 _4056_ (.A(\device.configuration[0] ),
    .B(\device.uartRx.delayCounter[0] ),
    .X(_2184_));
 sky130_fd_sc_hd__a21o_1 _4057_ (.A1(\device.uartRx.delayCounter[1] ),
    .A2(\device.uartRx.delayCounter[0] ),
    .B1(\device.uartRx.delayCounter[2] ),
    .X(_2185_));
 sky130_fd_sc_hd__nand2_1 _4058_ (.A(_2132_),
    .B(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hd__and3_1 _4059_ (.A(\device.configuration[2] ),
    .B(_2132_),
    .C(_2185_),
    .X(_2187_));
 sky130_fd_sc_hd__a21oi_1 _4060_ (.A1(_2132_),
    .A2(_2185_),
    .B1(\device.configuration[2] ),
    .Y(_2188_));
 sky130_fd_sc_hd__o211a_1 _4061_ (.A1(_2187_),
    .A2(_2188_),
    .B1(_2183_),
    .C1(_2184_),
    .X(_2189_));
 sky130_fd_sc_hd__a31o_1 _4062_ (.A1(\device.uartRx.delayCounter[2] ),
    .A2(\device.uartRx.delayCounter[1] ),
    .A3(\device.uartRx.delayCounter[0] ),
    .B1(\device.uartRx.delayCounter[3] ),
    .X(_2190_));
 sky130_fd_sc_hd__nand2_2 _4063_ (.A(_2134_),
    .B(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__xor2_2 _4064_ (.A(\device.configuration[3] ),
    .B(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__xnor2_4 _4065_ (.A(\device.uartRx.delayCounter[4] ),
    .B(net552),
    .Y(_2193_));
 sky130_fd_sc_hd__xor2_2 _4066_ (.A(\device.configuration[4] ),
    .B(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__and4_1 _4067_ (.A(_2180_),
    .B(_2189_),
    .C(_2192_),
    .D(_2194_),
    .X(_2195_));
 sky130_fd_sc_hd__a31o_1 _4068_ (.A1(_2130_),
    .A2(_2133_),
    .A3(_2137_),
    .B1(\device.uartRx.delayCounter[10] ),
    .X(_2196_));
 sky130_fd_sc_hd__nand2_1 _4069_ (.A(_2149_),
    .B(_2196_),
    .Y(_2197_));
 sky130_fd_sc_hd__a21oi_1 _4070_ (.A1(_2149_),
    .A2(_2196_),
    .B1(\device.configuration[10] ),
    .Y(_2198_));
 sky130_fd_sc_hd__and3_1 _4071_ (.A(\device.configuration[10] ),
    .B(_2149_),
    .C(_2196_),
    .X(_2199_));
 sky130_fd_sc_hd__o2bb2a_1 _4072_ (.A1_N(\device.configuration[13] ),
    .A2_N(_2160_),
    .B1(_2198_),
    .B2(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__and4b_1 _4073_ (.A_N(_2170_),
    .B(_2179_),
    .C(_2195_),
    .D(_2200_),
    .X(_2201_));
 sky130_fd_sc_hd__and4bb_1 _4074_ (.A_N(_2154_),
    .B_N(_2161_),
    .C(_2201_),
    .D(_2144_),
    .X(_2202_));
 sky130_fd_sc_hd__or4bb_4 _4075_ (.A(_2154_),
    .B(_2161_),
    .C_N(_2201_),
    .D_N(_2144_),
    .X(_2203_));
 sky130_fd_sc_hd__and2b_1 _4076_ (.A_N(\device.uartRx.state[0] ),
    .B(\device.uartRx.state[1] ),
    .X(_2204_));
 sky130_fd_sc_hd__nand2b_4 _4077_ (.A_N(\device.uartRx.state[0] ),
    .B(\device.uartRx.state[1] ),
    .Y(_2205_));
 sky130_fd_sc_hd__nor2_4 _4078_ (.A(_2203_),
    .B(_2205_),
    .Y(_2206_));
 sky130_fd_sc_hd__nand2_1 _4079_ (.A(\device.uartRx.bitCounter[1] ),
    .B(\device.uartRx.bitCounter[0] ),
    .Y(_2207_));
 sky130_fd_sc_hd__nor2_1 _4080_ (.A(_1344_),
    .B(_2207_),
    .Y(_2208_));
 sky130_fd_sc_hd__and3_2 _4081_ (.A(_2202_),
    .B(_2204_),
    .C(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__and2_1 _4082_ (.A(net420),
    .B(_2209_),
    .X(_1297_));
 sky130_fd_sc_hd__and2_1 _4083_ (.A(\device.uartRx.savedData[0] ),
    .B(net439),
    .X(_1306_));
 sky130_fd_sc_hd__and2_1 _4084_ (.A(\device.uartRx.savedData[1] ),
    .B(net439),
    .X(_1307_));
 sky130_fd_sc_hd__and2_1 _4085_ (.A(\device.uartRx.savedData[2] ),
    .B(net439),
    .X(_1308_));
 sky130_fd_sc_hd__and2_1 _4086_ (.A(\device.uartRx.savedData[3] ),
    .B(net439),
    .X(_1309_));
 sky130_fd_sc_hd__and2_1 _4087_ (.A(\device.uartRx.savedData[4] ),
    .B(net439),
    .X(_1310_));
 sky130_fd_sc_hd__and2_1 _4088_ (.A(\device.uartRx.savedData[5] ),
    .B(net439),
    .X(_1311_));
 sky130_fd_sc_hd__and2_1 _4089_ (.A(\device.uartRx.savedData[6] ),
    .B(_1442_),
    .X(_1312_));
 sky130_fd_sc_hd__and2_1 _4090_ (.A(\device.uartRx.savedData[7] ),
    .B(_1442_),
    .X(_1313_));
 sky130_fd_sc_hd__and2_4 _4091_ (.A(_1419_),
    .B(_2117_),
    .X(_2210_));
 sky130_fd_sc_hd__o2111a_1 _4092_ (.A1(_1342_),
    .A2(_1393_),
    .B1(net559),
    .C1(_2210_),
    .D1(net628),
    .X(_1333_));
 sky130_fd_sc_hd__and4b_1 _4093_ (.A_N(\device.txSendBusy ),
    .B(net440),
    .C(_1722_),
    .D(\device.configuration[17] ),
    .X(_1334_));
 sky130_fd_sc_hd__and3_1 _4094_ (.A(\device.configuration[17] ),
    .B(\device.uartRx.newData ),
    .C(_1442_),
    .X(_0581_));
 sky130_fd_sc_hd__and2_1 _4095_ (.A(net3447),
    .B(_2066_),
    .X(_0582_));
 sky130_fd_sc_hd__and2_1 _4096_ (.A(\device.uartTx.bitCounter[1] ),
    .B(\device.uartTx.bitCounter[0] ),
    .X(_2211_));
 sky130_fd_sc_hd__and3_1 _4097_ (.A(\device.uartTx.bitCounter[2] ),
    .B(\device.uartTx.state[1] ),
    .C(_2211_),
    .X(_2212_));
 sky130_fd_sc_hd__nand3_4 _4098_ (.A(\device.uartTx.delayCounter[2] ),
    .B(\device.uartTx.delayCounter[1] ),
    .C(\device.uartTx.delayCounter[0] ),
    .Y(_2213_));
 sky130_fd_sc_hd__and4_2 _4099_ (.A(\device.uartTx.delayCounter[3] ),
    .B(\device.uartTx.delayCounter[2] ),
    .C(\device.uartTx.delayCounter[1] ),
    .D(\device.uartTx.delayCounter[0] ),
    .X(_2214_));
 sky130_fd_sc_hd__and4_4 _4100_ (.A(\device.uartTx.delayCounter[7] ),
    .B(\device.uartTx.delayCounter[6] ),
    .C(\device.uartTx.delayCounter[5] ),
    .D(\device.uartTx.delayCounter[4] ),
    .X(_2215_));
 sky130_fd_sc_hd__nand2_1 _4101_ (.A(net550),
    .B(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__and2_2 _4102_ (.A(\device.uartTx.delayCounter[9] ),
    .B(\device.uartTx.delayCounter[8] ),
    .X(_2217_));
 sky130_fd_sc_hd__and4_2 _4103_ (.A(\device.uartTx.delayCounter[11] ),
    .B(\device.uartTx.delayCounter[10] ),
    .C(\device.uartTx.delayCounter[9] ),
    .D(\device.uartTx.delayCounter[8] ),
    .X(_2218_));
 sky130_fd_sc_hd__and4_4 _4104_ (.A(\device.uartTx.delayCounter[12] ),
    .B(net551),
    .C(_2215_),
    .D(_2218_),
    .X(_2219_));
 sky130_fd_sc_hd__nand3_4 _4105_ (.A(\device.uartTx.delayCounter[14] ),
    .B(\device.uartTx.delayCounter[13] ),
    .C(_2219_),
    .Y(_2220_));
 sky130_fd_sc_hd__xor2_2 _4106_ (.A(\device.uartTx.delayCounter[15] ),
    .B(_2220_),
    .X(_2221_));
 sky130_fd_sc_hd__xor2_1 _4107_ (.A(\device.configuration[15] ),
    .B(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__nand4_4 _4108_ (.A(\device.uartTx.delayCounter[10] ),
    .B(net551),
    .C(_2215_),
    .D(_2217_),
    .Y(_2223_));
 sky130_fd_sc_hd__a32o_1 _4109_ (.A1(net550),
    .A2(_2215_),
    .A3(_2218_),
    .B1(_2223_),
    .B2(_1362_),
    .X(_2224_));
 sky130_fd_sc_hd__xor2_1 _4110_ (.A(\device.configuration[11] ),
    .B(_2224_),
    .X(_2225_));
 sky130_fd_sc_hd__a31o_1 _4111_ (.A1(net551),
    .A2(_2215_),
    .A3(_2217_),
    .B1(\device.uartTx.delayCounter[10] ),
    .X(_2226_));
 sky130_fd_sc_hd__nand2_1 _4112_ (.A(_2223_),
    .B(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__a21bo_1 _4113_ (.A1(_2223_),
    .A2(_2226_),
    .B1_N(\device.configuration[10] ),
    .X(_2228_));
 sky130_fd_sc_hd__nand3b_1 _4114_ (.A_N(\device.configuration[10] ),
    .B(_2223_),
    .C(_2226_),
    .Y(_2229_));
 sky130_fd_sc_hd__a31oi_4 _4115_ (.A1(net551),
    .A2(_2215_),
    .A3(_2218_),
    .B1(\device.uartTx.delayCounter[12] ),
    .Y(_2230_));
 sky130_fd_sc_hd__or3_1 _4116_ (.A(\device.configuration[12] ),
    .B(_2219_),
    .C(_2230_),
    .X(_2231_));
 sky130_fd_sc_hd__o21ai_1 _4117_ (.A1(_2219_),
    .A2(_2230_),
    .B1(\device.configuration[12] ),
    .Y(_2232_));
 sky130_fd_sc_hd__and4_1 _4118_ (.A(_2228_),
    .B(_2229_),
    .C(_2231_),
    .D(_2232_),
    .X(_2233_));
 sky130_fd_sc_hd__nand3_2 _4119_ (.A(\device.uartTx.delayCounter[8] ),
    .B(net550),
    .C(_2215_),
    .Y(_2234_));
 sky130_fd_sc_hd__a21o_1 _4120_ (.A1(net550),
    .A2(_2215_),
    .B1(\device.uartTx.delayCounter[8] ),
    .X(_2235_));
 sky130_fd_sc_hd__nand2_1 _4121_ (.A(_2234_),
    .B(_2235_),
    .Y(_2236_));
 sky130_fd_sc_hd__and3_1 _4122_ (.A(\device.configuration[8] ),
    .B(_2234_),
    .C(_2235_),
    .X(_2237_));
 sky130_fd_sc_hd__a21oi_2 _4123_ (.A1(_2234_),
    .A2(_2235_),
    .B1(\device.configuration[8] ),
    .Y(_2238_));
 sky130_fd_sc_hd__nand3_1 _4124_ (.A(\device.uartTx.delayCounter[5] ),
    .B(\device.uartTx.delayCounter[4] ),
    .C(net550),
    .Y(_2239_));
 sky130_fd_sc_hd__nand4_2 _4125_ (.A(\device.uartTx.delayCounter[6] ),
    .B(\device.uartTx.delayCounter[5] ),
    .C(\device.uartTx.delayCounter[4] ),
    .D(net550),
    .Y(_2240_));
 sky130_fd_sc_hd__a31o_1 _4126_ (.A1(\device.uartTx.delayCounter[5] ),
    .A2(\device.uartTx.delayCounter[4] ),
    .A3(net550),
    .B1(\device.uartTx.delayCounter[6] ),
    .X(_2241_));
 sky130_fd_sc_hd__nand2_1 _4127_ (.A(_2240_),
    .B(_2241_),
    .Y(_2242_));
 sky130_fd_sc_hd__nand3b_1 _4128_ (.A_N(\device.configuration[6] ),
    .B(_2240_),
    .C(_2241_),
    .Y(_2243_));
 sky130_fd_sc_hd__a21o_1 _4129_ (.A1(\device.uartTx.delayCounter[4] ),
    .A2(net550),
    .B1(\device.uartTx.delayCounter[5] ),
    .X(_2244_));
 sky130_fd_sc_hd__nand2_1 _4130_ (.A(_2239_),
    .B(_2244_),
    .Y(_2245_));
 sky130_fd_sc_hd__o221a_1 _4131_ (.A1(_2237_),
    .A2(_2238_),
    .B1(_2245_),
    .B2(\device.configuration[5] ),
    .C1(_2243_),
    .X(_2246_));
 sky130_fd_sc_hd__xnor2_2 _4132_ (.A(\device.uartTx.delayCounter[4] ),
    .B(net550),
    .Y(_2247_));
 sky130_fd_sc_hd__xor2_1 _4133_ (.A(\device.configuration[4] ),
    .B(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__xor2_2 _4134_ (.A(\device.uartTx.delayCounter[3] ),
    .B(_2213_),
    .X(_2249_));
 sky130_fd_sc_hd__xor2_1 _4135_ (.A(\device.configuration[3] ),
    .B(_2249_),
    .X(_2250_));
 sky130_fd_sc_hd__xor2_4 _4136_ (.A(\device.uartTx.delayCounter[1] ),
    .B(\device.uartTx.delayCounter[0] ),
    .X(_2251_));
 sky130_fd_sc_hd__xnor2_1 _4137_ (.A(\device.configuration[1] ),
    .B(_2251_),
    .Y(_2252_));
 sky130_fd_sc_hd__nand2_1 _4138_ (.A(\device.configuration[0] ),
    .B(\device.uartTx.delayCounter[0] ),
    .Y(_2253_));
 sky130_fd_sc_hd__or2_1 _4139_ (.A(\device.configuration[0] ),
    .B(\device.uartTx.delayCounter[0] ),
    .X(_2254_));
 sky130_fd_sc_hd__a21o_1 _4140_ (.A1(\device.uartTx.delayCounter[1] ),
    .A2(\device.uartTx.delayCounter[0] ),
    .B1(\device.uartTx.delayCounter[2] ),
    .X(_2255_));
 sky130_fd_sc_hd__nand2_1 _4141_ (.A(_2213_),
    .B(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__and3_1 _4142_ (.A(\device.configuration[2] ),
    .B(_2213_),
    .C(_2255_),
    .X(_2257_));
 sky130_fd_sc_hd__a21oi_1 _4143_ (.A1(_2213_),
    .A2(_2255_),
    .B1(\device.configuration[2] ),
    .Y(_2258_));
 sky130_fd_sc_hd__o2111a_1 _4144_ (.A1(_2257_),
    .A2(_2258_),
    .B1(_2252_),
    .C1(_2253_),
    .D1(_2254_),
    .X(_2259_));
 sky130_fd_sc_hd__and3_1 _4145_ (.A(_2248_),
    .B(_2250_),
    .C(_2259_),
    .X(_2260_));
 sky130_fd_sc_hd__a21bo_1 _4146_ (.A1(_2239_),
    .A2(_2244_),
    .B1_N(\device.configuration[5] ),
    .X(_2261_));
 sky130_fd_sc_hd__a21bo_1 _4147_ (.A1(_2240_),
    .A2(_2241_),
    .B1_N(\device.configuration[6] ),
    .X(_2262_));
 sky130_fd_sc_hd__and2_1 _4148_ (.A(_2261_),
    .B(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__and4_1 _4149_ (.A(_2233_),
    .B(_2246_),
    .C(_2260_),
    .D(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__a21o_1 _4150_ (.A1(\device.uartTx.delayCounter[13] ),
    .A2(_2219_),
    .B1(\device.uartTx.delayCounter[14] ),
    .X(_2265_));
 sky130_fd_sc_hd__nand2_1 _4151_ (.A(_2220_),
    .B(_2265_),
    .Y(_2266_));
 sky130_fd_sc_hd__a21oi_2 _4152_ (.A1(_2220_),
    .A2(_2265_),
    .B1(\device.configuration[14] ),
    .Y(_2267_));
 sky130_fd_sc_hd__and3_1 _4153_ (.A(\device.configuration[14] ),
    .B(_2220_),
    .C(_2265_),
    .X(_2268_));
 sky130_fd_sc_hd__xnor2_2 _4154_ (.A(\device.uartTx.delayCounter[13] ),
    .B(_2219_),
    .Y(_2269_));
 sky130_fd_sc_hd__xor2_1 _4155_ (.A(\device.configuration[13] ),
    .B(_2269_),
    .X(_2270_));
 sky130_fd_sc_hd__a32o_2 _4156_ (.A1(net551),
    .A2(_2215_),
    .A3(_2217_),
    .B1(_2234_),
    .B2(_1363_),
    .X(_2271_));
 sky130_fd_sc_hd__xor2_1 _4157_ (.A(\device.configuration[9] ),
    .B(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__a41o_1 _4158_ (.A1(\device.uartTx.delayCounter[6] ),
    .A2(\device.uartTx.delayCounter[5] ),
    .A3(\device.uartTx.delayCounter[4] ),
    .A4(net550),
    .B1(\device.uartTx.delayCounter[7] ),
    .X(_2273_));
 sky130_fd_sc_hd__nand2_1 _4159_ (.A(_2216_),
    .B(_2273_),
    .Y(_2274_));
 sky130_fd_sc_hd__xnor2_1 _4160_ (.A(_1340_),
    .B(_2274_),
    .Y(_2275_));
 sky130_fd_sc_hd__o2111a_1 _4161_ (.A1(_2267_),
    .A2(_2268_),
    .B1(_2270_),
    .C1(_2272_),
    .D1(_2275_),
    .X(_2276_));
 sky130_fd_sc_hd__and4_4 _4162_ (.A(_2222_),
    .B(_2225_),
    .C(_2264_),
    .D(_2276_),
    .X(_2277_));
 sky130_fd_sc_hd__nand2_8 _4163_ (.A(\device.configuration[17] ),
    .B(_2050_),
    .Y(_2278_));
 sky130_fd_sc_hd__nor2_4 _4164_ (.A(net418),
    .B(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__nor2_1 _4165_ (.A(\device.uartTx.state[0] ),
    .B(_2212_),
    .Y(_2280_));
 sky130_fd_sc_hd__a21o_1 _4166_ (.A1(_2216_),
    .A2(_2273_),
    .B1(_1340_),
    .X(_2281_));
 sky130_fd_sc_hd__nand3_1 _4167_ (.A(_1340_),
    .B(_2216_),
    .C(_2273_),
    .Y(_2282_));
 sky130_fd_sc_hd__o221a_1 _4168_ (.A1(_2237_),
    .A2(_2238_),
    .B1(_2271_),
    .B2(\device.configuration[9] ),
    .C1(_2231_),
    .X(_2283_));
 sky130_fd_sc_hd__and4_1 _4169_ (.A(_2228_),
    .B(_2232_),
    .C(_2281_),
    .D(_2282_),
    .X(_2284_));
 sky130_fd_sc_hd__and4_1 _4170_ (.A(_2225_),
    .B(_2270_),
    .C(_2283_),
    .D(_2284_),
    .X(_2285_));
 sky130_fd_sc_hd__and3_1 _4171_ (.A(_2243_),
    .B(_2250_),
    .C(_2261_),
    .X(_2286_));
 sky130_fd_sc_hd__o2111a_1 _4172_ (.A1(\device.configuration[5] ),
    .A2(_2245_),
    .B1(_2248_),
    .C1(_2259_),
    .D1(_2262_),
    .X(_2287_));
 sky130_fd_sc_hd__a21boi_1 _4173_ (.A1(\device.configuration[9] ),
    .A2(_2271_),
    .B1_N(_2229_),
    .Y(_2288_));
 sky130_fd_sc_hd__o2111a_1 _4174_ (.A1(_2267_),
    .A2(_2268_),
    .B1(_2286_),
    .C1(_2287_),
    .D1(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__a211o_1 _4175_ (.A1(_2212_),
    .A2(_2277_),
    .B1(_2279_),
    .C1(\device.uartTx.state[0] ),
    .X(_2290_));
 sky130_fd_sc_hd__nand2_1 _4176_ (.A(\device.uartTx.state[0] ),
    .B(_2277_),
    .Y(_2291_));
 sky130_fd_sc_hd__and4_1 _4177_ (.A(\device.uartTx.state[0] ),
    .B(_2222_),
    .C(_2285_),
    .D(_2289_),
    .X(_2292_));
 sky130_fd_sc_hd__and3_1 _4178_ (.A(net2023),
    .B(_2290_),
    .C(_2291_),
    .X(_0727_));
 sky130_fd_sc_hd__a31o_1 _4179_ (.A1(\device.uartTx.state[1] ),
    .A2(\device.uartTx.state[0] ),
    .A3(_2277_),
    .B1(net427),
    .X(_2293_));
 sky130_fd_sc_hd__a21oi_1 _4180_ (.A1(_1364_),
    .A2(_2291_),
    .B1(_2293_),
    .Y(_0728_));
 sky130_fd_sc_hd__nor2_1 _4181_ (.A(\device.configuration[17] ),
    .B(_2051_),
    .Y(_2294_));
 sky130_fd_sc_hd__a21o_1 _4182_ (.A1(\device.uartTx.state[1] ),
    .A2(_2292_),
    .B1(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__nor2_1 _4183_ (.A(\device.uartTx.delayCounter[0] ),
    .B(_2050_),
    .Y(_2296_));
 sky130_fd_sc_hd__nor2_2 _4184_ (.A(_2277_),
    .B(_2294_),
    .Y(_2297_));
 sky130_fd_sc_hd__o221a_1 _4185_ (.A1(net409),
    .A2(_2296_),
    .B1(_2297_),
    .B2(\device.uartTx.delayCounter[0] ),
    .C1(net2023),
    .X(_0737_));
 sky130_fd_sc_hd__or2_2 _4186_ (.A(_2050_),
    .B(_2277_),
    .X(_2298_));
 sky130_fd_sc_hd__a32oi_4 _4187_ (.A1(_2051_),
    .A2(_2251_),
    .A3(_2297_),
    .B1(net409),
    .B2(\device.uartTx.delayCounter[1] ),
    .Y(_2299_));
 sky130_fd_sc_hd__nor2_1 _4188_ (.A(net427),
    .B(_2299_),
    .Y(_0738_));
 sky130_fd_sc_hd__o2bb2a_1 _4189_ (.A1_N(\device.uartTx.delayCounter[2] ),
    .A2_N(net409),
    .B1(net408),
    .B2(_2256_),
    .X(_2300_));
 sky130_fd_sc_hd__nor2_1 _4190_ (.A(net1984),
    .B(_2300_),
    .Y(_0739_));
 sky130_fd_sc_hd__o2bb2a_1 _4191_ (.A1_N(\device.uartTx.delayCounter[3] ),
    .A2_N(net409),
    .B1(net408),
    .B2(_2249_),
    .X(_2301_));
 sky130_fd_sc_hd__nor2_1 _4192_ (.A(net1984),
    .B(_2301_),
    .Y(_0740_));
 sky130_fd_sc_hd__o2bb2a_1 _4193_ (.A1_N(\device.uartTx.delayCounter[4] ),
    .A2_N(net409),
    .B1(net408),
    .B2(_2247_),
    .X(_2302_));
 sky130_fd_sc_hd__nor2_1 _4194_ (.A(net1984),
    .B(_2302_),
    .Y(_0741_));
 sky130_fd_sc_hd__o2bb2a_1 _4195_ (.A1_N(\device.uartTx.delayCounter[5] ),
    .A2_N(net409),
    .B1(net408),
    .B2(_2245_),
    .X(_2303_));
 sky130_fd_sc_hd__nor2_1 _4196_ (.A(net1984),
    .B(_2303_),
    .Y(_0742_));
 sky130_fd_sc_hd__o2bb2a_1 _4197_ (.A1_N(\device.uartTx.delayCounter[6] ),
    .A2_N(net409),
    .B1(net408),
    .B2(_2242_),
    .X(_2304_));
 sky130_fd_sc_hd__nor2_1 _4198_ (.A(net1984),
    .B(_2304_),
    .Y(_0743_));
 sky130_fd_sc_hd__o2bb2a_1 _4199_ (.A1_N(\device.uartTx.delayCounter[7] ),
    .A2_N(net409),
    .B1(net408),
    .B2(_2274_),
    .X(_2305_));
 sky130_fd_sc_hd__nor2_1 _4200_ (.A(net1984),
    .B(_2305_),
    .Y(_0744_));
 sky130_fd_sc_hd__o2bb2a_1 _4201_ (.A1_N(\device.uartTx.delayCounter[8] ),
    .A2_N(net409),
    .B1(net408),
    .B2(_2236_),
    .X(_2306_));
 sky130_fd_sc_hd__nor2_1 _4202_ (.A(net1984),
    .B(_2306_),
    .Y(_0745_));
 sky130_fd_sc_hd__o2bb2a_1 _4203_ (.A1_N(\device.uartTx.delayCounter[9] ),
    .A2_N(net409),
    .B1(_2298_),
    .B2(_2271_),
    .X(_2307_));
 sky130_fd_sc_hd__nor2_1 _4204_ (.A(net1984),
    .B(_2307_),
    .Y(_0746_));
 sky130_fd_sc_hd__o2bb2a_1 _4205_ (.A1_N(\device.uartTx.delayCounter[10] ),
    .A2_N(net410),
    .B1(_2298_),
    .B2(_2227_),
    .X(_2308_));
 sky130_fd_sc_hd__nor2_1 _4206_ (.A(net427),
    .B(_2308_),
    .Y(_0747_));
 sky130_fd_sc_hd__o2bb2a_1 _4207_ (.A1_N(\device.uartTx.delayCounter[11] ),
    .A2_N(net410),
    .B1(_2298_),
    .B2(_2224_),
    .X(_2309_));
 sky130_fd_sc_hd__nor2_1 _4208_ (.A(net427),
    .B(_2309_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_1 _4209_ (.A(\device.uartTx.delayCounter[12] ),
    .B(net410),
    .Y(_2310_));
 sky130_fd_sc_hd__or3_1 _4210_ (.A(_2219_),
    .B(_2230_),
    .C(net408),
    .X(_2311_));
 sky130_fd_sc_hd__a21oi_1 _4211_ (.A1(_2310_),
    .A2(_2311_),
    .B1(net427),
    .Y(_0749_));
 sky130_fd_sc_hd__o2bb2a_1 _4212_ (.A1_N(\device.uartTx.delayCounter[13] ),
    .A2_N(net410),
    .B1(net408),
    .B2(_2269_),
    .X(_2312_));
 sky130_fd_sc_hd__nor2_1 _4213_ (.A(net427),
    .B(_2312_),
    .Y(_0750_));
 sky130_fd_sc_hd__o2bb2a_1 _4214_ (.A1_N(\device.uartTx.delayCounter[14] ),
    .A2_N(net410),
    .B1(net408),
    .B2(_2266_),
    .X(_2313_));
 sky130_fd_sc_hd__nor2_1 _4215_ (.A(net427),
    .B(_2313_),
    .Y(_0751_));
 sky130_fd_sc_hd__o2bb2a_1 _4216_ (.A1_N(\device.uartTx.delayCounter[15] ),
    .A2_N(net410),
    .B1(_2298_),
    .B2(_2221_),
    .X(_2314_));
 sky130_fd_sc_hd__nor2_1 _4217_ (.A(net427),
    .B(_2314_),
    .Y(_0752_));
 sky130_fd_sc_hd__o221a_2 _4218_ (.A1(\device.configuration[17] ),
    .A2(_2051_),
    .B1(_2277_),
    .B2(_1364_),
    .C1(_2280_),
    .X(_2315_));
 sky130_fd_sc_hd__a31o_1 _4219_ (.A1(\device.uartTx.state[1] ),
    .A2(_2277_),
    .A3(_2280_),
    .B1(\device.uartTx.bitCounter[0] ),
    .X(_2316_));
 sky130_fd_sc_hd__nand2_1 _4220_ (.A(\device.uartTx.bitCounter[0] ),
    .B(_2315_),
    .Y(_2317_));
 sky130_fd_sc_hd__and3_1 _4221_ (.A(net2023),
    .B(_2316_),
    .C(_2317_),
    .X(_0753_));
 sky130_fd_sc_hd__or2_1 _4222_ (.A(_2049_),
    .B(_2211_),
    .X(_2318_));
 sky130_fd_sc_hd__a21o_1 _4223_ (.A1(_2315_),
    .A2(_2318_),
    .B1(net427),
    .X(_2319_));
 sky130_fd_sc_hd__a21oi_1 _4224_ (.A1(_1361_),
    .A2(_2317_),
    .B1(_2319_),
    .Y(_0754_));
 sky130_fd_sc_hd__a21bo_1 _4225_ (.A1(_2315_),
    .A2(_2318_),
    .B1_N(\device.uartTx.bitCounter[2] ),
    .X(_2320_));
 sky130_fd_sc_hd__or4bb_1 _4226_ (.A(\device.uartTx.bitCounter[2] ),
    .B(_2049_),
    .C_N(_2211_),
    .D_N(_2315_),
    .X(_2321_));
 sky130_fd_sc_hd__a21oi_1 _4227_ (.A1(_2320_),
    .A2(_2321_),
    .B1(net427),
    .Y(_0755_));
 sky130_fd_sc_hd__or2_1 _4228_ (.A(\device.uartTx.savedData[0] ),
    .B(_2279_),
    .X(_2322_));
 sky130_fd_sc_hd__o311a_1 _4229_ (.A1(\device.txBuffer.dataOut[0] ),
    .A2(net418),
    .A3(_2278_),
    .B1(_2322_),
    .C1(net2023),
    .X(_0756_));
 sky130_fd_sc_hd__or2_1 _4230_ (.A(\device.uartTx.savedData[1] ),
    .B(_2279_),
    .X(_2323_));
 sky130_fd_sc_hd__o311a_1 _4231_ (.A1(\device.txBuffer.dataOut[1] ),
    .A2(net418),
    .A3(_2278_),
    .B1(_2323_),
    .C1(net2023),
    .X(_0757_));
 sky130_fd_sc_hd__or2_1 _4232_ (.A(\device.uartTx.savedData[2] ),
    .B(_2279_),
    .X(_2324_));
 sky130_fd_sc_hd__o311a_1 _4233_ (.A1(\device.txBuffer.dataOut[2] ),
    .A2(net418),
    .A3(_2278_),
    .B1(_2324_),
    .C1(net2023),
    .X(_0758_));
 sky130_fd_sc_hd__or2_1 _4234_ (.A(\device.uartTx.savedData[3] ),
    .B(_2279_),
    .X(_2325_));
 sky130_fd_sc_hd__o311a_1 _4235_ (.A1(\device.txBuffer.dataOut[3] ),
    .A2(net418),
    .A3(_2278_),
    .B1(_2325_),
    .C1(net2023),
    .X(_0759_));
 sky130_fd_sc_hd__or2_1 _4236_ (.A(\device.uartTx.savedData[4] ),
    .B(_2279_),
    .X(_2326_));
 sky130_fd_sc_hd__o311a_1 _4237_ (.A1(\device.txBuffer.dataOut[4] ),
    .A2(net418),
    .A3(_2278_),
    .B1(_2326_),
    .C1(net2023),
    .X(_0760_));
 sky130_fd_sc_hd__or2_1 _4238_ (.A(\device.uartTx.savedData[5] ),
    .B(_2279_),
    .X(_2327_));
 sky130_fd_sc_hd__o311a_1 _4239_ (.A1(\device.txBuffer.dataOut[5] ),
    .A2(_1723_),
    .A3(_2278_),
    .B1(_2327_),
    .C1(net2023),
    .X(_0761_));
 sky130_fd_sc_hd__or2_1 _4240_ (.A(\device.uartTx.savedData[6] ),
    .B(_2279_),
    .X(_2328_));
 sky130_fd_sc_hd__o311a_1 _4241_ (.A1(\device.txBuffer.dataOut[6] ),
    .A2(_1723_),
    .A3(_2278_),
    .B1(_2328_),
    .C1(net2022),
    .X(_0762_));
 sky130_fd_sc_hd__or2_1 _4242_ (.A(\device.uartTx.savedData[7] ),
    .B(_2279_),
    .X(_2329_));
 sky130_fd_sc_hd__o311a_1 _4243_ (.A1(\device.txBuffer.dataOut[7] ),
    .A2(_1723_),
    .A3(_2278_),
    .B1(_2329_),
    .C1(net2022),
    .X(_0763_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(\device.txSendBusy ),
    .A1(_2278_),
    .S(net2023),
    .X(_0764_));
 sky130_fd_sc_hd__nand2b_1 _4245_ (.A_N(\device.uartRx.state[1] ),
    .B(\device.uartRx.state[0] ),
    .Y(_2330_));
 sky130_fd_sc_hd__a21oi_1 _4246_ (.A1(_2141_),
    .A2(_2145_),
    .B1(\device.configuration[15] ),
    .Y(_2331_));
 sky130_fd_sc_hd__and3_1 _4247_ (.A(\device.configuration[15] ),
    .B(_2141_),
    .C(_2145_),
    .X(_2332_));
 sky130_fd_sc_hd__xor2_1 _4248_ (.A(\device.configuration[11] ),
    .B(_2197_),
    .X(_2333_));
 sky130_fd_sc_hd__xor2_1 _4249_ (.A(\device.configuration[10] ),
    .B(_2158_),
    .X(_2334_));
 sky130_fd_sc_hd__o2111a_1 _4250_ (.A1(_2331_),
    .A2(_2332_),
    .B1(_2333_),
    .C1(_2334_),
    .D1(_2143_),
    .X(_2335_));
 sky130_fd_sc_hd__a22o_1 _4251_ (.A1(\device.configuration[12] ),
    .A2(_2150_),
    .B1(_2160_),
    .B2(\device.configuration[14] ),
    .X(_2336_));
 sky130_fd_sc_hd__o21ba_1 _4252_ (.A1(\device.configuration[14] ),
    .A2(_2160_),
    .B1_N(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__xnor2_1 _4253_ (.A(_1340_),
    .B(_2172_),
    .Y(_2338_));
 sky130_fd_sc_hd__and3_1 _4254_ (.A(\device.configuration[6] ),
    .B(_2136_),
    .C(_2175_),
    .X(_2339_));
 sky130_fd_sc_hd__a21oi_1 _4255_ (.A1(_2136_),
    .A2(_2175_),
    .B1(\device.configuration[6] ),
    .Y(_2340_));
 sky130_fd_sc_hd__o22a_1 _4256_ (.A1(\device.configuration[9] ),
    .A2(_2167_),
    .B1(_2339_),
    .B2(_2340_),
    .X(_2341_));
 sky130_fd_sc_hd__a21boi_1 _4257_ (.A1(_2132_),
    .A2(_2185_),
    .B1_N(\device.configuration[3] ),
    .Y(_2342_));
 sky130_fd_sc_hd__xnor2_1 _4258_ (.A(\device.configuration[2] ),
    .B(_2182_),
    .Y(_2343_));
 sky130_fd_sc_hd__and3b_1 _4259_ (.A_N(\device.configuration[3] ),
    .B(_2132_),
    .C(_2185_),
    .X(_2344_));
 sky130_fd_sc_hd__or4_1 _4260_ (.A(_2181_),
    .B(_2342_),
    .C(_2343_),
    .D(_2344_),
    .X(_2345_));
 sky130_fd_sc_hd__xnor2_1 _4261_ (.A(\device.configuration[4] ),
    .B(_2191_),
    .Y(_2346_));
 sky130_fd_sc_hd__xnor2_1 _4262_ (.A(\device.configuration[5] ),
    .B(_2193_),
    .Y(_2347_));
 sky130_fd_sc_hd__a2111o_1 _4263_ (.A1(\device.configuration[9] ),
    .A2(_2167_),
    .B1(_2345_),
    .C1(_2346_),
    .D1(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__xor2_1 _4264_ (.A(\device.configuration[8] ),
    .B(_2164_),
    .X(_2349_));
 sky130_fd_sc_hd__and4b_1 _4265_ (.A_N(_2348_),
    .B(_2338_),
    .C(_2341_),
    .D(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__xor2_1 _4266_ (.A(\device.configuration[13] ),
    .B(_2155_),
    .X(_2351_));
 sky130_fd_sc_hd__o21a_1 _4267_ (.A1(\device.configuration[12] ),
    .A2(_2150_),
    .B1(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__and4_2 _4268_ (.A(_2335_),
    .B(_2337_),
    .C(_2350_),
    .D(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__nor2_1 _4269_ (.A(_2330_),
    .B(_2353_),
    .Y(_2354_));
 sky130_fd_sc_hd__xnor2_1 _4270_ (.A(\device.configuration[13] ),
    .B(_2160_),
    .Y(_2355_));
 sky130_fd_sc_hd__nand4_1 _4271_ (.A(_2173_),
    .B(_2174_),
    .C(_2189_),
    .D(_2194_),
    .Y(_2356_));
 sky130_fd_sc_hd__a211o_1 _4272_ (.A1(\device.configuration[12] ),
    .A2(_2155_),
    .B1(_2165_),
    .C1(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__o221a_1 _4273_ (.A1(\device.configuration[12] ),
    .A2(_2155_),
    .B1(_2177_),
    .B2(_2178_),
    .C1(_2169_),
    .X(_2358_));
 sky130_fd_sc_hd__or3b_1 _4274_ (.A(_2151_),
    .B(_2355_),
    .C_N(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__and3b_1 _4275_ (.A_N(_2168_),
    .B(_2180_),
    .C(_2192_),
    .X(_2360_));
 sky130_fd_sc_hd__o211a_1 _4276_ (.A1(_2198_),
    .A2(_2199_),
    .B1(_2360_),
    .C1(_2159_),
    .X(_2361_));
 sky130_fd_sc_hd__or4b_2 _4277_ (.A(_2153_),
    .B(_2357_),
    .C(_2359_),
    .D_N(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__o22a_2 _4278_ (.A1(_2202_),
    .A2(_2205_),
    .B1(_2330_),
    .B2(_2353_),
    .X(_2363_));
 sky130_fd_sc_hd__or2_1 _4279_ (.A(_2205_),
    .B(_2208_),
    .X(_2364_));
 sky130_fd_sc_hd__nor2_1 _4280_ (.A(_1343_),
    .B(net1),
    .Y(_2365_));
 sky130_fd_sc_hd__or2_1 _4281_ (.A(_1343_),
    .B(net1),
    .X(_2366_));
 sky130_fd_sc_hd__nand2_2 _4282_ (.A(\device.uartRx.state[1] ),
    .B(\device.uartRx.state[0] ),
    .Y(_2367_));
 sky130_fd_sc_hd__or3_1 _4283_ (.A(\device.uartRx.state[1] ),
    .B(\device.uartRx.state[0] ),
    .C(_2365_),
    .X(_2368_));
 sky130_fd_sc_hd__o211a_1 _4284_ (.A1(_2366_),
    .A2(net549),
    .B1(_2368_),
    .C1(_2364_),
    .X(_2369_));
 sky130_fd_sc_hd__a21o_1 _4285_ (.A1(net407),
    .A2(_2369_),
    .B1(\device.uartRx.state[0] ),
    .X(_2370_));
 sky130_fd_sc_hd__nand2_1 _4286_ (.A(\device.uartRx.state[0] ),
    .B(_2369_),
    .Y(_2371_));
 sky130_fd_sc_hd__o211a_1 _4287_ (.A1(_2354_),
    .A2(_2371_),
    .B1(_2370_),
    .C1(net420),
    .X(_0861_));
 sky130_fd_sc_hd__a21o_1 _4288_ (.A1(\device.uartRx.state[0] ),
    .A2(_2353_),
    .B1(\device.uartRx.state[1] ),
    .X(_2372_));
 sky130_fd_sc_hd__o211a_1 _4289_ (.A1(_2365_),
    .A2(net549),
    .B1(_2372_),
    .C1(net420),
    .X(_0862_));
 sky130_fd_sc_hd__a21bo_1 _4290_ (.A1(\device.uartRx.delayCounter[0] ),
    .A2(net548),
    .B1_N(net419),
    .X(_2373_));
 sky130_fd_sc_hd__a21oi_1 _4291_ (.A1(_1360_),
    .A2(net406),
    .B1(_2373_),
    .Y(_0863_));
 sky130_fd_sc_hd__o22a_1 _4292_ (.A1(_2182_),
    .A2(net406),
    .B1(net548),
    .B2(_1359_),
    .X(_2374_));
 sky130_fd_sc_hd__and2b_1 _4293_ (.A_N(_2374_),
    .B(net419),
    .X(_0864_));
 sky130_fd_sc_hd__o22a_1 _4294_ (.A1(_2186_),
    .A2(net406),
    .B1(net548),
    .B2(_1358_),
    .X(_2375_));
 sky130_fd_sc_hd__and2b_1 _4295_ (.A_N(_2375_),
    .B(net419),
    .X(_0865_));
 sky130_fd_sc_hd__o22a_1 _4296_ (.A1(_2191_),
    .A2(net406),
    .B1(net548),
    .B2(_1357_),
    .X(_2376_));
 sky130_fd_sc_hd__and2b_1 _4297_ (.A_N(_2376_),
    .B(net419),
    .X(_0866_));
 sky130_fd_sc_hd__o22a_1 _4298_ (.A1(_2193_),
    .A2(net406),
    .B1(net548),
    .B2(_1356_),
    .X(_2377_));
 sky130_fd_sc_hd__and2b_1 _4299_ (.A_N(_2377_),
    .B(net419),
    .X(_0867_));
 sky130_fd_sc_hd__o22a_1 _4300_ (.A1(_2176_),
    .A2(net406),
    .B1(net548),
    .B2(_1355_),
    .X(_2378_));
 sky130_fd_sc_hd__and2b_1 _4301_ (.A_N(_2378_),
    .B(net419),
    .X(_0868_));
 sky130_fd_sc_hd__o22a_1 _4302_ (.A1(_2172_),
    .A2(net406),
    .B1(net548),
    .B2(_1354_),
    .X(_2379_));
 sky130_fd_sc_hd__and2b_1 _4303_ (.A_N(_2379_),
    .B(net419),
    .X(_0869_));
 sky130_fd_sc_hd__o22a_1 _4304_ (.A1(_2164_),
    .A2(net406),
    .B1(net548),
    .B2(_1353_),
    .X(_2380_));
 sky130_fd_sc_hd__and2b_1 _4305_ (.A_N(_2380_),
    .B(net419),
    .X(_0870_));
 sky130_fd_sc_hd__o22a_1 _4306_ (.A1(_2167_),
    .A2(net406),
    .B1(net548),
    .B2(_1352_),
    .X(_2381_));
 sky130_fd_sc_hd__and2b_1 _4307_ (.A_N(_2381_),
    .B(net419),
    .X(_0871_));
 sky130_fd_sc_hd__o22a_1 _4308_ (.A1(_2158_),
    .A2(net406),
    .B1(net548),
    .B2(_1351_),
    .X(_2382_));
 sky130_fd_sc_hd__and2b_1 _4309_ (.A_N(_2382_),
    .B(net419),
    .X(_0872_));
 sky130_fd_sc_hd__o22a_1 _4310_ (.A1(_2197_),
    .A2(net407),
    .B1(net549),
    .B2(_1350_),
    .X(_2383_));
 sky130_fd_sc_hd__and2b_1 _4311_ (.A_N(_2383_),
    .B(net1764),
    .X(_0873_));
 sky130_fd_sc_hd__o22a_1 _4312_ (.A1(_2150_),
    .A2(net407),
    .B1(net549),
    .B2(_1349_),
    .X(_2384_));
 sky130_fd_sc_hd__and2b_1 _4313_ (.A_N(_2384_),
    .B(net1787),
    .X(_0874_));
 sky130_fd_sc_hd__o22a_1 _4314_ (.A1(_2155_),
    .A2(net407),
    .B1(net549),
    .B2(_1348_),
    .X(_2385_));
 sky130_fd_sc_hd__and2b_1 _4315_ (.A_N(_2385_),
    .B(net1787),
    .X(_0875_));
 sky130_fd_sc_hd__o22a_1 _4316_ (.A1(_2160_),
    .A2(net407),
    .B1(net549),
    .B2(_1347_),
    .X(_2386_));
 sky130_fd_sc_hd__and2b_1 _4317_ (.A_N(_2386_),
    .B(net1764),
    .X(_0876_));
 sky130_fd_sc_hd__o22a_1 _4318_ (.A1(_2146_),
    .A2(net407),
    .B1(net549),
    .B2(_1346_),
    .X(_2387_));
 sky130_fd_sc_hd__and2b_1 _4319_ (.A_N(_2387_),
    .B(net1764),
    .X(_0877_));
 sky130_fd_sc_hd__and3_1 _4320_ (.A(\device.uartRx.delayCounter[15] ),
    .B(\device.uartRx.state[1] ),
    .C(\device.uartRx.state[0] ),
    .X(_2388_));
 sky130_fd_sc_hd__a21o_2 _4321_ (.A1(\device.uartRx.state[1] ),
    .A2(_2203_),
    .B1(\device.uartRx.state[0] ),
    .X(_2389_));
 sky130_fd_sc_hd__and3b_1 _4322_ (.A_N(_2143_),
    .B(net549),
    .C(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__o21a_1 _4323_ (.A1(_2388_),
    .A2(_2390_),
    .B1(net1764),
    .X(_0878_));
 sky130_fd_sc_hd__or3b_4 _4324_ (.A(_2205_),
    .B(_2362_),
    .C_N(_2144_),
    .X(_2391_));
 sky130_fd_sc_hd__nor2_1 _4325_ (.A(_2209_),
    .B(_2389_),
    .Y(_2392_));
 sky130_fd_sc_hd__a211o_1 _4326_ (.A1(_1345_),
    .A2(\device.uartRx.state[1] ),
    .B1(_2209_),
    .C1(_2389_),
    .X(_2393_));
 sky130_fd_sc_hd__o211a_1 _4327_ (.A1(\device.uartRx.bitCounter[0] ),
    .A2(_2392_),
    .B1(_2393_),
    .C1(net1764),
    .X(_0879_));
 sky130_fd_sc_hd__or2_1 _4328_ (.A(\device.uartRx.bitCounter[1] ),
    .B(\device.uartRx.bitCounter[0] ),
    .X(_2394_));
 sky130_fd_sc_hd__a311o_1 _4329_ (.A1(_2204_),
    .A2(_2207_),
    .A3(_2394_),
    .B1(_2389_),
    .C1(_2209_),
    .X(_2395_));
 sky130_fd_sc_hd__o211a_1 _4330_ (.A1(\device.uartRx.bitCounter[1] ),
    .A2(_2392_),
    .B1(_2395_),
    .C1(net1764),
    .X(_0880_));
 sky130_fd_sc_hd__a21o_1 _4331_ (.A1(_1344_),
    .A2(_2207_),
    .B1(_2364_),
    .X(_2396_));
 sky130_fd_sc_hd__a21bo_1 _4332_ (.A1(_1344_),
    .A2(_2389_),
    .B1_N(net420),
    .X(_2397_));
 sky130_fd_sc_hd__a21oi_1 _4333_ (.A1(_2392_),
    .A2(_2396_),
    .B1(_2397_),
    .Y(_0881_));
 sky130_fd_sc_hd__or2_1 _4334_ (.A(\device.uartRx.savedData[0] ),
    .B(_2206_),
    .X(_2398_));
 sky130_fd_sc_hd__o211a_1 _4335_ (.A1(\device.uartRx.savedData[1] ),
    .A2(_2391_),
    .B1(_2398_),
    .C1(net420),
    .X(_0882_));
 sky130_fd_sc_hd__or2_1 _4336_ (.A(\device.uartRx.savedData[1] ),
    .B(_2206_),
    .X(_2399_));
 sky130_fd_sc_hd__o211a_1 _4337_ (.A1(\device.uartRx.savedData[2] ),
    .A2(_2391_),
    .B1(_2399_),
    .C1(net420),
    .X(_0883_));
 sky130_fd_sc_hd__or2_1 _4338_ (.A(\device.uartRx.savedData[2] ),
    .B(_2206_),
    .X(_2400_));
 sky130_fd_sc_hd__o211a_1 _4339_ (.A1(\device.uartRx.savedData[3] ),
    .A2(_2391_),
    .B1(_2400_),
    .C1(net420),
    .X(_0884_));
 sky130_fd_sc_hd__or2_1 _4340_ (.A(\device.uartRx.savedData[3] ),
    .B(_2206_),
    .X(_2401_));
 sky130_fd_sc_hd__o211a_1 _4341_ (.A1(\device.uartRx.savedData[4] ),
    .A2(_2391_),
    .B1(_2401_),
    .C1(net420),
    .X(_0885_));
 sky130_fd_sc_hd__or2_1 _4342_ (.A(\device.uartRx.savedData[4] ),
    .B(_2206_),
    .X(_2402_));
 sky130_fd_sc_hd__o211a_1 _4343_ (.A1(\device.uartRx.savedData[5] ),
    .A2(_2391_),
    .B1(_2402_),
    .C1(net420),
    .X(_0886_));
 sky130_fd_sc_hd__or2_1 _4344_ (.A(\device.uartRx.savedData[5] ),
    .B(_2206_),
    .X(_2403_));
 sky130_fd_sc_hd__o211a_1 _4345_ (.A1(\device.uartRx.savedData[6] ),
    .A2(_2391_),
    .B1(_2403_),
    .C1(net1764),
    .X(_0887_));
 sky130_fd_sc_hd__or2_1 _4346_ (.A(\device.uartRx.savedData[6] ),
    .B(_2206_),
    .X(_2404_));
 sky130_fd_sc_hd__o211a_1 _4347_ (.A1(\device.uartRx.savedData[7] ),
    .A2(_2391_),
    .B1(_2404_),
    .C1(net1764),
    .X(_0888_));
 sky130_fd_sc_hd__or2_1 _4348_ (.A(\device.uartRx.savedData[7] ),
    .B(_2206_),
    .X(_2405_));
 sky130_fd_sc_hd__o211a_1 _4349_ (.A1(_2366_),
    .A2(_2391_),
    .B1(_2405_),
    .C1(net420),
    .X(_0889_));
 sky130_fd_sc_hd__and3_1 _4350_ (.A(net168),
    .B(net1286),
    .C(_2210_),
    .X(_0890_));
 sky130_fd_sc_hd__and4_1 _4351_ (.A(net2924),
    .B(net179),
    .C(net502),
    .D(_2210_),
    .X(_0891_));
 sky130_fd_sc_hd__and3_1 _4352_ (.A(net190),
    .B(net1286),
    .C(_2210_),
    .X(_0892_));
 sky130_fd_sc_hd__and3_1 _4353_ (.A(net193),
    .B(net1286),
    .C(_2210_),
    .X(_0893_));
 sky130_fd_sc_hd__and3_1 _4354_ (.A(net194),
    .B(net1286),
    .C(_2210_),
    .X(_0894_));
 sky130_fd_sc_hd__and3_1 _4355_ (.A(net195),
    .B(net1286),
    .C(_2210_),
    .X(_0895_));
 sky130_fd_sc_hd__and3_1 _4356_ (.A(net196),
    .B(net1971),
    .C(_2210_),
    .X(_0896_));
 sky130_fd_sc_hd__and3_1 _4357_ (.A(net197),
    .B(net1971),
    .C(_2210_),
    .X(_0897_));
 sky130_fd_sc_hd__nor2_2 _4358_ (.A(net4150),
    .B(_1457_),
    .Y(_0922_));
 sky130_fd_sc_hd__and2_1 _4359_ (.A(\device.rxBuffer.lastWriteLostData ),
    .B(net1992),
    .X(_0923_));
 sky130_fd_sc_hd__nor2_1 _4360_ (.A(net1466),
    .B(net418),
    .Y(_0924_));
 sky130_fd_sc_hd__nor2_1 _4361_ (.A(net3863),
    .B(_1393_),
    .Y(_0925_));
 sky130_fd_sc_hd__and2_1 _4362_ (.A(\device.txBuffer.lastWriteLostData ),
    .B(net632),
    .X(_0926_));
 sky130_fd_sc_hd__and2_1 _4363_ (.A(net632),
    .B(\device.rxDataAvailableBuffered ),
    .X(_0927_));
 sky130_fd_sc_hd__and2_1 _4364_ (.A(net1992),
    .B(\device.rxBufferFullBuffered ),
    .X(_0928_));
 sky130_fd_sc_hd__and2_1 _4365_ (.A(net1992),
    .B(\device.rxDataLostBuffered ),
    .X(_0929_));
 sky130_fd_sc_hd__and2_1 _4366_ (.A(net632),
    .B(\device.txDataAvailableBuffered ),
    .X(_0930_));
 sky130_fd_sc_hd__and2_1 _4367_ (.A(net632),
    .B(\device.txBufferFullBuffered ),
    .X(_0931_));
 sky130_fd_sc_hd__and2_1 _4368_ (.A(net632),
    .B(\device.txDataLostBuffered ),
    .X(_0932_));
 sky130_fd_sc_hd__nor4_2 _4369_ (.A(_1397_),
    .B(_1410_),
    .C(_1418_),
    .D(_2060_),
    .Y(_2406_));
 sky130_fd_sc_hd__and2_4 _4370_ (.A(\wbPeripheralBusInterface.currentByteSelect[2] ),
    .B(net460),
    .X(_2407_));
 sky130_fd_sc_hd__a21bo_1 _4371_ (.A1(net180),
    .A2(net488),
    .B1_N(_2407_),
    .X(_2408_));
 sky130_fd_sc_hd__o211a_1 _4372_ (.A1(\device.configuration[20] ),
    .A2(_2407_),
    .B1(net3104),
    .C1(net634),
    .X(_0933_));
 sky130_fd_sc_hd__a21bo_1 _4373_ (.A1(net178),
    .A2(net488),
    .B1_N(_2407_),
    .X(_2409_));
 sky130_fd_sc_hd__o211a_1 _4374_ (.A1(\device.configuration[19] ),
    .A2(_2407_),
    .B1(net3232),
    .C1(net634),
    .X(_0934_));
 sky130_fd_sc_hd__a21bo_1 _4375_ (.A1(net177),
    .A2(net488),
    .B1_N(_2407_),
    .X(_2410_));
 sky130_fd_sc_hd__o211a_1 _4376_ (.A1(\device.configuration[18] ),
    .A2(_2407_),
    .B1(net3210),
    .C1(net2156),
    .X(_0935_));
 sky130_fd_sc_hd__a21bo_1 _4377_ (.A1(net176),
    .A2(net487),
    .B1_N(_2407_),
    .X(_2411_));
 sky130_fd_sc_hd__o211a_1 _4378_ (.A1(\device.configuration[17] ),
    .A2(_2407_),
    .B1(net3127),
    .C1(net634),
    .X(_0936_));
 sky130_fd_sc_hd__a21bo_1 _4379_ (.A1(net175),
    .A2(net488),
    .B1_N(_2407_),
    .X(_2412_));
 sky130_fd_sc_hd__o211a_1 _4380_ (.A1(\device.configuration[16] ),
    .A2(_2407_),
    .B1(net3155),
    .C1(net2156),
    .X(_0937_));
 sky130_fd_sc_hd__and2_1 _4381_ (.A(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .B(net460),
    .X(_2413_));
 sky130_fd_sc_hd__a21bo_1 _4382_ (.A1(net174),
    .A2(net487),
    .B1_N(net444),
    .X(_2414_));
 sky130_fd_sc_hd__o211a_1 _4383_ (.A1(\device.configuration[15] ),
    .A2(net445),
    .B1(net3221),
    .C1(net634),
    .X(_0938_));
 sky130_fd_sc_hd__a21bo_1 _4384_ (.A1(net173),
    .A2(net487),
    .B1_N(net444),
    .X(_2415_));
 sky130_fd_sc_hd__o211a_1 _4385_ (.A1(\device.configuration[14] ),
    .A2(net445),
    .B1(net3199),
    .C1(net634),
    .X(_0939_));
 sky130_fd_sc_hd__a21bo_1 _4386_ (.A1(net172),
    .A2(net487),
    .B1_N(net445),
    .X(_2416_));
 sky130_fd_sc_hd__o211a_1 _4387_ (.A1(\device.configuration[13] ),
    .A2(net445),
    .B1(net3177),
    .C1(net634),
    .X(_0940_));
 sky130_fd_sc_hd__and2b_1 _4388_ (.A_N(net445),
    .B(\device.configuration[12] ),
    .X(_2417_));
 sky130_fd_sc_hd__and3_1 _4389_ (.A(net171),
    .B(net487),
    .C(net445),
    .X(_2418_));
 sky130_fd_sc_hd__or3_1 _4390_ (.A(net1483),
    .B(_2417_),
    .C(net2585),
    .X(_0941_));
 sky130_fd_sc_hd__a21bo_1 _4391_ (.A1(net170),
    .A2(net487),
    .B1_N(net444),
    .X(_2419_));
 sky130_fd_sc_hd__o211a_1 _4392_ (.A1(\device.configuration[11] ),
    .A2(net444),
    .B1(net3188),
    .C1(net634),
    .X(_0942_));
 sky130_fd_sc_hd__a21bo_1 _4393_ (.A1(net169),
    .A2(net487),
    .B1_N(net444),
    .X(_2420_));
 sky130_fd_sc_hd__o211a_1 _4394_ (.A1(\device.configuration[10] ),
    .A2(net444),
    .B1(net3166),
    .C1(net634),
    .X(_0943_));
 sky130_fd_sc_hd__a21bo_1 _4395_ (.A1(net199),
    .A2(net1971),
    .B1_N(net444),
    .X(_2421_));
 sky130_fd_sc_hd__o211a_1 _4396_ (.A1(\device.configuration[9] ),
    .A2(net444),
    .B1(_2421_),
    .C1(net634),
    .X(_0944_));
 sky130_fd_sc_hd__a21bo_1 _4397_ (.A1(net198),
    .A2(net1971),
    .B1_N(net444),
    .X(_2422_));
 sky130_fd_sc_hd__o211a_1 _4398_ (.A1(\device.configuration[8] ),
    .A2(net444),
    .B1(_2422_),
    .C1(net1954),
    .X(_0945_));
 sky130_fd_sc_hd__nor4_2 _4399_ (.A(_1375_),
    .B(net507),
    .C(_1410_),
    .D(_2055_),
    .Y(_2423_));
 sky130_fd_sc_hd__a21bo_1 _4400_ (.A1(net197),
    .A2(net1971),
    .B1_N(net443),
    .X(_2424_));
 sky130_fd_sc_hd__nand2_2 _4401_ (.A(net628),
    .B(_2406_),
    .Y(_2425_));
 sky130_fd_sc_hd__o211a_1 _4402_ (.A1(\device.configuration[7] ),
    .A2(net443),
    .B1(net1972),
    .C1(net1954),
    .X(_0946_));
 sky130_fd_sc_hd__a31o_1 _4403_ (.A1(net196),
    .A2(net1971),
    .A3(net443),
    .B1(net2731),
    .X(_2426_));
 sky130_fd_sc_hd__a21o_1 _4404_ (.A1(\device.configuration[6] ),
    .A2(_2425_),
    .B1(net1750),
    .X(_0947_));
 sky130_fd_sc_hd__a21bo_1 _4405_ (.A1(net195),
    .A2(net484),
    .B1_N(net443),
    .X(_2427_));
 sky130_fd_sc_hd__o211a_1 _4406_ (.A1(\device.configuration[5] ),
    .A2(net443),
    .B1(_2427_),
    .C1(net632),
    .X(_0948_));
 sky130_fd_sc_hd__a21bo_1 _4407_ (.A1(net194),
    .A2(net484),
    .B1_N(net443),
    .X(_2428_));
 sky130_fd_sc_hd__o211a_1 _4408_ (.A1(\device.configuration[4] ),
    .A2(net443),
    .B1(_2428_),
    .C1(net632),
    .X(_0949_));
 sky130_fd_sc_hd__or2_1 _4409_ (.A(\device.configuration[3] ),
    .B(_2423_),
    .X(_2429_));
 sky130_fd_sc_hd__o211a_1 _4410_ (.A1(net4170),
    .A2(_2425_),
    .B1(_2429_),
    .C1(net632),
    .X(_0950_));
 sky130_fd_sc_hd__a31o_1 _4411_ (.A1(net190),
    .A2(net484),
    .A3(net443),
    .B1(net1734),
    .X(_2430_));
 sky130_fd_sc_hd__a21o_1 _4412_ (.A1(\device.configuration[2] ),
    .A2(_2425_),
    .B1(_2430_),
    .X(_0951_));
 sky130_fd_sc_hd__a41o_1 _4413_ (.A1(net2924),
    .A2(net179),
    .A3(net502),
    .A4(net443),
    .B1(net1734),
    .X(_2431_));
 sky130_fd_sc_hd__a21o_1 _4414_ (.A1(\device.configuration[1] ),
    .A2(_2425_),
    .B1(net2928),
    .X(_0952_));
 sky130_fd_sc_hd__a31o_1 _4415_ (.A1(net168),
    .A2(net484),
    .A3(net443),
    .B1(net1734),
    .X(_2432_));
 sky130_fd_sc_hd__a21o_1 _4416_ (.A1(\device.configuration[0] ),
    .A2(_2425_),
    .B1(_2432_),
    .X(_0953_));
 sky130_fd_sc_hd__inv_2 _4417__2 (.A(clknet_leaf_31_wb_clk_i),
    .Y(net733));
 sky130_fd_sc_hd__inv_2 _4418__3 (.A(clknet_leaf_31_wb_clk_i),
    .Y(net734));
 sky130_fd_sc_hd__inv_2 _4419__4 (.A(clknet_leaf_35_wb_clk_i),
    .Y(net735));
 sky130_fd_sc_hd__inv_2 _4420__5 (.A(clknet_leaf_30_wb_clk_i),
    .Y(net736));
 sky130_fd_sc_hd__inv_2 _4421__6 (.A(clknet_leaf_29_wb_clk_i),
    .Y(net737));
 sky130_fd_sc_hd__inv_2 _4422__7 (.A(clknet_leaf_28_wb_clk_i),
    .Y(net738));
 sky130_fd_sc_hd__inv_2 _4423__8 (.A(clknet_leaf_30_wb_clk_i),
    .Y(net739));
 sky130_fd_sc_hd__inv_2 _4424__9 (.A(clknet_leaf_39_wb_clk_i),
    .Y(net740));
 sky130_fd_sc_hd__inv_2 _4425__10 (.A(clknet_leaf_43_wb_clk_i),
    .Y(net741));
 sky130_fd_sc_hd__inv_2 _4426__11 (.A(clknet_leaf_51_wb_clk_i),
    .Y(net742));
 sky130_fd_sc_hd__inv_2 _4427__12 (.A(clknet_leaf_51_wb_clk_i),
    .Y(net743));
 sky130_fd_sc_hd__inv_2 _4428__13 (.A(clknet_leaf_40_wb_clk_i),
    .Y(net744));
 sky130_fd_sc_hd__inv_2 _4429__14 (.A(clknet_leaf_39_wb_clk_i),
    .Y(net745));
 sky130_fd_sc_hd__inv_2 _4430__15 (.A(clknet_leaf_52_wb_clk_i),
    .Y(net746));
 sky130_fd_sc_hd__inv_2 _4431__16 (.A(clknet_leaf_51_wb_clk_i),
    .Y(net747));
 sky130_fd_sc_hd__inv_2 _4432__17 (.A(clknet_leaf_41_wb_clk_i),
    .Y(net748));
 sky130_fd_sc_hd__inv_2 _4433__18 (.A(clknet_leaf_24_wb_clk_i),
    .Y(net749));
 sky130_fd_sc_hd__inv_2 _4434__19 (.A(clknet_leaf_23_wb_clk_i),
    .Y(net750));
 sky130_fd_sc_hd__inv_2 _4435__20 (.A(clknet_leaf_15_wb_clk_i),
    .Y(net751));
 sky130_fd_sc_hd__inv_2 _4436__21 (.A(clknet_leaf_18_wb_clk_i),
    .Y(net752));
 sky130_fd_sc_hd__inv_2 _4437__22 (.A(clknet_leaf_19_wb_clk_i),
    .Y(net753));
 sky130_fd_sc_hd__inv_2 _4438__23 (.A(clknet_leaf_20_wb_clk_i),
    .Y(net754));
 sky130_fd_sc_hd__inv_2 _4439__24 (.A(clknet_leaf_23_wb_clk_i),
    .Y(net755));
 sky130_fd_sc_hd__inv_2 _4440__25 (.A(clknet_leaf_39_wb_clk_i),
    .Y(net756));
 sky130_fd_sc_hd__inv_2 _4441__26 (.A(clknet_leaf_47_wb_clk_i),
    .Y(net757));
 sky130_fd_sc_hd__inv_2 _4442__27 (.A(clknet_leaf_47_wb_clk_i),
    .Y(net758));
 sky130_fd_sc_hd__inv_2 _4443__28 (.A(clknet_leaf_47_wb_clk_i),
    .Y(net759));
 sky130_fd_sc_hd__inv_2 _4444__29 (.A(clknet_leaf_38_wb_clk_i),
    .Y(net760));
 sky130_fd_sc_hd__inv_2 _4445__30 (.A(clknet_leaf_38_wb_clk_i),
    .Y(net761));
 sky130_fd_sc_hd__inv_2 _4446__31 (.A(clknet_leaf_52_wb_clk_i),
    .Y(net762));
 sky130_fd_sc_hd__inv_2 _4447__32 (.A(clknet_leaf_50_wb_clk_i),
    .Y(net763));
 sky130_fd_sc_hd__inv_2 _4448__33 (.A(clknet_leaf_87_wb_clk_i),
    .Y(net764));
 sky130_fd_sc_hd__inv_2 _4449__34 (.A(clknet_leaf_87_wb_clk_i),
    .Y(net765));
 sky130_fd_sc_hd__inv_2 _4450__35 (.A(clknet_leaf_86_wb_clk_i),
    .Y(net766));
 sky130_fd_sc_hd__inv_2 _4451__36 (.A(clknet_leaf_86_wb_clk_i),
    .Y(net767));
 sky130_fd_sc_hd__inv_2 _4452__37 (.A(clknet_leaf_88_wb_clk_i),
    .Y(net768));
 sky130_fd_sc_hd__inv_2 _4453__38 (.A(clknet_leaf_89_wb_clk_i),
    .Y(net769));
 sky130_fd_sc_hd__inv_2 _4454__39 (.A(clknet_leaf_88_wb_clk_i),
    .Y(net770));
 sky130_fd_sc_hd__inv_2 _4455__40 (.A(clknet_leaf_93_wb_clk_i),
    .Y(net771));
 sky130_fd_sc_hd__inv_2 _4456__41 (.A(clknet_leaf_77_wb_clk_i),
    .Y(net772));
 sky130_fd_sc_hd__inv_2 _4457__42 (.A(clknet_leaf_85_wb_clk_i),
    .Y(net773));
 sky130_fd_sc_hd__inv_2 _4458__43 (.A(clknet_leaf_76_wb_clk_i),
    .Y(net774));
 sky130_fd_sc_hd__inv_2 _4459__44 (.A(clknet_leaf_102_wb_clk_i),
    .Y(net775));
 sky130_fd_sc_hd__inv_2 _4460__45 (.A(clknet_leaf_78_wb_clk_i),
    .Y(net776));
 sky130_fd_sc_hd__inv_2 _4461__46 (.A(clknet_leaf_74_wb_clk_i),
    .Y(net777));
 sky130_fd_sc_hd__inv_2 _4462__47 (.A(clknet_leaf_79_wb_clk_i),
    .Y(net778));
 sky130_fd_sc_hd__inv_2 _4463__48 (.A(clknet_leaf_79_wb_clk_i),
    .Y(net779));
 sky130_fd_sc_hd__inv_2 _4464__49 (.A(clknet_leaf_39_wb_clk_i),
    .Y(net780));
 sky130_fd_sc_hd__inv_2 _4465__50 (.A(clknet_leaf_39_wb_clk_i),
    .Y(net781));
 sky130_fd_sc_hd__inv_2 _4466__51 (.A(clknet_leaf_51_wb_clk_i),
    .Y(net782));
 sky130_fd_sc_hd__inv_2 _4467__52 (.A(clknet_leaf_51_wb_clk_i),
    .Y(net783));
 sky130_fd_sc_hd__inv_2 _4468__53 (.A(clknet_leaf_38_wb_clk_i),
    .Y(net784));
 sky130_fd_sc_hd__inv_2 _4469__54 (.A(clknet_leaf_51_wb_clk_i),
    .Y(net785));
 sky130_fd_sc_hd__inv_2 _4470__55 (.A(clknet_leaf_52_wb_clk_i),
    .Y(net786));
 sky130_fd_sc_hd__inv_2 _4471__56 (.A(clknet_leaf_50_wb_clk_i),
    .Y(net787));
 sky130_fd_sc_hd__inv_2 _4472__57 (.A(clknet_leaf_40_wb_clk_i),
    .Y(net788));
 sky130_fd_sc_hd__inv_2 _4473__58 (.A(clknet_leaf_32_wb_clk_i),
    .Y(net789));
 sky130_fd_sc_hd__inv_2 _4474__59 (.A(clknet_leaf_25_wb_clk_i),
    .Y(net790));
 sky130_fd_sc_hd__inv_2 _4475__60 (.A(clknet_leaf_33_wb_clk_i),
    .Y(net791));
 sky130_fd_sc_hd__inv_2 _4476__61 (.A(clknet_leaf_22_wb_clk_i),
    .Y(net792));
 sky130_fd_sc_hd__inv_2 _4477__62 (.A(clknet_leaf_21_wb_clk_i),
    .Y(net793));
 sky130_fd_sc_hd__inv_2 _4478__63 (.A(clknet_leaf_22_wb_clk_i),
    .Y(net794));
 sky130_fd_sc_hd__inv_2 _4479__64 (.A(clknet_leaf_26_wb_clk_i),
    .Y(net795));
 sky130_fd_sc_hd__inv_2 _4480__65 (.A(clknet_leaf_48_wb_clk_i),
    .Y(net796));
 sky130_fd_sc_hd__inv_2 _4481__66 (.A(clknet_leaf_49_wb_clk_i),
    .Y(net797));
 sky130_fd_sc_hd__inv_2 _4482__67 (.A(clknet_leaf_49_wb_clk_i),
    .Y(net798));
 sky130_fd_sc_hd__inv_2 _4483__68 (.A(clknet_leaf_58_wb_clk_i),
    .Y(net799));
 sky130_fd_sc_hd__inv_2 _4484__69 (.A(clknet_leaf_64_wb_clk_i),
    .Y(net800));
 sky130_fd_sc_hd__inv_2 _4485__70 (.A(clknet_leaf_68_wb_clk_i),
    .Y(net801));
 sky130_fd_sc_hd__inv_2 _4486__71 (.A(clknet_leaf_64_wb_clk_i),
    .Y(net802));
 sky130_fd_sc_hd__inv_2 _4487__72 (.A(clknet_leaf_65_wb_clk_i),
    .Y(net803));
 sky130_fd_sc_hd__inv_2 _4488__73 (.A(clknet_leaf_34_wb_clk_i),
    .Y(net804));
 sky130_fd_sc_hd__inv_2 _4489__74 (.A(clknet_leaf_32_wb_clk_i),
    .Y(net805));
 sky130_fd_sc_hd__inv_2 _4490__75 (.A(clknet_leaf_32_wb_clk_i),
    .Y(net806));
 sky130_fd_sc_hd__inv_2 _4491__76 (.A(clknet_leaf_34_wb_clk_i),
    .Y(net807));
 sky130_fd_sc_hd__inv_2 _4492__77 (.A(clknet_leaf_27_wb_clk_i),
    .Y(net808));
 sky130_fd_sc_hd__inv_2 _4493__78 (.A(clknet_leaf_26_wb_clk_i),
    .Y(net809));
 sky130_fd_sc_hd__inv_2 _4494__79 (.A(clknet_leaf_25_wb_clk_i),
    .Y(net810));
 sky130_fd_sc_hd__inv_2 _4495__80 (.A(clknet_leaf_28_wb_clk_i),
    .Y(net811));
 sky130_fd_sc_hd__inv_2 _4496__81 (.A(clknet_leaf_34_wb_clk_i),
    .Y(net812));
 sky130_fd_sc_hd__inv_2 _4497__82 (.A(clknet_leaf_32_wb_clk_i),
    .Y(net813));
 sky130_fd_sc_hd__inv_2 _4498__83 (.A(clknet_leaf_32_wb_clk_i),
    .Y(net814));
 sky130_fd_sc_hd__inv_2 _4499__84 (.A(clknet_leaf_34_wb_clk_i),
    .Y(net815));
 sky130_fd_sc_hd__inv_2 _4500__85 (.A(clknet_leaf_27_wb_clk_i),
    .Y(net816));
 sky130_fd_sc_hd__inv_2 _4501__86 (.A(clknet_leaf_26_wb_clk_i),
    .Y(net817));
 sky130_fd_sc_hd__inv_2 _4502__87 (.A(clknet_leaf_25_wb_clk_i),
    .Y(net818));
 sky130_fd_sc_hd__inv_2 _4503__88 (.A(clknet_leaf_28_wb_clk_i),
    .Y(net819));
 sky130_fd_sc_hd__inv_2 _4504__89 (.A(clknet_leaf_34_wb_clk_i),
    .Y(net820));
 sky130_fd_sc_hd__inv_2 _4505__90 (.A(clknet_leaf_32_wb_clk_i),
    .Y(net821));
 sky130_fd_sc_hd__inv_2 _4506__91 (.A(clknet_leaf_32_wb_clk_i),
    .Y(net822));
 sky130_fd_sc_hd__inv_2 _4507__92 (.A(clknet_leaf_33_wb_clk_i),
    .Y(net823));
 sky130_fd_sc_hd__inv_2 _4508__93 (.A(clknet_leaf_27_wb_clk_i),
    .Y(net824));
 sky130_fd_sc_hd__inv_2 _4509__94 (.A(clknet_leaf_26_wb_clk_i),
    .Y(net825));
 sky130_fd_sc_hd__inv_2 _4510__95 (.A(clknet_leaf_25_wb_clk_i),
    .Y(net826));
 sky130_fd_sc_hd__inv_2 _4511__96 (.A(clknet_leaf_28_wb_clk_i),
    .Y(net827));
 sky130_fd_sc_hd__inv_2 _4512__97 (.A(clknet_leaf_48_wb_clk_i),
    .Y(net828));
 sky130_fd_sc_hd__inv_2 _4513__98 (.A(clknet_leaf_70_wb_clk_i),
    .Y(net829));
 sky130_fd_sc_hd__inv_2 _4514__99 (.A(clknet_leaf_69_wb_clk_i),
    .Y(net830));
 sky130_fd_sc_hd__inv_2 _4515__100 (.A(clknet_leaf_70_wb_clk_i),
    .Y(net831));
 sky130_fd_sc_hd__inv_2 _4516__101 (.A(clknet_leaf_68_wb_clk_i),
    .Y(net832));
 sky130_fd_sc_hd__inv_2 _4517__102 (.A(clknet_leaf_68_wb_clk_i),
    .Y(net833));
 sky130_fd_sc_hd__inv_2 _4518__103 (.A(clknet_leaf_64_wb_clk_i),
    .Y(net834));
 sky130_fd_sc_hd__inv_2 _4519__104 (.A(clknet_leaf_65_wb_clk_i),
    .Y(net835));
 sky130_fd_sc_hd__inv_2 _4520__105 (.A(clknet_leaf_41_wb_clk_i),
    .Y(net836));
 sky130_fd_sc_hd__inv_2 _4521__106 (.A(clknet_leaf_24_wb_clk_i),
    .Y(net837));
 sky130_fd_sc_hd__inv_2 _4522__107 (.A(clknet_leaf_23_wb_clk_i),
    .Y(net838));
 sky130_fd_sc_hd__inv_2 _4523__108 (.A(clknet_leaf_15_wb_clk_i),
    .Y(net839));
 sky130_fd_sc_hd__inv_2 _4524__109 (.A(clknet_leaf_22_wb_clk_i),
    .Y(net840));
 sky130_fd_sc_hd__inv_2 _4525__110 (.A(clknet_leaf_21_wb_clk_i),
    .Y(net841));
 sky130_fd_sc_hd__inv_2 _4526__111 (.A(clknet_leaf_25_wb_clk_i),
    .Y(net842));
 sky130_fd_sc_hd__inv_2 _4527__112 (.A(clknet_leaf_26_wb_clk_i),
    .Y(net843));
 sky130_fd_sc_hd__inv_2 _4528__113 (.A(clknet_leaf_14_wb_clk_i),
    .Y(net844));
 sky130_fd_sc_hd__inv_2 _4529__114 (.A(clknet_leaf_15_wb_clk_i),
    .Y(net845));
 sky130_fd_sc_hd__inv_2 _4530__115 (.A(clknet_leaf_23_wb_clk_i),
    .Y(net846));
 sky130_fd_sc_hd__inv_2 _4531__116 (.A(clknet_leaf_15_wb_clk_i),
    .Y(net847));
 sky130_fd_sc_hd__inv_2 _4532__117 (.A(clknet_leaf_18_wb_clk_i),
    .Y(net848));
 sky130_fd_sc_hd__inv_2 _4533__118 (.A(clknet_leaf_19_wb_clk_i),
    .Y(net849));
 sky130_fd_sc_hd__inv_2 _4534__119 (.A(clknet_leaf_20_wb_clk_i),
    .Y(net850));
 sky130_fd_sc_hd__inv_2 _4535__120 (.A(clknet_leaf_22_wb_clk_i),
    .Y(net851));
 sky130_fd_sc_hd__inv_2 _4536__121 (.A(clknet_leaf_35_wb_clk_i),
    .Y(net852));
 sky130_fd_sc_hd__inv_2 _4537__122 (.A(clknet_leaf_31_wb_clk_i),
    .Y(net853));
 sky130_fd_sc_hd__inv_2 _4538__123 (.A(clknet_leaf_31_wb_clk_i),
    .Y(net854));
 sky130_fd_sc_hd__inv_2 _4539__124 (.A(clknet_leaf_35_wb_clk_i),
    .Y(net855));
 sky130_fd_sc_hd__inv_2 _4540__125 (.A(clknet_leaf_30_wb_clk_i),
    .Y(net856));
 sky130_fd_sc_hd__inv_2 _4541__126 (.A(clknet_leaf_29_wb_clk_i),
    .Y(net857));
 sky130_fd_sc_hd__inv_2 _4542__127 (.A(clknet_leaf_29_wb_clk_i),
    .Y(net858));
 sky130_fd_sc_hd__inv_2 _4543__128 (.A(clknet_leaf_30_wb_clk_i),
    .Y(net859));
 sky130_fd_sc_hd__inv_2 _4544__129 (.A(clknet_leaf_36_wb_clk_i),
    .Y(net860));
 sky130_fd_sc_hd__inv_2 _4545__130 (.A(clknet_leaf_31_wb_clk_i),
    .Y(net861));
 sky130_fd_sc_hd__inv_2 _4546__131 (.A(clknet_leaf_31_wb_clk_i),
    .Y(net862));
 sky130_fd_sc_hd__inv_2 _4547__132 (.A(clknet_leaf_35_wb_clk_i),
    .Y(net863));
 sky130_fd_sc_hd__inv_2 _4548__133 (.A(clknet_leaf_30_wb_clk_i),
    .Y(net864));
 sky130_fd_sc_hd__inv_2 _4549__134 (.A(clknet_leaf_29_wb_clk_i),
    .Y(net865));
 sky130_fd_sc_hd__inv_2 _4550__135 (.A(clknet_leaf_28_wb_clk_i),
    .Y(net866));
 sky130_fd_sc_hd__inv_2 _4551__136 (.A(clknet_leaf_30_wb_clk_i),
    .Y(net867));
 sky130_fd_sc_hd__inv_2 _4552__137 (.A(clknet_leaf_36_wb_clk_i),
    .Y(net868));
 sky130_fd_sc_hd__inv_2 _4553__138 (.A(clknet_leaf_31_wb_clk_i),
    .Y(net869));
 sky130_fd_sc_hd__inv_2 _4554__139 (.A(clknet_leaf_31_wb_clk_i),
    .Y(net870));
 sky130_fd_sc_hd__inv_2 _4555__140 (.A(clknet_leaf_35_wb_clk_i),
    .Y(net871));
 sky130_fd_sc_hd__inv_2 _4556__141 (.A(clknet_leaf_31_wb_clk_i),
    .Y(net872));
 sky130_fd_sc_hd__inv_2 _4557__142 (.A(clknet_leaf_29_wb_clk_i),
    .Y(net873));
 sky130_fd_sc_hd__inv_2 _4558__143 (.A(clknet_leaf_29_wb_clk_i),
    .Y(net874));
 sky130_fd_sc_hd__inv_2 _4559__144 (.A(clknet_leaf_30_wb_clk_i),
    .Y(net875));
 sky130_fd_sc_hd__inv_2 _4560__145 (.A(clknet_leaf_34_wb_clk_i),
    .Y(net876));
 sky130_fd_sc_hd__inv_2 _4561__146 (.A(clknet_leaf_32_wb_clk_i),
    .Y(net877));
 sky130_fd_sc_hd__inv_2 _4562__147 (.A(clknet_leaf_32_wb_clk_i),
    .Y(net878));
 sky130_fd_sc_hd__inv_2 _4563__148 (.A(clknet_leaf_33_wb_clk_i),
    .Y(net879));
 sky130_fd_sc_hd__inv_2 _4564__149 (.A(clknet_leaf_27_wb_clk_i),
    .Y(net880));
 sky130_fd_sc_hd__inv_2 _4565__150 (.A(clknet_leaf_26_wb_clk_i),
    .Y(net881));
 sky130_fd_sc_hd__inv_2 _4566__151 (.A(clknet_leaf_27_wb_clk_i),
    .Y(net882));
 sky130_fd_sc_hd__inv_2 _4567__152 (.A(clknet_leaf_27_wb_clk_i),
    .Y(net883));
 sky130_fd_sc_hd__inv_2 _4568__153 (.A(clknet_leaf_41_wb_clk_i),
    .Y(net884));
 sky130_fd_sc_hd__inv_2 _4569__154 (.A(clknet_leaf_24_wb_clk_i),
    .Y(net885));
 sky130_fd_sc_hd__inv_2 _4570__155 (.A(clknet_leaf_24_wb_clk_i),
    .Y(net886));
 sky130_fd_sc_hd__inv_2 _4571__156 (.A(clknet_leaf_41_wb_clk_i),
    .Y(net887));
 sky130_fd_sc_hd__inv_2 _4572__157 (.A(clknet_leaf_19_wb_clk_i),
    .Y(net888));
 sky130_fd_sc_hd__inv_2 _4573__158 (.A(clknet_leaf_19_wb_clk_i),
    .Y(net889));
 sky130_fd_sc_hd__inv_2 _4574__159 (.A(clknet_leaf_20_wb_clk_i),
    .Y(net890));
 sky130_fd_sc_hd__inv_2 _4575__160 (.A(clknet_leaf_20_wb_clk_i),
    .Y(net891));
 sky130_fd_sc_hd__inv_2 _4576__161 (.A(clknet_leaf_41_wb_clk_i),
    .Y(net892));
 sky130_fd_sc_hd__inv_2 _4577__162 (.A(clknet_leaf_24_wb_clk_i),
    .Y(net893));
 sky130_fd_sc_hd__inv_2 _4578__163 (.A(clknet_leaf_25_wb_clk_i),
    .Y(net894));
 sky130_fd_sc_hd__inv_2 _4579__164 (.A(clknet_leaf_33_wb_clk_i),
    .Y(net895));
 sky130_fd_sc_hd__inv_2 _4580__165 (.A(clknet_leaf_21_wb_clk_i),
    .Y(net896));
 sky130_fd_sc_hd__inv_2 _4581__166 (.A(clknet_leaf_21_wb_clk_i),
    .Y(net897));
 sky130_fd_sc_hd__inv_2 _4582__167 (.A(clknet_leaf_25_wb_clk_i),
    .Y(net898));
 sky130_fd_sc_hd__inv_2 _4583__168 (.A(clknet_leaf_26_wb_clk_i),
    .Y(net899));
 sky130_fd_sc_hd__inv_2 _4584__169 (.A(clknet_leaf_14_wb_clk_i),
    .Y(net900));
 sky130_fd_sc_hd__inv_2 _4585__170 (.A(clknet_leaf_15_wb_clk_i),
    .Y(net901));
 sky130_fd_sc_hd__inv_2 _4586__171 (.A(clknet_leaf_23_wb_clk_i),
    .Y(net902));
 sky130_fd_sc_hd__inv_2 _4587__172 (.A(clknet_leaf_15_wb_clk_i),
    .Y(net903));
 sky130_fd_sc_hd__inv_2 _4588__173 (.A(clknet_leaf_19_wb_clk_i),
    .Y(net904));
 sky130_fd_sc_hd__inv_2 _4589__174 (.A(clknet_leaf_19_wb_clk_i),
    .Y(net905));
 sky130_fd_sc_hd__inv_2 _4590__175 (.A(clknet_leaf_20_wb_clk_i),
    .Y(net906));
 sky130_fd_sc_hd__inv_2 _4591__176 (.A(clknet_leaf_20_wb_clk_i),
    .Y(net907));
 sky130_fd_sc_hd__inv_2 _4592__177 (.A(clknet_leaf_83_wb_clk_i),
    .Y(net908));
 sky130_fd_sc_hd__inv_2 _4593__178 (.A(clknet_leaf_87_wb_clk_i),
    .Y(net909));
 sky130_fd_sc_hd__inv_2 _4594__179 (.A(clknet_leaf_84_wb_clk_i),
    .Y(net910));
 sky130_fd_sc_hd__inv_2 _4595__180 (.A(clknet_leaf_83_wb_clk_i),
    .Y(net911));
 sky130_fd_sc_hd__inv_2 _4596__181 (.A(clknet_leaf_78_wb_clk_i),
    .Y(net912));
 sky130_fd_sc_hd__inv_2 _4597__182 (.A(clknet_leaf_81_wb_clk_i),
    .Y(net913));
 sky130_fd_sc_hd__inv_2 _4598__183 (.A(clknet_leaf_81_wb_clk_i),
    .Y(net914));
 sky130_fd_sc_hd__inv_2 _4599__184 (.A(clknet_leaf_80_wb_clk_i),
    .Y(net915));
 sky130_fd_sc_hd__inv_2 _4600__185 (.A(clknet_leaf_84_wb_clk_i),
    .Y(net916));
 sky130_fd_sc_hd__inv_2 _4601__186 (.A(clknet_leaf_84_wb_clk_i),
    .Y(net917));
 sky130_fd_sc_hd__inv_2 _4602__187 (.A(clknet_leaf_77_wb_clk_i),
    .Y(net918));
 sky130_fd_sc_hd__inv_2 _4603__188 (.A(clknet_leaf_77_wb_clk_i),
    .Y(net919));
 sky130_fd_sc_hd__inv_2 _4604__189 (.A(clknet_leaf_75_wb_clk_i),
    .Y(net920));
 sky130_fd_sc_hd__inv_2 _4605__190 (.A(clknet_leaf_74_wb_clk_i),
    .Y(net921));
 sky130_fd_sc_hd__inv_2 _4606__191 (.A(clknet_leaf_79_wb_clk_i),
    .Y(net922));
 sky130_fd_sc_hd__inv_2 _4607__192 (.A(clknet_leaf_79_wb_clk_i),
    .Y(net923));
 sky130_fd_sc_hd__inv_2 _4608__193 (.A(clknet_leaf_0_wb_clk_i),
    .Y(net924));
 sky130_fd_sc_hd__inv_2 _4609__194 (.A(clknet_leaf_0_wb_clk_i),
    .Y(net925));
 sky130_fd_sc_hd__inv_2 _4610__195 (.A(clknet_leaf_118_wb_clk_i),
    .Y(net926));
 sky130_fd_sc_hd__inv_2 _4611__196 (.A(clknet_leaf_0_wb_clk_i),
    .Y(net927));
 sky130_fd_sc_hd__inv_2 _4612__197 (.A(clknet_leaf_0_wb_clk_i),
    .Y(net928));
 sky130_fd_sc_hd__inv_2 _4613__198 (.A(clknet_leaf_121_wb_clk_i),
    .Y(net929));
 sky130_fd_sc_hd__inv_2 _4614__199 (.A(clknet_leaf_120_wb_clk_i),
    .Y(net930));
 sky130_fd_sc_hd__inv_2 _4615__200 (.A(clknet_leaf_119_wb_clk_i),
    .Y(net931));
 sky130_fd_sc_hd__inv_2 _4616__201 (.A(clknet_leaf_83_wb_clk_i),
    .Y(net932));
 sky130_fd_sc_hd__inv_2 _4617__202 (.A(clknet_leaf_83_wb_clk_i),
    .Y(net933));
 sky130_fd_sc_hd__inv_2 _4618__203 (.A(clknet_leaf_84_wb_clk_i),
    .Y(net934));
 sky130_fd_sc_hd__inv_2 _4619__204 (.A(clknet_leaf_83_wb_clk_i),
    .Y(net935));
 sky130_fd_sc_hd__inv_2 _4620__205 (.A(clknet_leaf_80_wb_clk_i),
    .Y(net936));
 sky130_fd_sc_hd__inv_2 _4621__206 (.A(clknet_leaf_81_wb_clk_i),
    .Y(net937));
 sky130_fd_sc_hd__inv_2 _4622__207 (.A(clknet_leaf_81_wb_clk_i),
    .Y(net938));
 sky130_fd_sc_hd__inv_2 _4623__208 (.A(clknet_leaf_80_wb_clk_i),
    .Y(net939));
 sky130_fd_sc_hd__inv_2 _4624__209 (.A(clknet_leaf_77_wb_clk_i),
    .Y(net940));
 sky130_fd_sc_hd__inv_2 _4625__210 (.A(clknet_leaf_85_wb_clk_i),
    .Y(net941));
 sky130_fd_sc_hd__inv_2 _4626__211 (.A(clknet_leaf_76_wb_clk_i),
    .Y(net942));
 sky130_fd_sc_hd__inv_2 _4627__212 (.A(clknet_leaf_102_wb_clk_i),
    .Y(net943));
 sky130_fd_sc_hd__inv_2 _4628__213 (.A(clknet_leaf_78_wb_clk_i),
    .Y(net944));
 sky130_fd_sc_hd__inv_2 _4629__214 (.A(clknet_leaf_74_wb_clk_i),
    .Y(net945));
 sky130_fd_sc_hd__inv_2 _4630__215 (.A(clknet_leaf_79_wb_clk_i),
    .Y(net946));
 sky130_fd_sc_hd__inv_2 _4631__216 (.A(clknet_leaf_78_wb_clk_i),
    .Y(net947));
 sky130_fd_sc_hd__inv_2 _4632__217 (.A(clknet_leaf_48_wb_clk_i),
    .Y(net948));
 sky130_fd_sc_hd__inv_2 _4633__218 (.A(clknet_leaf_70_wb_clk_i),
    .Y(net949));
 sky130_fd_sc_hd__inv_2 _4634__219 (.A(clknet_leaf_69_wb_clk_i),
    .Y(net950));
 sky130_fd_sc_hd__inv_2 _4635__220 (.A(clknet_leaf_70_wb_clk_i),
    .Y(net951));
 sky130_fd_sc_hd__inv_2 _4636__221 (.A(clknet_leaf_69_wb_clk_i),
    .Y(net952));
 sky130_fd_sc_hd__inv_2 _4637__222 (.A(clknet_leaf_68_wb_clk_i),
    .Y(net953));
 sky130_fd_sc_hd__inv_2 _4638__223 (.A(clknet_leaf_64_wb_clk_i),
    .Y(net954));
 sky130_fd_sc_hd__inv_2 _4639__224 (.A(clknet_leaf_68_wb_clk_i),
    .Y(net955));
 sky130_fd_sc_hd__inv_2 _4640__225 (.A(clknet_leaf_94_wb_clk_i),
    .Y(net956));
 sky130_fd_sc_hd__inv_2 _4641__226 (.A(clknet_leaf_94_wb_clk_i),
    .Y(net957));
 sky130_fd_sc_hd__inv_2 _4642__227 (.A(clknet_leaf_94_wb_clk_i),
    .Y(net958));
 sky130_fd_sc_hd__inv_2 _4643__228 (.A(clknet_leaf_101_wb_clk_i),
    .Y(net959));
 sky130_fd_sc_hd__inv_2 _4644__229 (.A(clknet_leaf_101_wb_clk_i),
    .Y(net960));
 sky130_fd_sc_hd__inv_2 _4645__230 (.A(clknet_leaf_104_wb_clk_i),
    .Y(net961));
 sky130_fd_sc_hd__inv_2 _4646__231 (.A(clknet_leaf_104_wb_clk_i),
    .Y(net962));
 sky130_fd_sc_hd__inv_2 _4647__232 (.A(clknet_leaf_100_wb_clk_i),
    .Y(net963));
 sky130_fd_sc_hd__inv_2 _4648__233 (.A(clknet_leaf_100_wb_clk_i),
    .Y(net964));
 sky130_fd_sc_hd__inv_2 _4649__234 (.A(clknet_leaf_100_wb_clk_i),
    .Y(net965));
 sky130_fd_sc_hd__inv_2 _4650__235 (.A(clknet_leaf_9_wb_clk_i),
    .Y(net966));
 sky130_fd_sc_hd__inv_2 _4651__236 (.A(clknet_leaf_101_wb_clk_i),
    .Y(net967));
 sky130_fd_sc_hd__inv_2 _4652__237 (.A(clknet_leaf_102_wb_clk_i),
    .Y(net968));
 sky130_fd_sc_hd__inv_2 _4653__238 (.A(clknet_leaf_103_wb_clk_i),
    .Y(net969));
 sky130_fd_sc_hd__inv_2 _4654__239 (.A(clknet_leaf_103_wb_clk_i),
    .Y(net970));
 sky130_fd_sc_hd__inv_2 _4655__240 (.A(clknet_leaf_102_wb_clk_i),
    .Y(net971));
 sky130_fd_sc_hd__inv_2 _4656__241 (.A(clknet_leaf_102_wb_clk_i),
    .Y(net972));
 sky130_fd_sc_hd__inv_2 _4657__242 (.A(clknet_leaf_102_wb_clk_i),
    .Y(net973));
 sky130_fd_sc_hd__inv_2 _4658__243 (.A(clknet_leaf_101_wb_clk_i),
    .Y(net974));
 sky130_fd_sc_hd__inv_2 _4659__244 (.A(clknet_leaf_41_wb_clk_i),
    .Y(net975));
 sky130_fd_sc_hd__inv_2 _4660__245 (.A(clknet_leaf_24_wb_clk_i),
    .Y(net976));
 sky130_fd_sc_hd__inv_2 _4661__246 (.A(clknet_leaf_23_wb_clk_i),
    .Y(net977));
 sky130_fd_sc_hd__inv_2 _4662__247 (.A(clknet_leaf_15_wb_clk_i),
    .Y(net978));
 sky130_fd_sc_hd__inv_2 _4663__248 (.A(clknet_leaf_22_wb_clk_i),
    .Y(net979));
 sky130_fd_sc_hd__inv_2 _4664__249 (.A(clknet_leaf_21_wb_clk_i),
    .Y(net980));
 sky130_fd_sc_hd__inv_2 _4665__250 (.A(clknet_leaf_21_wb_clk_i),
    .Y(net981));
 sky130_fd_sc_hd__inv_2 _4666__251 (.A(clknet_leaf_21_wb_clk_i),
    .Y(net982));
 sky130_fd_sc_hd__inv_2 _4667__252 (.A(clknet_leaf_48_wb_clk_i),
    .Y(net983));
 sky130_fd_sc_hd__inv_2 _4668__253 (.A(clknet_leaf_49_wb_clk_i),
    .Y(net984));
 sky130_fd_sc_hd__inv_2 _4669__254 (.A(clknet_leaf_49_wb_clk_i),
    .Y(net985));
 sky130_fd_sc_hd__inv_2 _4670__255 (.A(clknet_leaf_58_wb_clk_i),
    .Y(net986));
 sky130_fd_sc_hd__inv_2 _4671__256 (.A(clknet_leaf_69_wb_clk_i),
    .Y(net987));
 sky130_fd_sc_hd__inv_2 _4672__257 (.A(clknet_leaf_68_wb_clk_i),
    .Y(net988));
 sky130_fd_sc_hd__inv_2 _4673__258 (.A(clknet_leaf_64_wb_clk_i),
    .Y(net989));
 sky130_fd_sc_hd__inv_2 _4674__259 (.A(clknet_leaf_68_wb_clk_i),
    .Y(net990));
 sky130_fd_sc_hd__inv_2 _4675__260 (.A(clknet_leaf_14_wb_clk_i),
    .Y(net991));
 sky130_fd_sc_hd__inv_2 _4676__261 (.A(clknet_4_9_0_wb_clk_i),
    .Y(net992));
 sky130_fd_sc_hd__inv_2 _4677__262 (.A(clknet_leaf_43_wb_clk_i),
    .Y(net993));
 sky130_fd_sc_hd__inv_2 _4678__263 (.A(clknet_leaf_43_wb_clk_i),
    .Y(net994));
 sky130_fd_sc_hd__inv_2 _4679__264 (.A(clknet_leaf_41_wb_clk_i),
    .Y(net995));
 sky130_fd_sc_hd__inv_2 _4680__265 (.A(clknet_leaf_44_wb_clk_i),
    .Y(net996));
 sky130_fd_sc_hd__inv_2 _4681__266 (.A(clknet_leaf_44_wb_clk_i),
    .Y(net997));
 sky130_fd_sc_hd__inv_2 _4682__267 (.A(clknet_leaf_43_wb_clk_i),
    .Y(net998));
 sky130_fd_sc_hd__inv_2 _4683__268 (.A(clknet_leaf_43_wb_clk_i),
    .Y(net999));
 sky130_fd_sc_hd__inv_2 _4684__269 (.A(clknet_leaf_43_wb_clk_i),
    .Y(net1000));
 sky130_fd_sc_hd__inv_2 _4685__270 (.A(clknet_leaf_14_wb_clk_i),
    .Y(net1001));
 sky130_fd_sc_hd__inv_2 _4686__271 (.A(clknet_leaf_14_wb_clk_i),
    .Y(net1002));
 sky130_fd_sc_hd__inv_2 _4687__272 (.A(clknet_leaf_16_wb_clk_i),
    .Y(net1003));
 sky130_fd_sc_hd__inv_2 _4688__273 (.A(clknet_leaf_16_wb_clk_i),
    .Y(net1004));
 sky130_fd_sc_hd__inv_2 _4689__274 (.A(clknet_leaf_14_wb_clk_i),
    .Y(net1005));
 sky130_fd_sc_hd__inv_2 _4690__275 (.A(clknet_leaf_16_wb_clk_i),
    .Y(net1006));
 sky130_fd_sc_hd__inv_2 _4691__276 (.A(clknet_leaf_16_wb_clk_i),
    .Y(net1007));
 sky130_fd_sc_hd__inv_2 _4692__277 (.A(clknet_leaf_14_wb_clk_i),
    .Y(net1008));
 sky130_fd_sc_hd__inv_2 _4693__278 (.A(clknet_leaf_14_wb_clk_i),
    .Y(net1009));
 sky130_fd_sc_hd__inv_2 _4694__279 (.A(clknet_leaf_115_wb_clk_i),
    .Y(net1010));
 sky130_fd_sc_hd__inv_2 _4695__280 (.A(clknet_leaf_111_wb_clk_i),
    .Y(net1011));
 sky130_fd_sc_hd__inv_2 _4696__281 (.A(clknet_leaf_110_wb_clk_i),
    .Y(net1012));
 sky130_fd_sc_hd__inv_2 _4697__282 (.A(clknet_leaf_115_wb_clk_i),
    .Y(net1013));
 sky130_fd_sc_hd__inv_2 _4698__283 (.A(clknet_leaf_114_wb_clk_i),
    .Y(net1014));
 sky130_fd_sc_hd__inv_2 _4699__284 (.A(clknet_leaf_113_wb_clk_i),
    .Y(net1015));
 sky130_fd_sc_hd__inv_2 _4700__285 (.A(clknet_leaf_114_wb_clk_i),
    .Y(net1016));
 sky130_fd_sc_hd__inv_2 _4701__286 (.A(clknet_leaf_112_wb_clk_i),
    .Y(net1017));
 sky130_fd_sc_hd__inv_2 _4702__287 (.A(clknet_leaf_50_wb_clk_i),
    .Y(net1018));
 sky130_fd_sc_hd__inv_2 _4703__288 (.A(clknet_leaf_54_wb_clk_i),
    .Y(net1019));
 sky130_fd_sc_hd__inv_2 _4704__289 (.A(clknet_leaf_56_wb_clk_i),
    .Y(net1020));
 sky130_fd_sc_hd__inv_2 _4705__290 (.A(clknet_leaf_55_wb_clk_i),
    .Y(net1021));
 sky130_fd_sc_hd__inv_2 _4706__291 (.A(clknet_leaf_59_wb_clk_i),
    .Y(net1022));
 sky130_fd_sc_hd__inv_2 _4707__292 (.A(clknet_leaf_58_wb_clk_i),
    .Y(net1023));
 sky130_fd_sc_hd__inv_2 _4708__293 (.A(clknet_leaf_59_wb_clk_i),
    .Y(net1024));
 sky130_fd_sc_hd__inv_2 _4709__294 (.A(clknet_leaf_63_wb_clk_i),
    .Y(net1025));
 sky130_fd_sc_hd__inv_2 _4710__295 (.A(clknet_leaf_50_wb_clk_i),
    .Y(net1026));
 sky130_fd_sc_hd__inv_2 _4711__296 (.A(clknet_leaf_54_wb_clk_i),
    .Y(net1027));
 sky130_fd_sc_hd__inv_2 _4712__297 (.A(clknet_leaf_56_wb_clk_i),
    .Y(net1028));
 sky130_fd_sc_hd__inv_2 _4713__298 (.A(clknet_leaf_60_wb_clk_i),
    .Y(net1029));
 sky130_fd_sc_hd__inv_2 _4714__299 (.A(clknet_leaf_59_wb_clk_i),
    .Y(net1030));
 sky130_fd_sc_hd__inv_2 _4715__300 (.A(clknet_leaf_59_wb_clk_i),
    .Y(net1031));
 sky130_fd_sc_hd__inv_2 _4716__301 (.A(clknet_leaf_61_wb_clk_i),
    .Y(net1032));
 sky130_fd_sc_hd__inv_2 _4717__302 (.A(clknet_leaf_63_wb_clk_i),
    .Y(net1033));
 sky130_fd_sc_hd__inv_2 _4718__303 (.A(clknet_leaf_113_wb_clk_i),
    .Y(net1034));
 sky130_fd_sc_hd__inv_2 _4719__304 (.A(clknet_leaf_111_wb_clk_i),
    .Y(net1035));
 sky130_fd_sc_hd__inv_2 _4720__305 (.A(clknet_leaf_111_wb_clk_i),
    .Y(net1036));
 sky130_fd_sc_hd__inv_2 _4721__306 (.A(clknet_leaf_115_wb_clk_i),
    .Y(net1037));
 sky130_fd_sc_hd__inv_2 _4722__307 (.A(clknet_leaf_113_wb_clk_i),
    .Y(net1038));
 sky130_fd_sc_hd__inv_2 _4723__308 (.A(clknet_leaf_113_wb_clk_i),
    .Y(net1039));
 sky130_fd_sc_hd__inv_2 _4724__309 (.A(clknet_leaf_115_wb_clk_i),
    .Y(net1040));
 sky130_fd_sc_hd__inv_2 _4725__310 (.A(clknet_leaf_112_wb_clk_i),
    .Y(net1041));
 sky130_fd_sc_hd__inv_2 _4726__311 (.A(clknet_leaf_111_wb_clk_i),
    .Y(net1042));
 sky130_fd_sc_hd__inv_2 _4727__312 (.A(clknet_leaf_111_wb_clk_i),
    .Y(net1043));
 sky130_fd_sc_hd__inv_2 _4728__313 (.A(clknet_leaf_112_wb_clk_i),
    .Y(net1044));
 sky130_fd_sc_hd__inv_2 _4729__314 (.A(clknet_leaf_113_wb_clk_i),
    .Y(net1045));
 sky130_fd_sc_hd__inv_2 _4730__315 (.A(clknet_leaf_113_wb_clk_i),
    .Y(net1046));
 sky130_fd_sc_hd__inv_2 _4731__316 (.A(clknet_leaf_113_wb_clk_i),
    .Y(net1047));
 sky130_fd_sc_hd__inv_2 _4732__317 (.A(clknet_leaf_114_wb_clk_i),
    .Y(net1048));
 sky130_fd_sc_hd__inv_2 _4733__318 (.A(clknet_leaf_111_wb_clk_i),
    .Y(net1049));
 sky130_fd_sc_hd__inv_2 _4734__319 (.A(clknet_leaf_57_wb_clk_i),
    .Y(net1050));
 sky130_fd_sc_hd__inv_2 _4735__320 (.A(clknet_leaf_56_wb_clk_i),
    .Y(net1051));
 sky130_fd_sc_hd__inv_2 _4736__321 (.A(clknet_leaf_56_wb_clk_i),
    .Y(net1052));
 sky130_fd_sc_hd__inv_2 _4737__322 (.A(clknet_leaf_57_wb_clk_i),
    .Y(net1053));
 sky130_fd_sc_hd__inv_2 _4738__323 (.A(clknet_leaf_59_wb_clk_i),
    .Y(net1054));
 sky130_fd_sc_hd__inv_2 _4739__324 (.A(clknet_leaf_59_wb_clk_i),
    .Y(net1055));
 sky130_fd_sc_hd__inv_2 _4740__325 (.A(clknet_leaf_59_wb_clk_i),
    .Y(net1056));
 sky130_fd_sc_hd__inv_2 _4741__326 (.A(clknet_leaf_63_wb_clk_i),
    .Y(net1057));
 sky130_fd_sc_hd__inv_2 _4742__327 (.A(clknet_leaf_57_wb_clk_i),
    .Y(net1058));
 sky130_fd_sc_hd__inv_2 _4743__328 (.A(clknet_leaf_56_wb_clk_i),
    .Y(net1059));
 sky130_fd_sc_hd__inv_2 _4744__329 (.A(clknet_leaf_56_wb_clk_i),
    .Y(net1060));
 sky130_fd_sc_hd__inv_2 _4745__330 (.A(clknet_leaf_57_wb_clk_i),
    .Y(net1061));
 sky130_fd_sc_hd__inv_2 _4746__331 (.A(clknet_leaf_59_wb_clk_i),
    .Y(net1062));
 sky130_fd_sc_hd__inv_2 _4747__332 (.A(clknet_leaf_58_wb_clk_i),
    .Y(net1063));
 sky130_fd_sc_hd__inv_2 _4748__333 (.A(clknet_leaf_61_wb_clk_i),
    .Y(net1064));
 sky130_fd_sc_hd__inv_2 _4749__334 (.A(clknet_leaf_63_wb_clk_i),
    .Y(net1065));
 sky130_fd_sc_hd__inv_2 _4750__335 (.A(clknet_leaf_1_wb_clk_i),
    .Y(net1066));
 sky130_fd_sc_hd__inv_2 _4751__336 (.A(clknet_leaf_4_wb_clk_i),
    .Y(net1067));
 sky130_fd_sc_hd__inv_2 _4752__337 (.A(clknet_leaf_3_wb_clk_i),
    .Y(net1068));
 sky130_fd_sc_hd__inv_2 _4753__338 (.A(clknet_leaf_1_wb_clk_i),
    .Y(net1069));
 sky130_fd_sc_hd__inv_2 _4754__339 (.A(clknet_leaf_1_wb_clk_i),
    .Y(net1070));
 sky130_fd_sc_hd__inv_2 _4755__340 (.A(clknet_leaf_2_wb_clk_i),
    .Y(net1071));
 sky130_fd_sc_hd__inv_2 _4756__341 (.A(clknet_leaf_118_wb_clk_i),
    .Y(net1072));
 sky130_fd_sc_hd__inv_2 _4757__342 (.A(clknet_leaf_2_wb_clk_i),
    .Y(net1073));
 sky130_fd_sc_hd__inv_2 _4758__343 (.A(clknet_leaf_36_wb_clk_i),
    .Y(net1074));
 sky130_fd_sc_hd__inv_2 _4759__344 (.A(clknet_leaf_37_wb_clk_i),
    .Y(net1075));
 sky130_fd_sc_hd__inv_2 _4760__345 (.A(clknet_leaf_52_wb_clk_i),
    .Y(net1076));
 sky130_fd_sc_hd__inv_2 _4761__346 (.A(clknet_leaf_52_wb_clk_i),
    .Y(net1077));
 sky130_fd_sc_hd__inv_2 _4762__347 (.A(clknet_leaf_36_wb_clk_i),
    .Y(net1078));
 sky130_fd_sc_hd__inv_2 _4763__348 (.A(clknet_leaf_37_wb_clk_i),
    .Y(net1079));
 sky130_fd_sc_hd__inv_2 _4764__349 (.A(clknet_leaf_53_wb_clk_i),
    .Y(net1080));
 sky130_fd_sc_hd__inv_2 _4765__350 (.A(clknet_leaf_54_wb_clk_i),
    .Y(net1081));
 sky130_fd_sc_hd__inv_2 _4766__351 (.A(clknet_leaf_1_wb_clk_i),
    .Y(net1082));
 sky130_fd_sc_hd__inv_2 _4767__352 (.A(clknet_leaf_4_wb_clk_i),
    .Y(net1083));
 sky130_fd_sc_hd__inv_2 _4768__353 (.A(clknet_leaf_3_wb_clk_i),
    .Y(net1084));
 sky130_fd_sc_hd__inv_2 _4769__354 (.A(clknet_leaf_1_wb_clk_i),
    .Y(net1085));
 sky130_fd_sc_hd__inv_2 _4770__355 (.A(clknet_leaf_1_wb_clk_i),
    .Y(net1086));
 sky130_fd_sc_hd__inv_2 _4771__356 (.A(clknet_leaf_2_wb_clk_i),
    .Y(net1087));
 sky130_fd_sc_hd__inv_2 _4772__357 (.A(clknet_leaf_118_wb_clk_i),
    .Y(net1088));
 sky130_fd_sc_hd__inv_2 _4773__358 (.A(clknet_leaf_2_wb_clk_i),
    .Y(net1089));
 sky130_fd_sc_hd__inv_2 _4774__359 (.A(clknet_leaf_116_wb_clk_i),
    .Y(net1090));
 sky130_fd_sc_hd__inv_2 _4775__360 (.A(clknet_leaf_117_wb_clk_i),
    .Y(net1091));
 sky130_fd_sc_hd__inv_2 _4776__361 (.A(clknet_leaf_117_wb_clk_i),
    .Y(net1092));
 sky130_fd_sc_hd__inv_2 _4777__362 (.A(clknet_leaf_0_wb_clk_i),
    .Y(net1093));
 sky130_fd_sc_hd__inv_2 _4778__363 (.A(clknet_leaf_121_wb_clk_i),
    .Y(net1094));
 sky130_fd_sc_hd__inv_2 _4779__364 (.A(clknet_leaf_121_wb_clk_i),
    .Y(net1095));
 sky130_fd_sc_hd__inv_2 _4780__365 (.A(clknet_leaf_120_wb_clk_i),
    .Y(net1096));
 sky130_fd_sc_hd__inv_2 _4781__366 (.A(clknet_leaf_119_wb_clk_i),
    .Y(net1097));
 sky130_fd_sc_hd__inv_2 _4782__367 (.A(clknet_leaf_118_wb_clk_i),
    .Y(net1098));
 sky130_fd_sc_hd__inv_2 _4783__368 (.A(clknet_leaf_110_wb_clk_i),
    .Y(net1099));
 sky130_fd_sc_hd__inv_2 _4784__369 (.A(clknet_leaf_110_wb_clk_i),
    .Y(net1100));
 sky130_fd_sc_hd__inv_2 _4785__370 (.A(clknet_leaf_110_wb_clk_i),
    .Y(net1101));
 sky130_fd_sc_hd__inv_2 _4786__371 (.A(clknet_leaf_1_wb_clk_i),
    .Y(net1102));
 sky130_fd_sc_hd__inv_2 _4787__372 (.A(clknet_leaf_2_wb_clk_i),
    .Y(net1103));
 sky130_fd_sc_hd__inv_2 _4788__373 (.A(clknet_leaf_118_wb_clk_i),
    .Y(net1104));
 sky130_fd_sc_hd__inv_2 _4789__374 (.A(clknet_leaf_2_wb_clk_i),
    .Y(net1105));
 sky130_fd_sc_hd__inv_2 _4790__375 (.A(clknet_leaf_95_wb_clk_i),
    .Y(net1106));
 sky130_fd_sc_hd__inv_2 _4791__376 (.A(clknet_leaf_99_wb_clk_i),
    .Y(net1107));
 sky130_fd_sc_hd__inv_2 _4792__377 (.A(clknet_leaf_99_wb_clk_i),
    .Y(net1108));
 sky130_fd_sc_hd__inv_2 _4793__378 (.A(clknet_leaf_97_wb_clk_i),
    .Y(net1109));
 sky130_fd_sc_hd__inv_2 _4794__379 (.A(clknet_leaf_98_wb_clk_i),
    .Y(net1110));
 sky130_fd_sc_hd__inv_2 _4795__380 (.A(clknet_leaf_97_wb_clk_i),
    .Y(net1111));
 sky130_fd_sc_hd__inv_2 _4796__381 (.A(clknet_leaf_98_wb_clk_i),
    .Y(net1112));
 sky130_fd_sc_hd__inv_2 _4797__382 (.A(clknet_leaf_98_wb_clk_i),
    .Y(net1113));
 sky130_fd_sc_hd__inv_2 _4798__383 (.A(clknet_leaf_95_wb_clk_i),
    .Y(net1114));
 sky130_fd_sc_hd__inv_2 _4799__384 (.A(clknet_leaf_99_wb_clk_i),
    .Y(net1115));
 sky130_fd_sc_hd__inv_2 _4800__385 (.A(clknet_leaf_99_wb_clk_i),
    .Y(net1116));
 sky130_fd_sc_hd__inv_2 _4801__386 (.A(clknet_leaf_97_wb_clk_i),
    .Y(net1117));
 sky130_fd_sc_hd__inv_2 _4802__387 (.A(clknet_leaf_98_wb_clk_i),
    .Y(net1118));
 sky130_fd_sc_hd__inv_2 _4803__388 (.A(clknet_leaf_96_wb_clk_i),
    .Y(net1119));
 sky130_fd_sc_hd__inv_2 _4804__389 (.A(clknet_leaf_98_wb_clk_i),
    .Y(net1120));
 sky130_fd_sc_hd__inv_2 _4805__390 (.A(clknet_leaf_99_wb_clk_i),
    .Y(net1121));
 sky130_fd_sc_hd__inv_2 _4806__391 (.A(clknet_leaf_95_wb_clk_i),
    .Y(net1122));
 sky130_fd_sc_hd__inv_2 _4807__392 (.A(clknet_leaf_99_wb_clk_i),
    .Y(net1123));
 sky130_fd_sc_hd__inv_2 _4808__393 (.A(clknet_leaf_99_wb_clk_i),
    .Y(net1124));
 sky130_fd_sc_hd__inv_2 _4809__394 (.A(clknet_leaf_97_wb_clk_i),
    .Y(net1125));
 sky130_fd_sc_hd__inv_2 _4810__395 (.A(clknet_leaf_97_wb_clk_i),
    .Y(net1126));
 sky130_fd_sc_hd__inv_2 _4811__396 (.A(clknet_leaf_97_wb_clk_i),
    .Y(net1127));
 sky130_fd_sc_hd__inv_2 _4812__397 (.A(clknet_leaf_98_wb_clk_i),
    .Y(net1128));
 sky130_fd_sc_hd__inv_2 _4813__398 (.A(clknet_leaf_98_wb_clk_i),
    .Y(net1129));
 sky130_fd_sc_hd__inv_2 _4814__399 (.A(clknet_leaf_99_wb_clk_i),
    .Y(net1130));
 sky130_fd_sc_hd__inv_2 _4815__400 (.A(clknet_leaf_97_wb_clk_i),
    .Y(net1131));
 sky130_fd_sc_hd__inv_2 _4816__401 (.A(clknet_leaf_99_wb_clk_i),
    .Y(net1132));
 sky130_fd_sc_hd__inv_2 _4817__402 (.A(clknet_leaf_97_wb_clk_i),
    .Y(net1133));
 sky130_fd_sc_hd__inv_2 _4818__403 (.A(clknet_leaf_98_wb_clk_i),
    .Y(net1134));
 sky130_fd_sc_hd__inv_2 _4819__404 (.A(clknet_leaf_97_wb_clk_i),
    .Y(net1135));
 sky130_fd_sc_hd__inv_2 _4820__405 (.A(clknet_leaf_98_wb_clk_i),
    .Y(net1136));
 sky130_fd_sc_hd__inv_2 _4821__406 (.A(clknet_leaf_98_wb_clk_i),
    .Y(net1137));
 sky130_fd_sc_hd__inv_2 _4822__407 (.A(clknet_leaf_0_wb_clk_i),
    .Y(net1138));
 sky130_fd_sc_hd__inv_2 _4823__408 (.A(clknet_leaf_0_wb_clk_i),
    .Y(net1139));
 sky130_fd_sc_hd__inv_2 _4824__409 (.A(clknet_leaf_119_wb_clk_i),
    .Y(net1140));
 sky130_fd_sc_hd__inv_2 _4825__410 (.A(clknet_leaf_0_wb_clk_i),
    .Y(net1141));
 sky130_fd_sc_hd__inv_2 _4826__411 (.A(clknet_leaf_121_wb_clk_i),
    .Y(net1142));
 sky130_fd_sc_hd__inv_2 _4827__412 (.A(clknet_leaf_121_wb_clk_i),
    .Y(net1143));
 sky130_fd_sc_hd__inv_2 _4828__413 (.A(clknet_leaf_120_wb_clk_i),
    .Y(net1144));
 sky130_fd_sc_hd__inv_2 _4829__414 (.A(clknet_leaf_119_wb_clk_i),
    .Y(net1145));
 sky130_fd_sc_hd__inv_2 _4830__415 (.A(clknet_leaf_78_wb_clk_i),
    .Y(net1146));
 sky130_fd_sc_hd__inv_2 _4831__416 (.A(clknet_leaf_84_wb_clk_i),
    .Y(net1147));
 sky130_fd_sc_hd__inv_2 _4832__417 (.A(clknet_leaf_77_wb_clk_i),
    .Y(net1148));
 sky130_fd_sc_hd__inv_2 _4833__418 (.A(clknet_leaf_77_wb_clk_i),
    .Y(net1149));
 sky130_fd_sc_hd__inv_2 _4834__419 (.A(clknet_leaf_78_wb_clk_i),
    .Y(net1150));
 sky130_fd_sc_hd__inv_2 _4835__420 (.A(clknet_leaf_74_wb_clk_i),
    .Y(net1151));
 sky130_fd_sc_hd__inv_2 _4836__421 (.A(clknet_leaf_79_wb_clk_i),
    .Y(net1152));
 sky130_fd_sc_hd__inv_2 _4837__422 (.A(clknet_leaf_79_wb_clk_i),
    .Y(net1153));
 sky130_fd_sc_hd__inv_2 _4838__423 (.A(clknet_leaf_39_wb_clk_i),
    .Y(net1154));
 sky130_fd_sc_hd__inv_2 _4839__424 (.A(clknet_leaf_47_wb_clk_i),
    .Y(net1155));
 sky130_fd_sc_hd__inv_2 _4840__425 (.A(clknet_leaf_47_wb_clk_i),
    .Y(net1156));
 sky130_fd_sc_hd__inv_2 _4841__426 (.A(clknet_leaf_47_wb_clk_i),
    .Y(net1157));
 sky130_fd_sc_hd__inv_2 _4842__427 (.A(clknet_leaf_38_wb_clk_i),
    .Y(net1158));
 sky130_fd_sc_hd__inv_2 _4843__428 (.A(clknet_leaf_38_wb_clk_i),
    .Y(net1159));
 sky130_fd_sc_hd__inv_2 _4844__429 (.A(clknet_leaf_38_wb_clk_i),
    .Y(net1160));
 sky130_fd_sc_hd__inv_2 _4845__430 (.A(clknet_leaf_50_wb_clk_i),
    .Y(net1161));
 sky130_fd_sc_hd__inv_2 _4846__431 (.A(clknet_leaf_36_wb_clk_i),
    .Y(net1162));
 sky130_fd_sc_hd__inv_2 _4847__432 (.A(clknet_leaf_37_wb_clk_i),
    .Y(net1163));
 sky130_fd_sc_hd__inv_2 _4848__433 (.A(clknet_leaf_54_wb_clk_i),
    .Y(net1164));
 sky130_fd_sc_hd__inv_2 _4849__434 (.A(clknet_leaf_52_wb_clk_i),
    .Y(net1165));
 sky130_fd_sc_hd__inv_2 _4850__435 (.A(clknet_leaf_36_wb_clk_i),
    .Y(net1166));
 sky130_fd_sc_hd__inv_2 _4851__436 (.A(clknet_leaf_37_wb_clk_i),
    .Y(net1167));
 sky130_fd_sc_hd__inv_2 _4852__437 (.A(clknet_leaf_53_wb_clk_i),
    .Y(net1168));
 sky130_fd_sc_hd__inv_2 _4853__438 (.A(clknet_leaf_54_wb_clk_i),
    .Y(net1169));
 sky130_fd_sc_hd__inv_2 _4854__439 (.A(clknet_leaf_90_wb_clk_i),
    .Y(net1170));
 sky130_fd_sc_hd__inv_2 _4855__440 (.A(clknet_leaf_91_wb_clk_i),
    .Y(net1171));
 sky130_fd_sc_hd__inv_2 _4856__441 (.A(clknet_leaf_91_wb_clk_i),
    .Y(net1172));
 sky130_fd_sc_hd__inv_2 _4857__442 (.A(clknet_leaf_88_wb_clk_i),
    .Y(net1173));
 sky130_fd_sc_hd__inv_2 _4858__443 (.A(clknet_leaf_96_wb_clk_i),
    .Y(net1174));
 sky130_fd_sc_hd__inv_2 _4859__444 (.A(clknet_leaf_90_wb_clk_i),
    .Y(net1175));
 sky130_fd_sc_hd__inv_2 _4860__445 (.A(clknet_leaf_91_wb_clk_i),
    .Y(net1176));
 sky130_fd_sc_hd__inv_2 _4861__446 (.A(clknet_leaf_96_wb_clk_i),
    .Y(net1177));
 sky130_fd_sc_hd__inv_2 _4862__447 (.A(clknet_leaf_36_wb_clk_i),
    .Y(net1178));
 sky130_fd_sc_hd__inv_2 _4863__448 (.A(clknet_leaf_37_wb_clk_i),
    .Y(net1179));
 sky130_fd_sc_hd__inv_2 _4864__449 (.A(clknet_leaf_52_wb_clk_i),
    .Y(net1180));
 sky130_fd_sc_hd__inv_2 _4865__450 (.A(clknet_leaf_52_wb_clk_i),
    .Y(net1181));
 sky130_fd_sc_hd__inv_2 _4866__451 (.A(clknet_leaf_36_wb_clk_i),
    .Y(net1182));
 sky130_fd_sc_hd__inv_2 _4867__452 (.A(clknet_leaf_37_wb_clk_i),
    .Y(net1183));
 sky130_fd_sc_hd__inv_2 _4868__453 (.A(clknet_leaf_53_wb_clk_i),
    .Y(net1184));
 sky130_fd_sc_hd__inv_2 _4869__454 (.A(clknet_leaf_54_wb_clk_i),
    .Y(net1185));
 sky130_fd_sc_hd__inv_2 _4870__455 (.A(clknet_leaf_90_wb_clk_i),
    .Y(net1186));
 sky130_fd_sc_hd__inv_2 _4871__456 (.A(clknet_leaf_90_wb_clk_i),
    .Y(net1187));
 sky130_fd_sc_hd__inv_2 _4872__457 (.A(clknet_leaf_91_wb_clk_i),
    .Y(net1188));
 sky130_fd_sc_hd__inv_2 _4873__458 (.A(clknet_leaf_90_wb_clk_i),
    .Y(net1189));
 sky130_fd_sc_hd__inv_2 _4874__459 (.A(clknet_leaf_96_wb_clk_i),
    .Y(net1190));
 sky130_fd_sc_hd__inv_2 _4875__460 (.A(clknet_leaf_90_wb_clk_i),
    .Y(net1191));
 sky130_fd_sc_hd__inv_2 _4876__461 (.A(clknet_leaf_91_wb_clk_i),
    .Y(net1192));
 sky130_fd_sc_hd__inv_2 _4877__462 (.A(clknet_leaf_92_wb_clk_i),
    .Y(net1193));
 sky130_fd_sc_hd__inv_2 _4878__463 (.A(clknet_leaf_36_wb_clk_i),
    .Y(net1194));
 sky130_fd_sc_hd__inv_2 _4879__464 (.A(clknet_leaf_37_wb_clk_i),
    .Y(net1195));
 sky130_fd_sc_hd__inv_2 _4880__465 (.A(clknet_leaf_52_wb_clk_i),
    .Y(net1196));
 sky130_fd_sc_hd__inv_2 _4881__466 (.A(clknet_leaf_52_wb_clk_i),
    .Y(net1197));
 sky130_fd_sc_hd__inv_2 _4882__467 (.A(clknet_leaf_36_wb_clk_i),
    .Y(net1198));
 sky130_fd_sc_hd__inv_2 _4883__468 (.A(clknet_leaf_37_wb_clk_i),
    .Y(net1199));
 sky130_fd_sc_hd__inv_2 _4884__469 (.A(clknet_leaf_53_wb_clk_i),
    .Y(net1200));
 sky130_fd_sc_hd__inv_2 _4885__470 (.A(clknet_leaf_53_wb_clk_i),
    .Y(net1201));
 sky130_fd_sc_hd__inv_2 _4886__471 (.A(clknet_leaf_95_wb_clk_i),
    .Y(net1202));
 sky130_fd_sc_hd__inv_2 _4887__472 (.A(clknet_leaf_92_wb_clk_i),
    .Y(net1203));
 sky130_fd_sc_hd__inv_2 _4888__473 (.A(clknet_leaf_94_wb_clk_i),
    .Y(net1204));
 sky130_fd_sc_hd__inv_2 _4889__474 (.A(clknet_leaf_95_wb_clk_i),
    .Y(net1205));
 sky130_fd_sc_hd__inv_2 _4890__475 (.A(clknet_leaf_96_wb_clk_i),
    .Y(net1206));
 sky130_fd_sc_hd__inv_2 _4891__476 (.A(clknet_leaf_91_wb_clk_i),
    .Y(net1207));
 sky130_fd_sc_hd__inv_2 _4892__477 (.A(clknet_leaf_91_wb_clk_i),
    .Y(net1208));
 sky130_fd_sc_hd__inv_2 _4893__478 (.A(clknet_leaf_92_wb_clk_i),
    .Y(net1209));
 sky130_fd_sc_hd__inv_2 _4894__479 (.A(clknet_leaf_95_wb_clk_i),
    .Y(net1210));
 sky130_fd_sc_hd__inv_2 _4895__480 (.A(clknet_leaf_92_wb_clk_i),
    .Y(net1211));
 sky130_fd_sc_hd__inv_2 _4896__481 (.A(clknet_leaf_94_wb_clk_i),
    .Y(net1212));
 sky130_fd_sc_hd__inv_2 _4897__482 (.A(clknet_leaf_95_wb_clk_i),
    .Y(net1213));
 sky130_fd_sc_hd__inv_2 _4898__483 (.A(clknet_leaf_96_wb_clk_i),
    .Y(net1214));
 sky130_fd_sc_hd__inv_2 _4899__484 (.A(clknet_leaf_92_wb_clk_i),
    .Y(net1215));
 sky130_fd_sc_hd__inv_2 _4900__485 (.A(clknet_leaf_92_wb_clk_i),
    .Y(net1216));
 sky130_fd_sc_hd__inv_2 _4901__486 (.A(clknet_leaf_92_wb_clk_i),
    .Y(net1217));
 sky130_fd_sc_hd__inv_2 _4902__487 (.A(clknet_leaf_116_wb_clk_i),
    .Y(net1218));
 sky130_fd_sc_hd__inv_2 _4903__488 (.A(clknet_leaf_117_wb_clk_i),
    .Y(net1219));
 sky130_fd_sc_hd__inv_2 _4904__489 (.A(clknet_leaf_117_wb_clk_i),
    .Y(net1220));
 sky130_fd_sc_hd__inv_2 _4905__490 (.A(clknet_leaf_0_wb_clk_i),
    .Y(net1221));
 sky130_fd_sc_hd__inv_2 _4906__491 (.A(clknet_leaf_121_wb_clk_i),
    .Y(net1222));
 sky130_fd_sc_hd__inv_2 _4907__492 (.A(clknet_leaf_120_wb_clk_i),
    .Y(net1223));
 sky130_fd_sc_hd__inv_2 _4908__493 (.A(clknet_leaf_120_wb_clk_i),
    .Y(net1224));
 sky130_fd_sc_hd__inv_2 _4909__494 (.A(clknet_leaf_119_wb_clk_i),
    .Y(net1225));
 sky130_fd_sc_hd__inv_2 _4910__495 (.A(clknet_leaf_87_wb_clk_i),
    .Y(net1226));
 sky130_fd_sc_hd__inv_2 _4911__496 (.A(clknet_leaf_87_wb_clk_i),
    .Y(net1227));
 sky130_fd_sc_hd__inv_2 _4912__497 (.A(clknet_leaf_86_wb_clk_i),
    .Y(net1228));
 sky130_fd_sc_hd__inv_2 _4913__498 (.A(clknet_leaf_86_wb_clk_i),
    .Y(net1229));
 sky130_fd_sc_hd__inv_2 _4914__499 (.A(clknet_leaf_88_wb_clk_i),
    .Y(net1230));
 sky130_fd_sc_hd__inv_2 _4915__500 (.A(clknet_leaf_88_wb_clk_i),
    .Y(net1231));
 sky130_fd_sc_hd__inv_2 _4916__501 (.A(clknet_leaf_89_wb_clk_i),
    .Y(net1232));
 sky130_fd_sc_hd__inv_2 _4917__502 (.A(clknet_leaf_93_wb_clk_i),
    .Y(net1233));
 sky130_fd_sc_hd__inv_2 _4918__503 (.A(clknet_leaf_85_wb_clk_i),
    .Y(net1234));
 sky130_fd_sc_hd__inv_2 _4919__504 (.A(clknet_leaf_86_wb_clk_i),
    .Y(net1235));
 sky130_fd_sc_hd__inv_2 _4920__505 (.A(clknet_leaf_94_wb_clk_i),
    .Y(net1236));
 sky130_fd_sc_hd__inv_2 _4921__506 (.A(clknet_leaf_94_wb_clk_i),
    .Y(net1237));
 sky130_fd_sc_hd__inv_2 _4922__507 (.A(clknet_leaf_88_wb_clk_i),
    .Y(net1238));
 sky130_fd_sc_hd__inv_2 _4923__508 (.A(clknet_leaf_89_wb_clk_i),
    .Y(net1239));
 sky130_fd_sc_hd__inv_2 _4924__509 (.A(clknet_leaf_88_wb_clk_i),
    .Y(net1240));
 sky130_fd_sc_hd__inv_2 _4925__510 (.A(clknet_leaf_93_wb_clk_i),
    .Y(net1241));
 sky130_fd_sc_hd__inv_2 _4926__511 (.A(clknet_leaf_86_wb_clk_i),
    .Y(net1242));
 sky130_fd_sc_hd__inv_2 _4927__512 (.A(clknet_leaf_86_wb_clk_i),
    .Y(net1243));
 sky130_fd_sc_hd__inv_2 _4928__513 (.A(clknet_leaf_93_wb_clk_i),
    .Y(net1244));
 sky130_fd_sc_hd__inv_2 _4929__514 (.A(clknet_leaf_86_wb_clk_i),
    .Y(net1245));
 sky130_fd_sc_hd__inv_2 _4930__515 (.A(clknet_leaf_86_wb_clk_i),
    .Y(net1246));
 sky130_fd_sc_hd__inv_2 _4931__516 (.A(clknet_leaf_88_wb_clk_i),
    .Y(net1247));
 sky130_fd_sc_hd__inv_2 _4932__517 (.A(clknet_leaf_88_wb_clk_i),
    .Y(net1248));
 sky130_fd_sc_hd__inv_2 _4933__518 (.A(clknet_leaf_93_wb_clk_i),
    .Y(net1249));
 sky130_fd_sc_hd__inv_2 _4934__519 (.A(clknet_leaf_115_wb_clk_i),
    .Y(net1250));
 sky130_fd_sc_hd__inv_2 _4935__520 (.A(clknet_leaf_117_wb_clk_i),
    .Y(net1251));
 sky130_fd_sc_hd__inv_2 _4936__521 (.A(clknet_leaf_110_wb_clk_i),
    .Y(net1252));
 sky130_fd_sc_hd__inv_2 _4937__522 (.A(clknet_leaf_117_wb_clk_i),
    .Y(net1253));
 sky130_fd_sc_hd__inv_2 _4938__523 (.A(clknet_leaf_114_wb_clk_i),
    .Y(net1254));
 sky130_fd_sc_hd__inv_2 _4939__524 (.A(clknet_leaf_114_wb_clk_i),
    .Y(net1255));
 sky130_fd_sc_hd__inv_2 _4940__525 (.A(clknet_leaf_115_wb_clk_i),
    .Y(net1256));
 sky130_fd_sc_hd__inv_2 _4941__526 (.A(clknet_leaf_111_wb_clk_i),
    .Y(net1257));
 sky130_fd_sc_hd__inv_2 _4942__527 (.A(clknet_leaf_83_wb_clk_i),
    .Y(net1258));
 sky130_fd_sc_hd__inv_2 _4943__528 (.A(clknet_leaf_83_wb_clk_i),
    .Y(net1259));
 sky130_fd_sc_hd__inv_2 _4944__529 (.A(clknet_leaf_84_wb_clk_i),
    .Y(net1260));
 sky130_fd_sc_hd__inv_2 _4945__530 (.A(clknet_leaf_84_wb_clk_i),
    .Y(net1261));
 sky130_fd_sc_hd__inv_2 _4946__531 (.A(clknet_leaf_80_wb_clk_i),
    .Y(net1262));
 sky130_fd_sc_hd__inv_2 _4947__532 (.A(clknet_leaf_80_wb_clk_i),
    .Y(net1263));
 sky130_fd_sc_hd__inv_2 _4948__533 (.A(clknet_leaf_81_wb_clk_i),
    .Y(net1264));
 sky130_fd_sc_hd__inv_2 _4949__534 (.A(clknet_leaf_80_wb_clk_i),
    .Y(net1265));
 sky130_fd_sc_hd__inv_2 _4950__535 (.A(clknet_leaf_118_wb_clk_i),
    .Y(net1266));
 sky130_fd_sc_hd__inv_2 _4951__536 (.A(clknet_leaf_110_wb_clk_i),
    .Y(net1267));
 sky130_fd_sc_hd__inv_2 _4952__537 (.A(clknet_leaf_110_wb_clk_i),
    .Y(net1268));
 sky130_fd_sc_hd__inv_2 _4953__538 (.A(clknet_leaf_110_wb_clk_i),
    .Y(net1269));
 sky130_fd_sc_hd__inv_2 _4954__539 (.A(clknet_leaf_118_wb_clk_i),
    .Y(net1270));
 sky130_fd_sc_hd__inv_2 _4955__540 (.A(clknet_leaf_118_wb_clk_i),
    .Y(net1271));
 sky130_fd_sc_hd__inv_2 _4956__541 (.A(clknet_leaf_118_wb_clk_i),
    .Y(net1272));
 sky130_fd_sc_hd__inv_2 _4957__542 (.A(clknet_leaf_2_wb_clk_i),
    .Y(net1273));
 sky130_fd_sc_hd__inv_2 _4958__543 (.A(clknet_leaf_83_wb_clk_i),
    .Y(net1274));
 sky130_fd_sc_hd__inv_2 _4959__544 (.A(clknet_leaf_83_wb_clk_i),
    .Y(net1275));
 sky130_fd_sc_hd__inv_2 _4960__545 (.A(clknet_leaf_84_wb_clk_i),
    .Y(net1276));
 sky130_fd_sc_hd__inv_2 _4961__546 (.A(clknet_leaf_83_wb_clk_i),
    .Y(net1277));
 sky130_fd_sc_hd__inv_2 _4962__547 (.A(clknet_4_7_0_wb_clk_i),
    .Y(net1278));
 sky130_fd_sc_hd__inv_2 _4963__548 (.A(clknet_leaf_81_wb_clk_i),
    .Y(net1279));
 sky130_fd_sc_hd__inv_2 _4964__549 (.A(clknet_leaf_81_wb_clk_i),
    .Y(net1280));
 sky130_fd_sc_hd__inv_2 _4965__550 (.A(clknet_leaf_80_wb_clk_i),
    .Y(net1281));
 sky130_fd_sc_hd__dfxtp_2 _4966_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(net3490),
    .Q(hostConfigLatch));
 sky130_fd_sc_hd__dfxtp_1 _4967_ (.CLK(net732),
    .D(_0955_),
    .Q(\device.rxBuffer.buffer[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4968_ (.CLK(net733),
    .D(_0956_),
    .Q(\device.rxBuffer.buffer[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4969_ (.CLK(net734),
    .D(_0957_),
    .Q(\device.rxBuffer.buffer[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4970_ (.CLK(net735),
    .D(_0958_),
    .Q(\device.rxBuffer.buffer[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4971_ (.CLK(net736),
    .D(_0959_),
    .Q(\device.rxBuffer.buffer[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4972_ (.CLK(net737),
    .D(_0960_),
    .Q(\device.rxBuffer.buffer[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4973_ (.CLK(net738),
    .D(_0961_),
    .Q(\device.rxBuffer.buffer[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4974_ (.CLK(net739),
    .D(_0962_),
    .Q(\device.rxBuffer.buffer[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4975_ (.CLK(net740),
    .D(_0963_),
    .Q(\device.rxBuffer.buffer[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4976_ (.CLK(net741),
    .D(_0964_),
    .Q(\device.rxBuffer.buffer[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4977_ (.CLK(net742),
    .D(_0965_),
    .Q(\device.rxBuffer.buffer[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4978_ (.CLK(net743),
    .D(_0966_),
    .Q(\device.rxBuffer.buffer[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4979_ (.CLK(net744),
    .D(_0967_),
    .Q(\device.rxBuffer.buffer[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4980_ (.CLK(net745),
    .D(_0968_),
    .Q(\device.rxBuffer.buffer[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4981_ (.CLK(net746),
    .D(_0969_),
    .Q(\device.rxBuffer.buffer[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4982_ (.CLK(net747),
    .D(_0970_),
    .Q(\device.rxBuffer.buffer[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4983_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(net3386),
    .Q(\wbAddressExtension.dataRead_buffered[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4984_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(net3393),
    .Q(\wbAddressExtension.dataRead_buffered[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4985_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net1735),
    .Q(\wbAddressExtension.dataRead_buffered[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4986_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(net3365),
    .Q(\wbAddressExtension.dataRead_buffered[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4987_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(net3358),
    .Q(\wbAddressExtension.dataRead_buffered[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4988_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(net3379),
    .Q(\wbAddressExtension.dataRead_buffered[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4989_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(net3372),
    .Q(\wbAddressExtension.dataRead_buffered[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4990_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(net3311),
    .Q(\wbAddressExtension.dataRead_buffered[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4991_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(net3323),
    .Q(\wbAddressExtension.dataRead_buffered[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4992_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(net3317),
    .Q(\wbAddressExtension.dataRead_buffered[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4993_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(net3282),
    .Q(\wbAddressExtension.dataRead_buffered[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4994_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(net3294),
    .Q(\wbAddressExtension.dataRead_buffered[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4995_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(net3288),
    .Q(\wbAddressExtension.dataRead_buffered[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4996_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(net3340),
    .Q(\wbAddressExtension.dataRead_buffered[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4997_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(net3479),
    .Q(\wbAddressExtension.dataRead_buffered[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4998_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0986_),
    .Q(\wbAddressExtension.dataRead_buffered[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4999_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0987_),
    .Q(\wbAddressExtension.dataRead_buffered[16] ));
 sky130_fd_sc_hd__dfxtp_1 _5000_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0988_),
    .Q(\wbAddressExtension.dataRead_buffered[17] ));
 sky130_fd_sc_hd__dfxtp_1 _5001_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0989_),
    .Q(\wbAddressExtension.dataRead_buffered[18] ));
 sky130_fd_sc_hd__dfxtp_1 _5002_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1540),
    .Q(\wbAddressExtension.dataRead_buffered[19] ));
 sky130_fd_sc_hd__dfxtp_1 _5003_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0991_),
    .Q(\wbAddressExtension.dataRead_buffered[20] ));
 sky130_fd_sc_hd__dfxtp_1 _5004_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0992_),
    .Q(\wbAddressExtension.dataRead_buffered[21] ));
 sky130_fd_sc_hd__dfxtp_1 _5005_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net1531),
    .Q(\wbAddressExtension.dataRead_buffered[22] ));
 sky130_fd_sc_hd__dfxtp_1 _5006_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(net1527),
    .Q(\wbAddressExtension.dataRead_buffered[23] ));
 sky130_fd_sc_hd__dfxtp_1 _5007_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(net1559),
    .Q(\wbAddressExtension.dataRead_buffered[24] ));
 sky130_fd_sc_hd__dfxtp_1 _5008_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(net1563),
    .Q(\wbAddressExtension.dataRead_buffered[25] ));
 sky130_fd_sc_hd__dfxtp_1 _5009_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(net1569),
    .Q(\wbAddressExtension.dataRead_buffered[26] ));
 sky130_fd_sc_hd__dfxtp_1 _5010_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(net1549),
    .Q(\wbAddressExtension.dataRead_buffered[27] ));
 sky130_fd_sc_hd__dfxtp_1 _5011_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(net1646),
    .Q(\wbAddressExtension.dataRead_buffered[28] ));
 sky130_fd_sc_hd__dfxtp_1 _5012_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_1000_),
    .Q(\wbAddressExtension.dataRead_buffered[29] ));
 sky130_fd_sc_hd__dfxtp_1 _5013_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(net1640),
    .Q(\wbAddressExtension.dataRead_buffered[30] ));
 sky130_fd_sc_hd__dfxtp_1 _5014_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_1002_),
    .Q(\wbAddressExtension.dataRead_buffered[31] ));
 sky130_fd_sc_hd__dfxtp_1 _5015_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_1003_),
    .Q(\wbAddressExtension.currentAddress[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5016_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_1004_),
    .Q(\wbAddressExtension.currentAddress[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5017_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net1340),
    .Q(\wbAddressExtension.currentAddress[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5018_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(net1353),
    .Q(\wbAddressExtension.currentAddress[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5019_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_1007_),
    .Q(\wbAddressExtension.currentAddress[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5020_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_1008_),
    .Q(\wbAddressExtension.currentAddress[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5021_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_1009_),
    .Q(\wbAddressExtension.currentAddress[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5022_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(net1362),
    .Q(\wbAddressExtension.currentAddress[7] ));
 sky130_fd_sc_hd__dfxtp_2 _5023_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net3120),
    .Q(\wbAddressExtension.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5024_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net3148),
    .Q(\wbAddressExtension.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5025_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_1013_),
    .Q(net206));
 sky130_fd_sc_hd__dfxtp_1 _5026_ (.CLK(net748),
    .D(_1014_),
    .Q(\device.rxBuffer.buffer[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5027_ (.CLK(net749),
    .D(_1015_),
    .Q(\device.rxBuffer.buffer[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5028_ (.CLK(net750),
    .D(_1016_),
    .Q(\device.rxBuffer.buffer[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5029_ (.CLK(net751),
    .D(_1017_),
    .Q(\device.rxBuffer.buffer[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5030_ (.CLK(net752),
    .D(_1018_),
    .Q(\device.rxBuffer.buffer[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5031_ (.CLK(net753),
    .D(_1019_),
    .Q(\device.rxBuffer.buffer[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5032_ (.CLK(net754),
    .D(_1020_),
    .Q(\device.rxBuffer.buffer[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5033_ (.CLK(net755),
    .D(_1021_),
    .Q(\device.rxBuffer.buffer[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5034_ (.CLK(net756),
    .D(_1022_),
    .Q(\device.rxBuffer.buffer[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5035_ (.CLK(net757),
    .D(_1023_),
    .Q(\device.rxBuffer.buffer[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5036_ (.CLK(net758),
    .D(_1024_),
    .Q(\device.rxBuffer.buffer[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5037_ (.CLK(net759),
    .D(_1025_),
    .Q(\device.rxBuffer.buffer[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5038_ (.CLK(net760),
    .D(_1026_),
    .Q(\device.rxBuffer.buffer[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5039_ (.CLK(net761),
    .D(_1027_),
    .Q(\device.rxBuffer.buffer[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5040_ (.CLK(net762),
    .D(_1028_),
    .Q(\device.rxBuffer.buffer[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5041_ (.CLK(net763),
    .D(_1029_),
    .Q(\device.rxBuffer.buffer[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5042_ (.CLK(net764),
    .D(_1030_),
    .Q(\device.txBuffer.buffer[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5043_ (.CLK(net765),
    .D(_1031_),
    .Q(\device.txBuffer.buffer[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5044_ (.CLK(net766),
    .D(_1032_),
    .Q(\device.txBuffer.buffer[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5045_ (.CLK(net767),
    .D(_1033_),
    .Q(\device.txBuffer.buffer[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5046_ (.CLK(net768),
    .D(_1034_),
    .Q(\device.txBuffer.buffer[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5047_ (.CLK(net769),
    .D(_1035_),
    .Q(\device.txBuffer.buffer[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5048_ (.CLK(net770),
    .D(_1036_),
    .Q(\device.txBuffer.buffer[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5049_ (.CLK(net771),
    .D(_1037_),
    .Q(\device.txBuffer.buffer[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5050_ (.CLK(net772),
    .D(_1038_),
    .Q(\device.txBuffer.buffer[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5051_ (.CLK(net773),
    .D(_1039_),
    .Q(\device.txBuffer.buffer[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5052_ (.CLK(net774),
    .D(_1040_),
    .Q(\device.txBuffer.buffer[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5053_ (.CLK(net775),
    .D(_1041_),
    .Q(\device.txBuffer.buffer[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5054_ (.CLK(net776),
    .D(_1042_),
    .Q(\device.txBuffer.buffer[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5055_ (.CLK(net777),
    .D(_1043_),
    .Q(\device.txBuffer.buffer[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5056_ (.CLK(net778),
    .D(_1044_),
    .Q(\device.txBuffer.buffer[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5057_ (.CLK(net779),
    .D(_1045_),
    .Q(\device.txBuffer.buffer[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5058_ (.CLK(net780),
    .D(_1046_),
    .Q(\device.rxBuffer.buffer[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5059_ (.CLK(net781),
    .D(_1047_),
    .Q(\device.rxBuffer.buffer[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5060_ (.CLK(net782),
    .D(_1048_),
    .Q(\device.rxBuffer.buffer[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5061_ (.CLK(net783),
    .D(_1049_),
    .Q(\device.rxBuffer.buffer[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5062_ (.CLK(net784),
    .D(_1050_),
    .Q(\device.rxBuffer.buffer[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5063_ (.CLK(net785),
    .D(_1051_),
    .Q(\device.rxBuffer.buffer[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5064_ (.CLK(net786),
    .D(_1052_),
    .Q(\device.rxBuffer.buffer[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5065_ (.CLK(net787),
    .D(_1053_),
    .Q(\device.rxBuffer.buffer[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5066_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net2677),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5067_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net2656),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5068_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net2649),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5069_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net2663),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5070_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net1808),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5071_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net2670),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5072_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net1818),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5073_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net1837),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5074_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_1062_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[8] ));
 sky130_fd_sc_hd__dfxtp_1 _5075_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_1063_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[9] ));
 sky130_fd_sc_hd__dfxtp_1 _5076_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_1064_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[10] ));
 sky130_fd_sc_hd__dfxtp_1 _5077_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_1065_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[11] ));
 sky130_fd_sc_hd__dfxtp_1 _5078_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_1066_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[12] ));
 sky130_fd_sc_hd__dfxtp_1 _5079_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_1067_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[13] ));
 sky130_fd_sc_hd__dfxtp_1 _5080_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_1068_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[14] ));
 sky130_fd_sc_hd__dfxtp_1 _5081_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_1069_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[15] ));
 sky130_fd_sc_hd__dfxtp_1 _5082_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_1070_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[16] ));
 sky130_fd_sc_hd__dfxtp_1 _5083_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_1071_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[17] ));
 sky130_fd_sc_hd__dfxtp_1 _5084_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_1072_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[18] ));
 sky130_fd_sc_hd__dfxtp_1 _5085_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_1073_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[19] ));
 sky130_fd_sc_hd__dfxtp_1 _5086_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_1074_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[20] ));
 sky130_fd_sc_hd__dfxtp_1 _5087_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_1075_),
    .Q(\wbPeripheralBusInterface.dataRead_buffered[21] ));
 sky130_fd_sc_hd__dfxtp_1 _5088_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net1955),
    .Q(\wbPeripheralBusInterface.acknowledge ));
 sky130_fd_sc_hd__dfxtp_1 _5089_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net2852),
    .Q(\wbPeripheralBusInterface.currentAddress[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5090_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net2864),
    .Q(\wbPeripheralBusInterface.currentAddress[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5091_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net2756),
    .Q(\wbPeripheralBusInterface.currentAddress[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5092_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net2768),
    .Q(\wbPeripheralBusInterface.currentAddress[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5093_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net2780),
    .Q(\wbPeripheralBusInterface.currentAddress[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5094_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net2792),
    .Q(\wbPeripheralBusInterface.currentAddress[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5095_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net2804),
    .Q(\wbPeripheralBusInterface.currentAddress[8] ));
 sky130_fd_sc_hd__dfxtp_1 _5096_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net2816),
    .Q(\wbPeripheralBusInterface.currentAddress[9] ));
 sky130_fd_sc_hd__dfxtp_1 _5097_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net2828),
    .Q(\wbPeripheralBusInterface.currentAddress[10] ));
 sky130_fd_sc_hd__dfxtp_1 _5098_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net2840),
    .Q(\wbPeripheralBusInterface.currentAddress[11] ));
 sky130_fd_sc_hd__dfxtp_1 _5099_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net2876),
    .Q(\wbPeripheralBusInterface.currentAddress[12] ));
 sky130_fd_sc_hd__dfxtp_1 _5100_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net2900),
    .Q(\wbPeripheralBusInterface.currentAddress[13] ));
 sky130_fd_sc_hd__dfxtp_1 _5101_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net2888),
    .Q(\wbPeripheralBusInterface.currentAddress[14] ));
 sky130_fd_sc_hd__dfxtp_1 _5102_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_1090_),
    .Q(\wbPeripheralBusInterface.currentAddress[15] ));
 sky130_fd_sc_hd__dfxtp_1 _5103_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net1584),
    .Q(\wbPeripheralBusInterface.currentAddress[16] ));
 sky130_fd_sc_hd__dfxtp_1 _5104_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_1092_),
    .Q(\wbPeripheralBusInterface.currentAddress[17] ));
 sky130_fd_sc_hd__dfxtp_1 _5105_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net1592),
    .Q(\wbPeripheralBusInterface.currentAddress[18] ));
 sky130_fd_sc_hd__dfxtp_1 _5106_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_1094_),
    .Q(\wbPeripheralBusInterface.currentAddress[19] ));
 sky130_fd_sc_hd__dfxtp_1 _5107_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(net1603),
    .Q(\wbPeripheralBusInterface.currentAddress[20] ));
 sky130_fd_sc_hd__dfxtp_1 _5108_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_1096_),
    .Q(\wbPeripheralBusInterface.currentAddress[21] ));
 sky130_fd_sc_hd__dfxtp_1 _5109_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_1097_),
    .Q(\wbPeripheralBusInterface.currentAddress[22] ));
 sky130_fd_sc_hd__dfxtp_1 _5110_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_1098_),
    .Q(\wbPeripheralBusInterface.currentAddress[23] ));
 sky130_fd_sc_hd__dfxtp_2 _5111_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net3248),
    .Q(\wbPeripheralBusInterface.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5112_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net3334),
    .Q(\wbPeripheralBusInterface.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5113_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net2733),
    .Q(\wbAddressExtension.acknowledge ));
 sky130_fd_sc_hd__dfxtp_1 _5114_ (.CLK(net788),
    .D(_1102_),
    .Q(\device.rxBuffer.buffer[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5115_ (.CLK(net789),
    .D(_1103_),
    .Q(\device.rxBuffer.buffer[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5116_ (.CLK(net790),
    .D(_1104_),
    .Q(\device.rxBuffer.buffer[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5117_ (.CLK(net791),
    .D(_1105_),
    .Q(\device.rxBuffer.buffer[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5118_ (.CLK(net792),
    .D(_1106_),
    .Q(\device.rxBuffer.buffer[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5119_ (.CLK(net793),
    .D(_1107_),
    .Q(\device.rxBuffer.buffer[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5120_ (.CLK(net794),
    .D(_1108_),
    .Q(\device.rxBuffer.buffer[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5121_ (.CLK(net795),
    .D(_1109_),
    .Q(\device.rxBuffer.buffer[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5122_ (.CLK(net796),
    .D(_1110_),
    .Q(\device.rxBuffer.buffer[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5123_ (.CLK(net797),
    .D(_1111_),
    .Q(\device.rxBuffer.buffer[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5124_ (.CLK(net798),
    .D(_1112_),
    .Q(\device.rxBuffer.buffer[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5125_ (.CLK(net799),
    .D(_1113_),
    .Q(\device.rxBuffer.buffer[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5126_ (.CLK(net800),
    .D(_1114_),
    .Q(\device.rxBuffer.buffer[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5127_ (.CLK(net801),
    .D(_1115_),
    .Q(\device.rxBuffer.buffer[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5128_ (.CLK(net802),
    .D(_1116_),
    .Q(\device.rxBuffer.buffer[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5129_ (.CLK(net803),
    .D(_1117_),
    .Q(\device.rxBuffer.buffer[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5130_ (.CLK(net804),
    .D(_1118_),
    .Q(\device.rxBuffer.buffer[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5131_ (.CLK(net805),
    .D(_1119_),
    .Q(\device.rxBuffer.buffer[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5132_ (.CLK(net806),
    .D(_1120_),
    .Q(\device.rxBuffer.buffer[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5133_ (.CLK(net807),
    .D(_1121_),
    .Q(\device.rxBuffer.buffer[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5134_ (.CLK(net808),
    .D(_1122_),
    .Q(\device.rxBuffer.buffer[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5135_ (.CLK(net809),
    .D(_1123_),
    .Q(\device.rxBuffer.buffer[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5136_ (.CLK(net810),
    .D(_1124_),
    .Q(\device.rxBuffer.buffer[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5137_ (.CLK(net811),
    .D(_1125_),
    .Q(\device.rxBuffer.buffer[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5138_ (.CLK(net812),
    .D(_1126_),
    .Q(\device.rxBuffer.buffer[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5139_ (.CLK(net813),
    .D(_1127_),
    .Q(\device.rxBuffer.buffer[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5140_ (.CLK(net814),
    .D(_1128_),
    .Q(\device.rxBuffer.buffer[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5141_ (.CLK(net815),
    .D(_1129_),
    .Q(\device.rxBuffer.buffer[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5142_ (.CLK(net816),
    .D(_1130_),
    .Q(\device.rxBuffer.buffer[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5143_ (.CLK(net817),
    .D(_1131_),
    .Q(\device.rxBuffer.buffer[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5144_ (.CLK(net818),
    .D(_1132_),
    .Q(\device.rxBuffer.buffer[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5145_ (.CLK(net819),
    .D(_1133_),
    .Q(\device.rxBuffer.buffer[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5146_ (.CLK(net820),
    .D(_1134_),
    .Q(\device.rxBuffer.buffer[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5147_ (.CLK(net821),
    .D(_1135_),
    .Q(\device.rxBuffer.buffer[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5148_ (.CLK(net822),
    .D(_1136_),
    .Q(\device.rxBuffer.buffer[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5149_ (.CLK(net823),
    .D(_1137_),
    .Q(\device.rxBuffer.buffer[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5150_ (.CLK(net824),
    .D(_1138_),
    .Q(\device.rxBuffer.buffer[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5151_ (.CLK(net825),
    .D(_1139_),
    .Q(\device.rxBuffer.buffer[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5152_ (.CLK(net826),
    .D(_1140_),
    .Q(\device.rxBuffer.buffer[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5153_ (.CLK(net827),
    .D(_1141_),
    .Q(\device.rxBuffer.buffer[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5154_ (.CLK(net828),
    .D(_1142_),
    .Q(\device.rxBuffer.buffer[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5155_ (.CLK(net829),
    .D(_1143_),
    .Q(\device.rxBuffer.buffer[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5156_ (.CLK(net830),
    .D(_1144_),
    .Q(\device.rxBuffer.buffer[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5157_ (.CLK(net831),
    .D(_1145_),
    .Q(\device.rxBuffer.buffer[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5158_ (.CLK(net832),
    .D(_1146_),
    .Q(\device.rxBuffer.buffer[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5159_ (.CLK(net833),
    .D(_1147_),
    .Q(\device.rxBuffer.buffer[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5160_ (.CLK(net834),
    .D(_1148_),
    .Q(\device.rxBuffer.buffer[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5161_ (.CLK(net835),
    .D(_1149_),
    .Q(\device.rxBuffer.buffer[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5162_ (.CLK(net836),
    .D(_1150_),
    .Q(\device.rxBuffer.buffer[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5163_ (.CLK(net837),
    .D(_1151_),
    .Q(\device.rxBuffer.buffer[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5164_ (.CLK(net838),
    .D(_1152_),
    .Q(\device.rxBuffer.buffer[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5165_ (.CLK(net839),
    .D(_1153_),
    .Q(\device.rxBuffer.buffer[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5166_ (.CLK(net840),
    .D(_1154_),
    .Q(\device.rxBuffer.buffer[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5167_ (.CLK(net841),
    .D(_1155_),
    .Q(\device.rxBuffer.buffer[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5168_ (.CLK(net842),
    .D(_1156_),
    .Q(\device.rxBuffer.buffer[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5169_ (.CLK(net843),
    .D(_1157_),
    .Q(\device.rxBuffer.buffer[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5170_ (.CLK(net844),
    .D(_1158_),
    .Q(\device.rxBuffer.buffer[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5171_ (.CLK(net845),
    .D(_1159_),
    .Q(\device.rxBuffer.buffer[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5172_ (.CLK(net846),
    .D(_1160_),
    .Q(\device.rxBuffer.buffer[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5173_ (.CLK(net847),
    .D(_1161_),
    .Q(\device.rxBuffer.buffer[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5174_ (.CLK(net848),
    .D(_1162_),
    .Q(\device.rxBuffer.buffer[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5175_ (.CLK(net849),
    .D(_1163_),
    .Q(\device.rxBuffer.buffer[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5176_ (.CLK(net850),
    .D(_1164_),
    .Q(\device.rxBuffer.buffer[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5177_ (.CLK(net851),
    .D(_1165_),
    .Q(\device.rxBuffer.buffer[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5178_ (.CLK(net852),
    .D(_1166_),
    .Q(\device.rxBuffer.buffer[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5179_ (.CLK(net853),
    .D(_1167_),
    .Q(\device.rxBuffer.buffer[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5180_ (.CLK(net854),
    .D(_1168_),
    .Q(\device.rxBuffer.buffer[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5181_ (.CLK(net855),
    .D(_1169_),
    .Q(\device.rxBuffer.buffer[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5182_ (.CLK(net856),
    .D(_1170_),
    .Q(\device.rxBuffer.buffer[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5183_ (.CLK(net857),
    .D(_1171_),
    .Q(\device.rxBuffer.buffer[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5184_ (.CLK(net858),
    .D(_1172_),
    .Q(\device.rxBuffer.buffer[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5185_ (.CLK(net859),
    .D(_1173_),
    .Q(\device.rxBuffer.buffer[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5186_ (.CLK(net860),
    .D(_1174_),
    .Q(\device.rxBuffer.buffer[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5187_ (.CLK(net861),
    .D(_1175_),
    .Q(\device.rxBuffer.buffer[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5188_ (.CLK(net862),
    .D(_1176_),
    .Q(\device.rxBuffer.buffer[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5189_ (.CLK(net863),
    .D(_1177_),
    .Q(\device.rxBuffer.buffer[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5190_ (.CLK(net864),
    .D(_1178_),
    .Q(\device.rxBuffer.buffer[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5191_ (.CLK(net865),
    .D(_1179_),
    .Q(\device.rxBuffer.buffer[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5192_ (.CLK(net866),
    .D(_1180_),
    .Q(\device.rxBuffer.buffer[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5193_ (.CLK(net867),
    .D(_1181_),
    .Q(\device.rxBuffer.buffer[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5194_ (.CLK(net868),
    .D(_1182_),
    .Q(\device.rxBuffer.buffer[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5195_ (.CLK(net869),
    .D(_1183_),
    .Q(\device.rxBuffer.buffer[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5196_ (.CLK(net870),
    .D(_1184_),
    .Q(\device.rxBuffer.buffer[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5197_ (.CLK(net871),
    .D(_1185_),
    .Q(\device.rxBuffer.buffer[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5198_ (.CLK(net872),
    .D(_1186_),
    .Q(\device.rxBuffer.buffer[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5199_ (.CLK(net873),
    .D(_1187_),
    .Q(\device.rxBuffer.buffer[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5200_ (.CLK(net874),
    .D(_1188_),
    .Q(\device.rxBuffer.buffer[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5201_ (.CLK(net875),
    .D(_1189_),
    .Q(\device.rxBuffer.buffer[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5202_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_1190_),
    .Q(\device.rxRegister.baseReadData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5203_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_1191_),
    .Q(\device.rxRegister.baseReadData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5204_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net1669),
    .Q(\device.rxRegister.baseReadData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5205_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net1676),
    .Q(\device.rxRegister.baseReadData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5206_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_1194_),
    .Q(\device.rxRegister.baseReadData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5207_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_1195_),
    .Q(\device.rxRegister.baseReadData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5208_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_1196_),
    .Q(\device.rxRegister.baseReadData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5209_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_1197_),
    .Q(\device.rxRegister.baseReadData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5210_ (.CLK(net876),
    .D(_1198_),
    .Q(\device.rxBuffer.buffer[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5211_ (.CLK(net877),
    .D(_1199_),
    .Q(\device.rxBuffer.buffer[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5212_ (.CLK(net878),
    .D(_1200_),
    .Q(\device.rxBuffer.buffer[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5213_ (.CLK(net879),
    .D(_1201_),
    .Q(\device.rxBuffer.buffer[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5214_ (.CLK(net880),
    .D(_1202_),
    .Q(\device.rxBuffer.buffer[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5215_ (.CLK(net881),
    .D(_1203_),
    .Q(\device.rxBuffer.buffer[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5216_ (.CLK(net882),
    .D(_1204_),
    .Q(\device.rxBuffer.buffer[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5217_ (.CLK(net883),
    .D(_1205_),
    .Q(\device.rxBuffer.buffer[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5218_ (.CLK(net884),
    .D(_1206_),
    .Q(\device.rxBuffer.buffer[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5219_ (.CLK(net885),
    .D(_1207_),
    .Q(\device.rxBuffer.buffer[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5220_ (.CLK(net886),
    .D(_1208_),
    .Q(\device.rxBuffer.buffer[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5221_ (.CLK(net887),
    .D(_1209_),
    .Q(\device.rxBuffer.buffer[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5222_ (.CLK(net888),
    .D(_1210_),
    .Q(\device.rxBuffer.buffer[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5223_ (.CLK(net889),
    .D(_1211_),
    .Q(\device.rxBuffer.buffer[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5224_ (.CLK(net890),
    .D(_1212_),
    .Q(\device.rxBuffer.buffer[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5225_ (.CLK(net891),
    .D(_1213_),
    .Q(\device.rxBuffer.buffer[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5226_ (.CLK(net892),
    .D(_1214_),
    .Q(\device.rxBuffer.buffer[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5227_ (.CLK(net893),
    .D(_1215_),
    .Q(\device.rxBuffer.buffer[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5228_ (.CLK(net894),
    .D(_1216_),
    .Q(\device.rxBuffer.buffer[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5229_ (.CLK(net895),
    .D(_1217_),
    .Q(\device.rxBuffer.buffer[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5230_ (.CLK(net896),
    .D(_1218_),
    .Q(\device.rxBuffer.buffer[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5231_ (.CLK(net897),
    .D(_1219_),
    .Q(\device.rxBuffer.buffer[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5232_ (.CLK(net898),
    .D(_1220_),
    .Q(\device.rxBuffer.buffer[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5233_ (.CLK(net899),
    .D(_1221_),
    .Q(\device.rxBuffer.buffer[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5234_ (.CLK(net900),
    .D(_1222_),
    .Q(\device.rxBuffer.buffer[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5235_ (.CLK(net901),
    .D(_1223_),
    .Q(\device.rxBuffer.buffer[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5236_ (.CLK(net902),
    .D(_1224_),
    .Q(\device.rxBuffer.buffer[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5237_ (.CLK(net903),
    .D(_1225_),
    .Q(\device.rxBuffer.buffer[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5238_ (.CLK(net904),
    .D(_1226_),
    .Q(\device.rxBuffer.buffer[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5239_ (.CLK(net905),
    .D(_1227_),
    .Q(\device.rxBuffer.buffer[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5240_ (.CLK(net906),
    .D(_1228_),
    .Q(\device.rxBuffer.buffer[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5241_ (.CLK(net907),
    .D(_1229_),
    .Q(\device.rxBuffer.buffer[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5242_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_1230_),
    .Q(\wbAddressExtension.currentAddress[8] ));
 sky130_fd_sc_hd__dfxtp_1 _5243_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_1231_),
    .Q(\wbAddressExtension.currentAddress[9] ));
 sky130_fd_sc_hd__dfxtp_1 _5244_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_1232_),
    .Q(\wbAddressExtension.currentAddress[10] ));
 sky130_fd_sc_hd__dfxtp_1 _5245_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_1233_),
    .Q(\wbAddressExtension.currentAddress[11] ));
 sky130_fd_sc_hd__dfxtp_1 _5246_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(net1443),
    .Q(\wbAddressExtension.currentAddress[12] ));
 sky130_fd_sc_hd__dfxtp_1 _5247_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_1235_),
    .Q(\wbAddressExtension.currentAddress[13] ));
 sky130_fd_sc_hd__dfxtp_1 _5248_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(net1428),
    .Q(\wbAddressExtension.currentAddress[14] ));
 sky130_fd_sc_hd__dfxtp_2 _5249_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_1237_),
    .Q(\wbAddressExtension.currentAddress[15] ));
 sky130_fd_sc_hd__dfxtp_2 _5250_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_1238_),
    .Q(\wbAddressExtension.currentAddress[16] ));
 sky130_fd_sc_hd__dfxtp_2 _5251_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net1402),
    .Q(\wbAddressExtension.currentAddress[17] ));
 sky130_fd_sc_hd__dfxtp_2 _5252_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net1391),
    .Q(\wbAddressExtension.currentAddress[18] ));
 sky130_fd_sc_hd__dfxtp_2 _5253_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_1241_),
    .Q(\wbAddressExtension.currentAddress[19] ));
 sky130_fd_sc_hd__dfxtp_2 _5254_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_1242_),
    .Q(\wbAddressExtension.currentAddress[20] ));
 sky130_fd_sc_hd__dfxtp_2 _5255_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_1243_),
    .Q(\wbAddressExtension.currentAddress[21] ));
 sky130_fd_sc_hd__dfxtp_2 _5256_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_1244_),
    .Q(\wbAddressExtension.currentAddress[22] ));
 sky130_fd_sc_hd__dfxtp_2 _5257_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_1245_),
    .Q(\wbAddressExtension.currentAddress[23] ));
 sky130_fd_sc_hd__dfxtp_2 _5258_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_1246_),
    .Q(\wbAddressExtension.currentAddress[24] ));
 sky130_fd_sc_hd__dfxtp_2 _5259_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(net1514),
    .Q(\wbAddressExtension.currentAddress[25] ));
 sky130_fd_sc_hd__dfxtp_2 _5260_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(net1494),
    .Q(\wbAddressExtension.currentAddress[26] ));
 sky130_fd_sc_hd__dfxtp_2 _5261_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(net1501),
    .Q(\wbAddressExtension.currentAddress[27] ));
 sky130_fd_sc_hd__dfxtp_1 _5262_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_1250_),
    .Q(\wbAddressExtension.currentAddress[28] ));
 sky130_fd_sc_hd__dfxtp_1 _5263_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_1251_),
    .Q(\wbAddressExtension.currentAddress[29] ));
 sky130_fd_sc_hd__dfxtp_1 _5264_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_1252_),
    .Q(\wbAddressExtension.currentAddress[30] ));
 sky130_fd_sc_hd__dfxtp_1 _5265_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_1253_),
    .Q(\wbAddressExtension.currentAddress[31] ));
 sky130_fd_sc_hd__dfxtp_1 _5266_ (.CLK(net908),
    .D(_1254_),
    .Q(\device.txBuffer.buffer[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5267_ (.CLK(net909),
    .D(_1255_),
    .Q(\device.txBuffer.buffer[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5268_ (.CLK(net910),
    .D(_1256_),
    .Q(\device.txBuffer.buffer[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5269_ (.CLK(net911),
    .D(_1257_),
    .Q(\device.txBuffer.buffer[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5270_ (.CLK(net912),
    .D(_1258_),
    .Q(\device.txBuffer.buffer[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5271_ (.CLK(net913),
    .D(_1259_),
    .Q(\device.txBuffer.buffer[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5272_ (.CLK(net914),
    .D(_1260_),
    .Q(\device.txBuffer.buffer[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5273_ (.CLK(net915),
    .D(_1261_),
    .Q(\device.txBuffer.buffer[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5274_ (.CLK(net916),
    .D(_1262_),
    .Q(\device.txBuffer.buffer[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5275_ (.CLK(net917),
    .D(_1263_),
    .Q(\device.txBuffer.buffer[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5276_ (.CLK(net918),
    .D(_1264_),
    .Q(\device.txBuffer.buffer[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5277_ (.CLK(net919),
    .D(_1265_),
    .Q(\device.txBuffer.buffer[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5278_ (.CLK(net920),
    .D(_1266_),
    .Q(\device.txBuffer.buffer[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5279_ (.CLK(net921),
    .D(_1267_),
    .Q(\device.txBuffer.buffer[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5280_ (.CLK(net922),
    .D(_1268_),
    .Q(\device.txBuffer.buffer[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5281_ (.CLK(net923),
    .D(_1269_),
    .Q(\device.txBuffer.buffer[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5282_ (.CLK(net924),
    .D(_1270_),
    .Q(\device.txBuffer.buffer[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5283_ (.CLK(net925),
    .D(_1271_),
    .Q(\device.txBuffer.buffer[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5284_ (.CLK(net926),
    .D(_1272_),
    .Q(\device.txBuffer.buffer[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5285_ (.CLK(net927),
    .D(_1273_),
    .Q(\device.txBuffer.buffer[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5286_ (.CLK(net928),
    .D(_1274_),
    .Q(\device.txBuffer.buffer[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5287_ (.CLK(net929),
    .D(_1275_),
    .Q(\device.txBuffer.buffer[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5288_ (.CLK(net930),
    .D(_1276_),
    .Q(\device.txBuffer.buffer[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5289_ (.CLK(net931),
    .D(_1277_),
    .Q(\device.txBuffer.buffer[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5290_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net1292),
    .Q(\wbPeripheralBusInterface.currentByteSelect[0] ));
 sky130_fd_sc_hd__dfxtp_2 _5291_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net1316),
    .Q(\wbPeripheralBusInterface.currentByteSelect[1] ));
 sky130_fd_sc_hd__dfxtp_2 _5292_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net1334),
    .Q(\wbPeripheralBusInterface.currentByteSelect[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5293_ (.CLK(net932),
    .D(_1281_),
    .Q(\device.txBuffer.buffer[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5294_ (.CLK(net933),
    .D(_1282_),
    .Q(\device.txBuffer.buffer[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5295_ (.CLK(net934),
    .D(_1283_),
    .Q(\device.txBuffer.buffer[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5296_ (.CLK(net935),
    .D(_1284_),
    .Q(\device.txBuffer.buffer[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5297_ (.CLK(net936),
    .D(_1285_),
    .Q(\device.txBuffer.buffer[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5298_ (.CLK(net937),
    .D(_1286_),
    .Q(\device.txBuffer.buffer[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5299_ (.CLK(net938),
    .D(_1287_),
    .Q(\device.txBuffer.buffer[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5300_ (.CLK(net939),
    .D(_1288_),
    .Q(\device.txBuffer.buffer[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5301_ (.CLK(net940),
    .D(_1289_),
    .Q(\device.txBuffer.buffer[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5302_ (.CLK(net941),
    .D(_1290_),
    .Q(\device.txBuffer.buffer[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5303_ (.CLK(net942),
    .D(_1291_),
    .Q(\device.txBuffer.buffer[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5304_ (.CLK(net943),
    .D(_1292_),
    .Q(\device.txBuffer.buffer[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5305_ (.CLK(net944),
    .D(_1293_),
    .Q(\device.txBuffer.buffer[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5306_ (.CLK(net945),
    .D(_1294_),
    .Q(\device.txBuffer.buffer[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5307_ (.CLK(net946),
    .D(_1295_),
    .Q(\device.txBuffer.buffer[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5308_ (.CLK(net947),
    .D(_1296_),
    .Q(\device.txBuffer.buffer[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5309_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_1297_),
    .Q(\device.uartRx.newData ));
 sky130_fd_sc_hd__dfxtp_1 _5310_ (.CLK(net948),
    .D(_1298_),
    .Q(\device.rxBuffer.buffer[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5311_ (.CLK(net949),
    .D(_1299_),
    .Q(\device.rxBuffer.buffer[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5312_ (.CLK(net950),
    .D(_1300_),
    .Q(\device.rxBuffer.buffer[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5313_ (.CLK(net951),
    .D(_1301_),
    .Q(\device.rxBuffer.buffer[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5314_ (.CLK(net952),
    .D(_1302_),
    .Q(\device.rxBuffer.buffer[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5315_ (.CLK(net953),
    .D(_1303_),
    .Q(\device.rxBuffer.buffer[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5316_ (.CLK(net954),
    .D(_1304_),
    .Q(\device.rxBuffer.buffer[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5317_ (.CLK(net955),
    .D(_1305_),
    .Q(\device.rxBuffer.buffer[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5318_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(net3759),
    .Q(\device.rxBuffer.dataIn_buffered[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5319_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(net3772),
    .Q(\device.rxBuffer.dataIn_buffered[1] ));
 sky130_fd_sc_hd__dfxtp_4 _5320_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(net3785),
    .Q(\device.rxBuffer.dataIn_buffered[2] ));
 sky130_fd_sc_hd__dfxtp_4 _5321_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(net3824),
    .Q(\device.rxBuffer.dataIn_buffered[3] ));
 sky130_fd_sc_hd__dfxtp_2 _5322_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(net3811),
    .Q(\device.rxBuffer.dataIn_buffered[4] ));
 sky130_fd_sc_hd__dfxtp_4 _5323_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(net3798),
    .Q(\device.rxBuffer.dataIn_buffered[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5324_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(net3502),
    .Q(\device.rxBuffer.dataIn_buffered[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5325_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(net3514),
    .Q(\device.rxBuffer.dataIn_buffered[7] ));
 sky130_fd_sc_hd__dfxtp_2 _5326_ (.CLK(net956),
    .D(_1314_),
    .Q(\device.txBuffer.startPointer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5327_ (.CLK(net957),
    .D(_1315_),
    .Q(\device.txBuffer.startPointer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5328_ (.CLK(net958),
    .D(_1316_),
    .Q(\device.txBuffer.startPointer[2] ));
 sky130_fd_sc_hd__dfxtp_2 _5329_ (.CLK(net959),
    .D(_1317_),
    .Q(\device.txBuffer.startPointer[3] ));
 sky130_fd_sc_hd__dfxtp_4 _5330_ (.CLK(net960),
    .D(_1318_),
    .Q(\device.txBuffer.startPointer[4] ));
 sky130_fd_sc_hd__dfxtp_2 _5331_ (.CLK(net961),
    .D(_1319_),
    .Q(\device.txBuffer.endPointer[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5332_ (.CLK(net962),
    .D(_1320_),
    .Q(\device.txBuffer.endPointer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5333_ (.CLK(net963),
    .D(_1321_),
    .Q(\device.txBuffer.endPointer[2] ));
 sky130_fd_sc_hd__dfxtp_4 _5334_ (.CLK(net964),
    .D(_1322_),
    .Q(\device.txBuffer.endPointer[3] ));
 sky130_fd_sc_hd__dfxtp_4 _5335_ (.CLK(net965),
    .D(_1323_),
    .Q(\device.txBuffer.endPointer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5336_ (.CLK(net966),
    .D(_1324_),
    .Q(\device.txBuffer.lastWriteLostData ));
 sky130_fd_sc_hd__dfxtp_1 _5337_ (.CLK(net967),
    .D(_1325_),
    .Q(\device.txBuffer.dataOut[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5338_ (.CLK(net968),
    .D(_1326_),
    .Q(\device.txBuffer.dataOut[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5339_ (.CLK(net969),
    .D(_1327_),
    .Q(\device.txBuffer.dataOut[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5340_ (.CLK(net970),
    .D(_1328_),
    .Q(\device.txBuffer.dataOut[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5341_ (.CLK(net971),
    .D(_1329_),
    .Q(\device.txBuffer.dataOut[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5342_ (.CLK(net972),
    .D(_1330_),
    .Q(\device.txBuffer.dataOut[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5343_ (.CLK(net973),
    .D(_1331_),
    .Q(\device.txBuffer.dataOut[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5344_ (.CLK(net974),
    .D(_1332_),
    .Q(\device.txBuffer.dataOut[7] ));
 sky130_fd_sc_hd__dfxtp_4 _5345_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net3305),
    .Q(\device.txBuffer.we_buffered ));
 sky130_fd_sc_hd__dfxtp_1 _5346_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(net3351),
    .Q(\device.txBuffer.oe_buffered ));
 sky130_fd_sc_hd__dfxtp_1 _5347_ (.CLK(net975),
    .D(_1335_),
    .Q(\device.rxBuffer.buffer[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5348_ (.CLK(net976),
    .D(_1336_),
    .Q(\device.rxBuffer.buffer[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5349_ (.CLK(net977),
    .D(_1337_),
    .Q(\device.rxBuffer.buffer[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5350_ (.CLK(net978),
    .D(_1338_),
    .Q(\device.rxBuffer.buffer[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5351_ (.CLK(net979),
    .D(_1339_),
    .Q(\device.rxBuffer.buffer[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5352_ (.CLK(net980),
    .D(_0550_),
    .Q(\device.rxBuffer.buffer[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5353_ (.CLK(net981),
    .D(_0551_),
    .Q(\device.rxBuffer.buffer[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5354_ (.CLK(net982),
    .D(_0552_),
    .Q(\device.rxBuffer.buffer[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5355_ (.CLK(net983),
    .D(_0553_),
    .Q(\device.rxBuffer.buffer[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5356_ (.CLK(net984),
    .D(_0554_),
    .Q(\device.rxBuffer.buffer[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5357_ (.CLK(net985),
    .D(_0555_),
    .Q(\device.rxBuffer.buffer[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5358_ (.CLK(net986),
    .D(_0556_),
    .Q(\device.rxBuffer.buffer[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5359_ (.CLK(net987),
    .D(_0557_),
    .Q(\device.rxBuffer.buffer[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5360_ (.CLK(net988),
    .D(_0558_),
    .Q(\device.rxBuffer.buffer[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5361_ (.CLK(net989),
    .D(_0559_),
    .Q(\device.rxBuffer.buffer[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5362_ (.CLK(net990),
    .D(_0560_),
    .Q(\device.rxBuffer.buffer[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5363_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net1686),
    .Q(\device.rxDataAvailableBuffered ));
 sky130_fd_sc_hd__dfxtp_2 _5364_ (.CLK(net991),
    .D(_0562_),
    .Q(\device.rxBuffer.startPointer[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5365_ (.CLK(net992),
    .D(_0563_),
    .Q(\device.rxBuffer.startPointer[1] ));
 sky130_fd_sc_hd__dfxtp_4 _5366_ (.CLK(net993),
    .D(_0564_),
    .Q(\device.rxBuffer.startPointer[2] ));
 sky130_fd_sc_hd__dfxtp_2 _5367_ (.CLK(net994),
    .D(_0565_),
    .Q(\device.rxBuffer.startPointer[3] ));
 sky130_fd_sc_hd__dfxtp_4 _5368_ (.CLK(net995),
    .D(_0566_),
    .Q(\device.rxBuffer.startPointer[4] ));
 sky130_fd_sc_hd__dfxtp_4 _5369_ (.CLK(net996),
    .D(_0567_),
    .Q(\device.rxBuffer.endPointer[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5370_ (.CLK(net997),
    .D(_0568_),
    .Q(\device.rxBuffer.endPointer[1] ));
 sky130_fd_sc_hd__dfxtp_2 _5371_ (.CLK(net998),
    .D(_0569_),
    .Q(\device.rxBuffer.endPointer[2] ));
 sky130_fd_sc_hd__dfxtp_2 _5372_ (.CLK(net999),
    .D(_0570_),
    .Q(\device.rxBuffer.endPointer[3] ));
 sky130_fd_sc_hd__dfxtp_4 _5373_ (.CLK(net1000),
    .D(_0571_),
    .Q(\device.rxBuffer.endPointer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5374_ (.CLK(net1001),
    .D(_0572_),
    .Q(\device.rxBuffer.lastWriteLostData ));
 sky130_fd_sc_hd__dfxtp_1 _5375_ (.CLK(net1002),
    .D(_0573_),
    .Q(\device.rxBuffer.dataOut[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5376_ (.CLK(net1003),
    .D(_0574_),
    .Q(\device.rxBuffer.dataOut[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5377_ (.CLK(net1004),
    .D(_0575_),
    .Q(\device.rxBuffer.dataOut[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5378_ (.CLK(net1005),
    .D(_0576_),
    .Q(\device.rxBuffer.dataOut[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5379_ (.CLK(net1006),
    .D(_0577_),
    .Q(\device.rxBuffer.dataOut[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5380_ (.CLK(net1007),
    .D(_0578_),
    .Q(\device.rxBuffer.dataOut[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5381_ (.CLK(net1008),
    .D(_0579_),
    .Q(\device.rxBuffer.dataOut[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5382_ (.CLK(net1009),
    .D(_0580_),
    .Q(\device.rxBuffer.dataOut[7] ));
 sky130_fd_sc_hd__dfxtp_4 _5383_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net3568),
    .Q(\device.rxBuffer.we_buffered ));
 sky130_fd_sc_hd__dfxtp_1 _5384_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net2686),
    .Q(\device.rxBuffer.oe_buffered ));
 sky130_fd_sc_hd__dfxtp_1 _5385_ (.CLK(net1010),
    .D(_0583_),
    .Q(\device.txBuffer.buffer[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5386_ (.CLK(net1011),
    .D(_0584_),
    .Q(\device.txBuffer.buffer[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5387_ (.CLK(net1012),
    .D(_0585_),
    .Q(\device.txBuffer.buffer[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5388_ (.CLK(net1013),
    .D(_0586_),
    .Q(\device.txBuffer.buffer[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5389_ (.CLK(net1014),
    .D(_0587_),
    .Q(\device.txBuffer.buffer[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5390_ (.CLK(net1015),
    .D(_0588_),
    .Q(\device.txBuffer.buffer[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5391_ (.CLK(net1016),
    .D(_0589_),
    .Q(\device.txBuffer.buffer[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5392_ (.CLK(net1017),
    .D(_0590_),
    .Q(\device.txBuffer.buffer[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5393_ (.CLK(net1018),
    .D(_0591_),
    .Q(\device.rxBuffer.buffer[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5394_ (.CLK(net1019),
    .D(_0592_),
    .Q(\device.rxBuffer.buffer[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5395_ (.CLK(net1020),
    .D(_0593_),
    .Q(\device.rxBuffer.buffer[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5396_ (.CLK(net1021),
    .D(_0594_),
    .Q(\device.rxBuffer.buffer[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5397_ (.CLK(net1022),
    .D(_0595_),
    .Q(\device.rxBuffer.buffer[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5398_ (.CLK(net1023),
    .D(_0596_),
    .Q(\device.rxBuffer.buffer[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5399_ (.CLK(net1024),
    .D(_0597_),
    .Q(\device.rxBuffer.buffer[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5400_ (.CLK(net1025),
    .D(_0598_),
    .Q(\device.rxBuffer.buffer[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5401_ (.CLK(net1026),
    .D(_0599_),
    .Q(\device.rxBuffer.buffer[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5402_ (.CLK(net1027),
    .D(_0600_),
    .Q(\device.rxBuffer.buffer[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5403_ (.CLK(net1028),
    .D(_0601_),
    .Q(\device.rxBuffer.buffer[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5404_ (.CLK(net1029),
    .D(_0602_),
    .Q(\device.rxBuffer.buffer[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5405_ (.CLK(net1030),
    .D(_0603_),
    .Q(\device.rxBuffer.buffer[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5406_ (.CLK(net1031),
    .D(_0604_),
    .Q(\device.rxBuffer.buffer[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5407_ (.CLK(net1032),
    .D(_0605_),
    .Q(\device.rxBuffer.buffer[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5408_ (.CLK(net1033),
    .D(_0606_),
    .Q(\device.rxBuffer.buffer[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5409_ (.CLK(net1034),
    .D(_0607_),
    .Q(\device.txBuffer.buffer[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5410_ (.CLK(net1035),
    .D(_0608_),
    .Q(\device.txBuffer.buffer[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5411_ (.CLK(net1036),
    .D(_0609_),
    .Q(\device.txBuffer.buffer[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5412_ (.CLK(net1037),
    .D(_0610_),
    .Q(\device.txBuffer.buffer[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5413_ (.CLK(net1038),
    .D(_0611_),
    .Q(\device.txBuffer.buffer[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5414_ (.CLK(net1039),
    .D(_0612_),
    .Q(\device.txBuffer.buffer[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5415_ (.CLK(net1040),
    .D(_0613_),
    .Q(\device.txBuffer.buffer[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5416_ (.CLK(net1041),
    .D(_0614_),
    .Q(\device.txBuffer.buffer[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5417_ (.CLK(net1042),
    .D(_0615_),
    .Q(\device.txBuffer.buffer[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5418_ (.CLK(net1043),
    .D(_0616_),
    .Q(\device.txBuffer.buffer[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5419_ (.CLK(net1044),
    .D(_0617_),
    .Q(\device.txBuffer.buffer[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5420_ (.CLK(net1045),
    .D(_0618_),
    .Q(\device.txBuffer.buffer[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5421_ (.CLK(net1046),
    .D(_0619_),
    .Q(\device.txBuffer.buffer[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5422_ (.CLK(net1047),
    .D(_0620_),
    .Q(\device.txBuffer.buffer[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5423_ (.CLK(net1048),
    .D(_0621_),
    .Q(\device.txBuffer.buffer[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5424_ (.CLK(net1049),
    .D(_0622_),
    .Q(\device.txBuffer.buffer[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5425_ (.CLK(net1050),
    .D(_0623_),
    .Q(\device.rxBuffer.buffer[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5426_ (.CLK(net1051),
    .D(_0624_),
    .Q(\device.rxBuffer.buffer[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5427_ (.CLK(net1052),
    .D(_0625_),
    .Q(\device.rxBuffer.buffer[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5428_ (.CLK(net1053),
    .D(_0626_),
    .Q(\device.rxBuffer.buffer[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5429_ (.CLK(net1054),
    .D(_0627_),
    .Q(\device.rxBuffer.buffer[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5430_ (.CLK(net1055),
    .D(_0628_),
    .Q(\device.rxBuffer.buffer[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5431_ (.CLK(net1056),
    .D(_0629_),
    .Q(\device.rxBuffer.buffer[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5432_ (.CLK(net1057),
    .D(_0630_),
    .Q(\device.rxBuffer.buffer[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5433_ (.CLK(net1058),
    .D(_0631_),
    .Q(\device.rxBuffer.buffer[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5434_ (.CLK(net1059),
    .D(_0632_),
    .Q(\device.rxBuffer.buffer[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5435_ (.CLK(net1060),
    .D(_0633_),
    .Q(\device.rxBuffer.buffer[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5436_ (.CLK(net1061),
    .D(_0634_),
    .Q(\device.rxBuffer.buffer[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5437_ (.CLK(net1062),
    .D(_0635_),
    .Q(\device.rxBuffer.buffer[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5438_ (.CLK(net1063),
    .D(_0636_),
    .Q(\device.rxBuffer.buffer[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5439_ (.CLK(net1064),
    .D(_0637_),
    .Q(\device.rxBuffer.buffer[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5440_ (.CLK(net1065),
    .D(_0638_),
    .Q(\device.rxBuffer.buffer[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5441_ (.CLK(net1066),
    .D(_0639_),
    .Q(\device.txBuffer.buffer[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5442_ (.CLK(net1067),
    .D(_0640_),
    .Q(\device.txBuffer.buffer[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5443_ (.CLK(net1068),
    .D(_0641_),
    .Q(\device.txBuffer.buffer[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5444_ (.CLK(net1069),
    .D(_0642_),
    .Q(\device.txBuffer.buffer[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5445_ (.CLK(net1070),
    .D(_0643_),
    .Q(\device.txBuffer.buffer[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5446_ (.CLK(net1071),
    .D(_0644_),
    .Q(\device.txBuffer.buffer[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5447_ (.CLK(net1072),
    .D(_0645_),
    .Q(\device.txBuffer.buffer[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5448_ (.CLK(net1073),
    .D(_0646_),
    .Q(\device.txBuffer.buffer[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5449_ (.CLK(net1074),
    .D(_0647_),
    .Q(\device.rxBuffer.buffer[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5450_ (.CLK(net1075),
    .D(_0648_),
    .Q(\device.rxBuffer.buffer[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5451_ (.CLK(net1076),
    .D(_0649_),
    .Q(\device.rxBuffer.buffer[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5452_ (.CLK(net1077),
    .D(_0650_),
    .Q(\device.rxBuffer.buffer[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5453_ (.CLK(net1078),
    .D(_0651_),
    .Q(\device.rxBuffer.buffer[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5454_ (.CLK(net1079),
    .D(_0652_),
    .Q(\device.rxBuffer.buffer[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5455_ (.CLK(net1080),
    .D(_0653_),
    .Q(\device.rxBuffer.buffer[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5456_ (.CLK(net1081),
    .D(_0654_),
    .Q(\device.rxBuffer.buffer[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5457_ (.CLK(net1082),
    .D(_0655_),
    .Q(\device.txBuffer.buffer[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5458_ (.CLK(net1083),
    .D(_0656_),
    .Q(\device.txBuffer.buffer[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5459_ (.CLK(net1084),
    .D(_0657_),
    .Q(\device.txBuffer.buffer[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5460_ (.CLK(net1085),
    .D(_0658_),
    .Q(\device.txBuffer.buffer[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5461_ (.CLK(net1086),
    .D(_0659_),
    .Q(\device.txBuffer.buffer[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5462_ (.CLK(net1087),
    .D(_0660_),
    .Q(\device.txBuffer.buffer[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5463_ (.CLK(net1088),
    .D(_0661_),
    .Q(\device.txBuffer.buffer[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5464_ (.CLK(net1089),
    .D(_0662_),
    .Q(\device.txBuffer.buffer[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5465_ (.CLK(net1090),
    .D(_0663_),
    .Q(\device.txBuffer.buffer[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5466_ (.CLK(net1091),
    .D(_0664_),
    .Q(\device.txBuffer.buffer[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5467_ (.CLK(net1092),
    .D(_0665_),
    .Q(\device.txBuffer.buffer[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5468_ (.CLK(net1093),
    .D(_0666_),
    .Q(\device.txBuffer.buffer[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5469_ (.CLK(net1094),
    .D(_0667_),
    .Q(\device.txBuffer.buffer[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5470_ (.CLK(net1095),
    .D(_0668_),
    .Q(\device.txBuffer.buffer[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5471_ (.CLK(net1096),
    .D(_0669_),
    .Q(\device.txBuffer.buffer[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5472_ (.CLK(net1097),
    .D(_0670_),
    .Q(\device.txBuffer.buffer[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5473_ (.CLK(net1098),
    .D(_0671_),
    .Q(\device.txBuffer.buffer[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5474_ (.CLK(net1099),
    .D(_0672_),
    .Q(\device.txBuffer.buffer[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5475_ (.CLK(net1100),
    .D(_0673_),
    .Q(\device.txBuffer.buffer[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5476_ (.CLK(net1101),
    .D(_0674_),
    .Q(\device.txBuffer.buffer[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5477_ (.CLK(net1102),
    .D(_0675_),
    .Q(\device.txBuffer.buffer[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5478_ (.CLK(net1103),
    .D(_0676_),
    .Q(\device.txBuffer.buffer[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5479_ (.CLK(net1104),
    .D(_0677_),
    .Q(\device.txBuffer.buffer[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5480_ (.CLK(net1105),
    .D(_0678_),
    .Q(\device.txBuffer.buffer[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5481_ (.CLK(net1106),
    .D(_0679_),
    .Q(\device.txBuffer.buffer[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5482_ (.CLK(net1107),
    .D(_0680_),
    .Q(\device.txBuffer.buffer[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5483_ (.CLK(net1108),
    .D(_0681_),
    .Q(\device.txBuffer.buffer[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5484_ (.CLK(net1109),
    .D(_0682_),
    .Q(\device.txBuffer.buffer[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5485_ (.CLK(net1110),
    .D(_0683_),
    .Q(\device.txBuffer.buffer[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5486_ (.CLK(net1111),
    .D(_0684_),
    .Q(\device.txBuffer.buffer[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5487_ (.CLK(net1112),
    .D(_0685_),
    .Q(\device.txBuffer.buffer[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5488_ (.CLK(net1113),
    .D(_0686_),
    .Q(\device.txBuffer.buffer[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5489_ (.CLK(net1114),
    .D(_0687_),
    .Q(\device.txBuffer.buffer[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5490_ (.CLK(net1115),
    .D(_0688_),
    .Q(\device.txBuffer.buffer[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5491_ (.CLK(net1116),
    .D(_0689_),
    .Q(\device.txBuffer.buffer[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5492_ (.CLK(net1117),
    .D(_0690_),
    .Q(\device.txBuffer.buffer[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5493_ (.CLK(net1118),
    .D(_0691_),
    .Q(\device.txBuffer.buffer[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5494_ (.CLK(net1119),
    .D(_0692_),
    .Q(\device.txBuffer.buffer[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5495_ (.CLK(net1120),
    .D(_0693_),
    .Q(\device.txBuffer.buffer[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5496_ (.CLK(net1121),
    .D(_0694_),
    .Q(\device.txBuffer.buffer[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5497_ (.CLK(net1122),
    .D(_0695_),
    .Q(\device.txBuffer.buffer[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5498_ (.CLK(net1123),
    .D(_0696_),
    .Q(\device.txBuffer.buffer[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5499_ (.CLK(net1124),
    .D(_0697_),
    .Q(\device.txBuffer.buffer[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5500_ (.CLK(net1125),
    .D(_0698_),
    .Q(\device.txBuffer.buffer[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5501_ (.CLK(net1126),
    .D(_0699_),
    .Q(\device.txBuffer.buffer[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5502_ (.CLK(net1127),
    .D(_0700_),
    .Q(\device.txBuffer.buffer[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5503_ (.CLK(net1128),
    .D(_0701_),
    .Q(\device.txBuffer.buffer[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5504_ (.CLK(net1129),
    .D(_0702_),
    .Q(\device.txBuffer.buffer[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5505_ (.CLK(net1130),
    .D(_0703_),
    .Q(\device.txBuffer.buffer[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5506_ (.CLK(net1131),
    .D(_0704_),
    .Q(\device.txBuffer.buffer[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5507_ (.CLK(net1132),
    .D(_0705_),
    .Q(\device.txBuffer.buffer[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5508_ (.CLK(net1133),
    .D(_0706_),
    .Q(\device.txBuffer.buffer[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5509_ (.CLK(net1134),
    .D(_0707_),
    .Q(\device.txBuffer.buffer[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5510_ (.CLK(net1135),
    .D(_0708_),
    .Q(\device.txBuffer.buffer[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5511_ (.CLK(net1136),
    .D(_0709_),
    .Q(\device.txBuffer.buffer[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5512_ (.CLK(net1137),
    .D(_0710_),
    .Q(\device.txBuffer.buffer[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5513_ (.CLK(net1138),
    .D(_0711_),
    .Q(\device.txBuffer.buffer[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5514_ (.CLK(net1139),
    .D(_0712_),
    .Q(\device.txBuffer.buffer[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5515_ (.CLK(net1140),
    .D(_0713_),
    .Q(\device.txBuffer.buffer[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5516_ (.CLK(net1141),
    .D(_0714_),
    .Q(\device.txBuffer.buffer[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5517_ (.CLK(net1142),
    .D(_0715_),
    .Q(\device.txBuffer.buffer[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5518_ (.CLK(net1143),
    .D(_0716_),
    .Q(\device.txBuffer.buffer[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5519_ (.CLK(net1144),
    .D(_0717_),
    .Q(\device.txBuffer.buffer[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5520_ (.CLK(net1145),
    .D(_0718_),
    .Q(\device.txBuffer.buffer[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5521_ (.CLK(net1146),
    .D(_0719_),
    .Q(\device.txBuffer.buffer[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5522_ (.CLK(net1147),
    .D(_0720_),
    .Q(\device.txBuffer.buffer[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5523_ (.CLK(net1148),
    .D(_0721_),
    .Q(\device.txBuffer.buffer[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5524_ (.CLK(net1149),
    .D(_0722_),
    .Q(\device.txBuffer.buffer[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5525_ (.CLK(net1150),
    .D(_0723_),
    .Q(\device.txBuffer.buffer[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5526_ (.CLK(net1151),
    .D(_0724_),
    .Q(\device.txBuffer.buffer[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5527_ (.CLK(net1152),
    .D(_0725_),
    .Q(\device.txBuffer.buffer[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5528_ (.CLK(net1153),
    .D(_0726_),
    .Q(\device.txBuffer.buffer[31][7] ));
 sky130_fd_sc_hd__dfxtp_4 _5529_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_0727_),
    .Q(\device.uartTx.state[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5530_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_0728_),
    .Q(\device.uartTx.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5531_ (.CLK(net1154),
    .D(_0729_),
    .Q(\device.rxBuffer.buffer[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5532_ (.CLK(net1155),
    .D(_0730_),
    .Q(\device.rxBuffer.buffer[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5533_ (.CLK(net1156),
    .D(_0731_),
    .Q(\device.rxBuffer.buffer[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5534_ (.CLK(net1157),
    .D(_0732_),
    .Q(\device.rxBuffer.buffer[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5535_ (.CLK(net1158),
    .D(_0733_),
    .Q(\device.rxBuffer.buffer[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5536_ (.CLK(net1159),
    .D(_0734_),
    .Q(\device.rxBuffer.buffer[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5537_ (.CLK(net1160),
    .D(_0735_),
    .Q(\device.rxBuffer.buffer[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5538_ (.CLK(net1161),
    .D(_0736_),
    .Q(\device.rxBuffer.buffer[18][7] ));
 sky130_fd_sc_hd__dfxtp_4 _5539_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_0737_),
    .Q(\device.uartTx.delayCounter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5540_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_0738_),
    .Q(\device.uartTx.delayCounter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _5541_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net1949),
    .Q(\device.uartTx.delayCounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5542_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net1985),
    .Q(\device.uartTx.delayCounter[3] ));
 sky130_fd_sc_hd__dfxtp_4 _5543_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_0741_),
    .Q(\device.uartTx.delayCounter[4] ));
 sky130_fd_sc_hd__dfxtp_2 _5544_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_0742_),
    .Q(\device.uartTx.delayCounter[5] ));
 sky130_fd_sc_hd__dfxtp_2 _5545_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_0743_),
    .Q(\device.uartTx.delayCounter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5546_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_0744_),
    .Q(\device.uartTx.delayCounter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5547_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_0745_),
    .Q(\device.uartTx.delayCounter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _5548_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_0746_),
    .Q(\device.uartTx.delayCounter[9] ));
 sky130_fd_sc_hd__dfxtp_2 _5549_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_0747_),
    .Q(\device.uartTx.delayCounter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _5550_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_0748_),
    .Q(\device.uartTx.delayCounter[11] ));
 sky130_fd_sc_hd__dfxtp_2 _5551_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_0749_),
    .Q(\device.uartTx.delayCounter[12] ));
 sky130_fd_sc_hd__dfxtp_2 _5552_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_0750_),
    .Q(\device.uartTx.delayCounter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _5553_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_0751_),
    .Q(\device.uartTx.delayCounter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _5554_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_0752_),
    .Q(\device.uartTx.delayCounter[15] ));
 sky130_fd_sc_hd__dfxtp_2 _5555_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_0753_),
    .Q(\device.uartTx.bitCounter[0] ));
 sky130_fd_sc_hd__dfxtp_2 _5556_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_0754_),
    .Q(\device.uartTx.bitCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5557_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_0755_),
    .Q(\device.uartTx.bitCounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5558_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_0756_),
    .Q(\device.uartTx.savedData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5559_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_0757_),
    .Q(\device.uartTx.savedData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5560_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_0758_),
    .Q(\device.uartTx.savedData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5561_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_0759_),
    .Q(\device.uartTx.savedData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5562_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_0760_),
    .Q(\device.uartTx.savedData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5563_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_0761_),
    .Q(\device.uartTx.savedData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5564_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(net1854),
    .Q(\device.uartTx.savedData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5565_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(net1877),
    .Q(\device.uartTx.savedData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5566_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_0764_),
    .Q(\device.txSendBusy ));
 sky130_fd_sc_hd__dfxtp_1 _5567_ (.CLK(net1162),
    .D(_0765_),
    .Q(\device.rxBuffer.buffer[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5568_ (.CLK(net1163),
    .D(_0766_),
    .Q(\device.rxBuffer.buffer[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5569_ (.CLK(net1164),
    .D(_0767_),
    .Q(\device.rxBuffer.buffer[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5570_ (.CLK(net1165),
    .D(_0768_),
    .Q(\device.rxBuffer.buffer[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5571_ (.CLK(net1166),
    .D(_0769_),
    .Q(\device.rxBuffer.buffer[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5572_ (.CLK(net1167),
    .D(_0770_),
    .Q(\device.rxBuffer.buffer[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5573_ (.CLK(net1168),
    .D(_0771_),
    .Q(\device.rxBuffer.buffer[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5574_ (.CLK(net1169),
    .D(_0772_),
    .Q(\device.rxBuffer.buffer[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5575_ (.CLK(net1170),
    .D(_0773_),
    .Q(\device.txBuffer.buffer[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5576_ (.CLK(net1171),
    .D(_0774_),
    .Q(\device.txBuffer.buffer[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5577_ (.CLK(net1172),
    .D(_0775_),
    .Q(\device.txBuffer.buffer[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5578_ (.CLK(net1173),
    .D(_0776_),
    .Q(\device.txBuffer.buffer[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5579_ (.CLK(net1174),
    .D(_0777_),
    .Q(\device.txBuffer.buffer[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5580_ (.CLK(net1175),
    .D(_0778_),
    .Q(\device.txBuffer.buffer[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5581_ (.CLK(net1176),
    .D(_0779_),
    .Q(\device.txBuffer.buffer[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5582_ (.CLK(net1177),
    .D(_0780_),
    .Q(\device.txBuffer.buffer[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5583_ (.CLK(net1178),
    .D(_0781_),
    .Q(\device.rxBuffer.buffer[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5584_ (.CLK(net1179),
    .D(_0782_),
    .Q(\device.rxBuffer.buffer[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5585_ (.CLK(net1180),
    .D(_0783_),
    .Q(\device.rxBuffer.buffer[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5586_ (.CLK(net1181),
    .D(_0784_),
    .Q(\device.rxBuffer.buffer[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5587_ (.CLK(net1182),
    .D(_0785_),
    .Q(\device.rxBuffer.buffer[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5588_ (.CLK(net1183),
    .D(_0786_),
    .Q(\device.rxBuffer.buffer[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5589_ (.CLK(net1184),
    .D(_0787_),
    .Q(\device.rxBuffer.buffer[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5590_ (.CLK(net1185),
    .D(_0788_),
    .Q(\device.rxBuffer.buffer[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5591_ (.CLK(net1186),
    .D(_0789_),
    .Q(\device.txBuffer.buffer[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5592_ (.CLK(net1187),
    .D(_0790_),
    .Q(\device.txBuffer.buffer[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5593_ (.CLK(net1188),
    .D(_0791_),
    .Q(\device.txBuffer.buffer[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5594_ (.CLK(net1189),
    .D(_0792_),
    .Q(\device.txBuffer.buffer[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5595_ (.CLK(net1190),
    .D(_0793_),
    .Q(\device.txBuffer.buffer[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5596_ (.CLK(net1191),
    .D(_0794_),
    .Q(\device.txBuffer.buffer[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5597_ (.CLK(net1192),
    .D(_0795_),
    .Q(\device.txBuffer.buffer[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5598_ (.CLK(net1193),
    .D(_0796_),
    .Q(\device.txBuffer.buffer[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5599_ (.CLK(net1194),
    .D(_0797_),
    .Q(\device.rxBuffer.buffer[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5600_ (.CLK(net1195),
    .D(_0798_),
    .Q(\device.rxBuffer.buffer[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5601_ (.CLK(net1196),
    .D(_0799_),
    .Q(\device.rxBuffer.buffer[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5602_ (.CLK(net1197),
    .D(_0800_),
    .Q(\device.rxBuffer.buffer[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5603_ (.CLK(net1198),
    .D(_0801_),
    .Q(\device.rxBuffer.buffer[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5604_ (.CLK(net1199),
    .D(_0802_),
    .Q(\device.rxBuffer.buffer[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5605_ (.CLK(net1200),
    .D(_0803_),
    .Q(\device.rxBuffer.buffer[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5606_ (.CLK(net1201),
    .D(_0804_),
    .Q(\device.rxBuffer.buffer[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5607_ (.CLK(net1202),
    .D(_0805_),
    .Q(\device.txBuffer.buffer[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5608_ (.CLK(net1203),
    .D(_0806_),
    .Q(\device.txBuffer.buffer[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5609_ (.CLK(net1204),
    .D(_0807_),
    .Q(\device.txBuffer.buffer[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5610_ (.CLK(net1205),
    .D(_0808_),
    .Q(\device.txBuffer.buffer[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5611_ (.CLK(net1206),
    .D(_0809_),
    .Q(\device.txBuffer.buffer[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5612_ (.CLK(net1207),
    .D(_0810_),
    .Q(\device.txBuffer.buffer[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5613_ (.CLK(net1208),
    .D(_0811_),
    .Q(\device.txBuffer.buffer[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5614_ (.CLK(net1209),
    .D(_0812_),
    .Q(\device.txBuffer.buffer[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5615_ (.CLK(net1210),
    .D(_0813_),
    .Q(\device.txBuffer.buffer[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5616_ (.CLK(net1211),
    .D(_0814_),
    .Q(\device.txBuffer.buffer[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5617_ (.CLK(net1212),
    .D(_0815_),
    .Q(\device.txBuffer.buffer[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5618_ (.CLK(net1213),
    .D(_0816_),
    .Q(\device.txBuffer.buffer[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5619_ (.CLK(net1214),
    .D(_0817_),
    .Q(\device.txBuffer.buffer[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5620_ (.CLK(net1215),
    .D(_0818_),
    .Q(\device.txBuffer.buffer[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5621_ (.CLK(net1216),
    .D(_0819_),
    .Q(\device.txBuffer.buffer[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5622_ (.CLK(net1217),
    .D(_0820_),
    .Q(\device.txBuffer.buffer[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5623_ (.CLK(net1218),
    .D(_0821_),
    .Q(\device.txBuffer.buffer[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5624_ (.CLK(net1219),
    .D(_0822_),
    .Q(\device.txBuffer.buffer[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5625_ (.CLK(net1220),
    .D(_0823_),
    .Q(\device.txBuffer.buffer[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5626_ (.CLK(net1221),
    .D(_0824_),
    .Q(\device.txBuffer.buffer[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5627_ (.CLK(net1222),
    .D(_0825_),
    .Q(\device.txBuffer.buffer[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5628_ (.CLK(net1223),
    .D(_0826_),
    .Q(\device.txBuffer.buffer[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5629_ (.CLK(net1224),
    .D(_0827_),
    .Q(\device.txBuffer.buffer[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5630_ (.CLK(net1225),
    .D(_0828_),
    .Q(\device.txBuffer.buffer[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5631_ (.CLK(net1226),
    .D(_0829_),
    .Q(\device.txBuffer.buffer[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5632_ (.CLK(net1227),
    .D(_0830_),
    .Q(\device.txBuffer.buffer[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5633_ (.CLK(net1228),
    .D(_0831_),
    .Q(\device.txBuffer.buffer[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5634_ (.CLK(net1229),
    .D(_0832_),
    .Q(\device.txBuffer.buffer[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5635_ (.CLK(net1230),
    .D(_0833_),
    .Q(\device.txBuffer.buffer[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5636_ (.CLK(net1231),
    .D(_0834_),
    .Q(\device.txBuffer.buffer[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5637_ (.CLK(net1232),
    .D(_0835_),
    .Q(\device.txBuffer.buffer[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5638_ (.CLK(net1233),
    .D(_0836_),
    .Q(\device.txBuffer.buffer[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5639_ (.CLK(net1234),
    .D(_0837_),
    .Q(\device.txBuffer.buffer[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5640_ (.CLK(net1235),
    .D(_0838_),
    .Q(\device.txBuffer.buffer[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5641_ (.CLK(net1236),
    .D(_0839_),
    .Q(\device.txBuffer.buffer[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5642_ (.CLK(net1237),
    .D(_0840_),
    .Q(\device.txBuffer.buffer[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5643_ (.CLK(net1238),
    .D(_0841_),
    .Q(\device.txBuffer.buffer[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5644_ (.CLK(net1239),
    .D(_0842_),
    .Q(\device.txBuffer.buffer[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5645_ (.CLK(net1240),
    .D(_0843_),
    .Q(\device.txBuffer.buffer[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5646_ (.CLK(net1241),
    .D(_0844_),
    .Q(\device.txBuffer.buffer[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5647_ (.CLK(net1242),
    .D(_0845_),
    .Q(\device.txBuffer.buffer[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5648_ (.CLK(net1243),
    .D(_0846_),
    .Q(\device.txBuffer.buffer[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5649_ (.CLK(net1244),
    .D(_0847_),
    .Q(\device.txBuffer.buffer[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5650_ (.CLK(net1245),
    .D(_0848_),
    .Q(\device.txBuffer.buffer[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5651_ (.CLK(net1246),
    .D(_0849_),
    .Q(\device.txBuffer.buffer[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5652_ (.CLK(net1247),
    .D(_0850_),
    .Q(\device.txBuffer.buffer[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5653_ (.CLK(net1248),
    .D(_0851_),
    .Q(\device.txBuffer.buffer[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5654_ (.CLK(net1249),
    .D(_0852_),
    .Q(\device.txBuffer.buffer[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5655_ (.CLK(net1250),
    .D(_0853_),
    .Q(\device.txBuffer.buffer[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5656_ (.CLK(net1251),
    .D(_0854_),
    .Q(\device.txBuffer.buffer[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5657_ (.CLK(net1252),
    .D(_0855_),
    .Q(\device.txBuffer.buffer[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5658_ (.CLK(net1253),
    .D(_0856_),
    .Q(\device.txBuffer.buffer[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5659_ (.CLK(net1254),
    .D(_0857_),
    .Q(\device.txBuffer.buffer[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5660_ (.CLK(net1255),
    .D(_0858_),
    .Q(\device.txBuffer.buffer[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5661_ (.CLK(net1256),
    .D(_0859_),
    .Q(\device.txBuffer.buffer[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5662_ (.CLK(net1257),
    .D(_0860_),
    .Q(\device.txBuffer.buffer[15][7] ));
 sky130_fd_sc_hd__dfxtp_4 _5663_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_0861_),
    .Q(\device.uartRx.state[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5664_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_0862_),
    .Q(\device.uartRx.state[1] ));
 sky130_fd_sc_hd__dfxtp_4 _5665_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0863_),
    .Q(\device.uartRx.delayCounter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5666_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0864_),
    .Q(\device.uartRx.delayCounter[1] ));
 sky130_fd_sc_hd__dfxtp_4 _5667_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0865_),
    .Q(\device.uartRx.delayCounter[2] ));
 sky130_fd_sc_hd__dfxtp_2 _5668_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0866_),
    .Q(\device.uartRx.delayCounter[3] ));
 sky130_fd_sc_hd__dfxtp_4 _5669_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0867_),
    .Q(\device.uartRx.delayCounter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5670_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0868_),
    .Q(\device.uartRx.delayCounter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5671_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0869_),
    .Q(\device.uartRx.delayCounter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5672_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0870_),
    .Q(\device.uartRx.delayCounter[7] ));
 sky130_fd_sc_hd__dfxtp_2 _5673_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0871_),
    .Q(\device.uartRx.delayCounter[8] ));
 sky130_fd_sc_hd__dfxtp_2 _5674_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0872_),
    .Q(\device.uartRx.delayCounter[9] ));
 sky130_fd_sc_hd__dfxtp_2 _5675_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_0873_),
    .Q(\device.uartRx.delayCounter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _5676_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(net1707),
    .Q(\device.uartRx.delayCounter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _5677_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net1714),
    .Q(\device.uartRx.delayCounter[12] ));
 sky130_fd_sc_hd__dfxtp_4 _5678_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_0876_),
    .Q(\device.uartRx.delayCounter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _5679_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_0877_),
    .Q(\device.uartRx.delayCounter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _5680_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(net1765),
    .Q(\device.uartRx.delayCounter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _5681_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_0879_),
    .Q(\device.uartRx.bitCounter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5682_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0880_),
    .Q(\device.uartRx.bitCounter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5683_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_0881_),
    .Q(\device.uartRx.bitCounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5684_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_0882_),
    .Q(\device.uartRx.savedData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5685_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_0883_),
    .Q(\device.uartRx.savedData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5686_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_0884_),
    .Q(\device.uartRx.savedData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5687_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0885_),
    .Q(\device.uartRx.savedData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5688_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0886_),
    .Q(\device.uartRx.savedData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5689_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0887_),
    .Q(\device.uartRx.savedData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5690_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0888_),
    .Q(\device.uartRx.savedData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _5691_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_0889_),
    .Q(\device.uartRx.savedData[7] ));
 sky130_fd_sc_hd__dfxtp_4 _5692_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net3653),
    .Q(\device.txBuffer.dataIn_buffered[0] ));
 sky130_fd_sc_hd__dfxtp_4 _5693_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net4075),
    .Q(\device.txBuffer.dataIn_buffered[1] ));
 sky130_fd_sc_hd__dfxtp_4 _5694_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net3640),
    .Q(\device.txBuffer.dataIn_buffered[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5695_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net3604),
    .Q(\device.txBuffer.dataIn_buffered[3] ));
 sky130_fd_sc_hd__dfxtp_4 _5696_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net3627),
    .Q(\device.txBuffer.dataIn_buffered[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5697_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net3591),
    .Q(\device.txBuffer.dataIn_buffered[5] ));
 sky130_fd_sc_hd__dfxtp_4 _5698_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net3270),
    .Q(\device.txBuffer.dataIn_buffered[6] ));
 sky130_fd_sc_hd__dfxtp_2 _5699_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net3259),
    .Q(\device.txBuffer.dataIn_buffered[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5700_ (.CLK(net1258),
    .D(_0898_),
    .Q(\device.txBuffer.buffer[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5701_ (.CLK(net1259),
    .D(_0899_),
    .Q(\device.txBuffer.buffer[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5702_ (.CLK(net1260),
    .D(_0900_),
    .Q(\device.txBuffer.buffer[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5703_ (.CLK(net1261),
    .D(_0901_),
    .Q(\device.txBuffer.buffer[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5704_ (.CLK(net1262),
    .D(_0902_),
    .Q(\device.txBuffer.buffer[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5705_ (.CLK(net1263),
    .D(_0903_),
    .Q(\device.txBuffer.buffer[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5706_ (.CLK(net1264),
    .D(_0904_),
    .Q(\device.txBuffer.buffer[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5707_ (.CLK(net1265),
    .D(_0905_),
    .Q(\device.txBuffer.buffer[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5708_ (.CLK(net1266),
    .D(_0906_),
    .Q(\device.txBuffer.buffer[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5709_ (.CLK(net1267),
    .D(_0907_),
    .Q(\device.txBuffer.buffer[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5710_ (.CLK(net1268),
    .D(_0908_),
    .Q(\device.txBuffer.buffer[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5711_ (.CLK(net1269),
    .D(_0909_),
    .Q(\device.txBuffer.buffer[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5712_ (.CLK(net1270),
    .D(_0910_),
    .Q(\device.txBuffer.buffer[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5713_ (.CLK(net1271),
    .D(_0911_),
    .Q(\device.txBuffer.buffer[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5714_ (.CLK(net1272),
    .D(_0912_),
    .Q(\device.txBuffer.buffer[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5715_ (.CLK(net1273),
    .D(_0913_),
    .Q(\device.txBuffer.buffer[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5716_ (.CLK(net1274),
    .D(_0914_),
    .Q(\device.txBuffer.buffer[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5717_ (.CLK(net1275),
    .D(_0915_),
    .Q(\device.txBuffer.buffer[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5718_ (.CLK(net1276),
    .D(_0916_),
    .Q(\device.txBuffer.buffer[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5719_ (.CLK(net1277),
    .D(_0917_),
    .Q(\device.txBuffer.buffer[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5720_ (.CLK(net1278),
    .D(_0918_),
    .Q(\device.txBuffer.buffer[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5721_ (.CLK(net1279),
    .D(_0919_),
    .Q(\device.txBuffer.buffer[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5722_ (.CLK(net1280),
    .D(_0920_),
    .Q(\device.txBuffer.buffer[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5723_ (.CLK(net1281),
    .D(_0921_),
    .Q(\device.txBuffer.buffer[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5724_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net3860),
    .Q(\device.rxBufferFullBuffered ));
 sky130_fd_sc_hd__dfxtp_1 _5725_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0923_),
    .Q(\device.rxDataLostBuffered ));
 sky130_fd_sc_hd__dfxtp_2 _5726_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(net3470),
    .Q(\device.txDataAvailableBuffered ));
 sky130_fd_sc_hd__dfxtp_1 _5727_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net3138),
    .Q(\device.txBufferFullBuffered ));
 sky130_fd_sc_hd__dfxtp_1 _5728_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0926_),
    .Q(\device.txDataLostBuffered ));
 sky130_fd_sc_hd__dfxtp_1 _5729_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0927_),
    .Q(\device.statusRegister.baseReadData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _5730_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0928_),
    .Q(\device.statusRegister.baseReadData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5731_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0929_),
    .Q(\device.statusRegister.baseReadData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5732_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0930_),
    .Q(\device.statusRegister.baseReadData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5733_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0931_),
    .Q(\device.statusRegister.baseReadData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _5734_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0932_),
    .Q(\device.statusRegister.baseReadData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5735_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(net3108),
    .Q(\device.configuration[20] ));
 sky130_fd_sc_hd__dfxtp_1 _5736_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(net3236),
    .Q(\device.configuration[19] ));
 sky130_fd_sc_hd__dfxtp_1 _5737_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(net3214),
    .Q(\device.configuration[18] ));
 sky130_fd_sc_hd__dfxtp_4 _5738_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(net3131),
    .Q(\device.configuration[17] ));
 sky130_fd_sc_hd__dfxtp_2 _5739_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net3159),
    .Q(\device.configuration[16] ));
 sky130_fd_sc_hd__dfxtp_4 _5740_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(net3225),
    .Q(\device.configuration[15] ));
 sky130_fd_sc_hd__dfxtp_4 _5741_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(net3203),
    .Q(\device.configuration[14] ));
 sky130_fd_sc_hd__dfxtp_4 _5742_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(net3181),
    .Q(\device.configuration[13] ));
 sky130_fd_sc_hd__dfxtp_4 _5743_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net3276),
    .Q(\device.configuration[12] ));
 sky130_fd_sc_hd__dfxtp_4 _5744_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net3192),
    .Q(\device.configuration[11] ));
 sky130_fd_sc_hd__dfxtp_4 _5745_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net3170),
    .Q(\device.configuration[10] ));
 sky130_fd_sc_hd__dfxtp_4 _5746_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net2108),
    .Q(\device.configuration[9] ));
 sky130_fd_sc_hd__dfxtp_4 _5747_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0945_),
    .Q(\device.configuration[8] ));
 sky130_fd_sc_hd__dfxtp_2 _5748_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net1973),
    .Q(\device.configuration[7] ));
 sky130_fd_sc_hd__dfxtp_4 _5749_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net1751),
    .Q(\device.configuration[6] ));
 sky130_fd_sc_hd__dfxtp_4 _5750_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net3666),
    .Q(\device.configuration[5] ));
 sky130_fd_sc_hd__dfxtp_4 _5751_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net3689),
    .Q(\device.configuration[4] ));
 sky130_fd_sc_hd__dfxtp_4 _5752_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net4181),
    .Q(\device.configuration[3] ));
 sky130_fd_sc_hd__dfxtp_4 _5753_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net3850),
    .Q(\device.configuration[2] ));
 sky130_fd_sc_hd__dfxtp_4 _5754_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net2932),
    .Q(\device.configuration[1] ));
 sky130_fd_sc_hd__dfxtp_2 _5755_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net3837),
    .Q(\device.configuration[0] ));
 sky130_fd_sc_hd__clkbuf_4 _5837_ (.A(net36),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 _5838_ (.A(net47),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_4 _5839_ (.A(net58),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_4 _5840_ (.A(net69),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_4 _5841_ (.A(net80),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_4 _5842_ (.A(net91),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_4 _5843_ (.A(net102),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_4 _5844_ (.A(net113),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_4 _5845_ (.A(net124),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_4 _5846_ (.A(net133),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_4 _5847_ (.A(net37),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 _5848_ (.A(net38),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_4 _5849_ (.A(net39),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 _5850_ (.A(net40),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 _5851_ (.A(net41),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 _5852_ (.A(net42),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_4 _5853_ (.A(net43),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_4 _5854_ (.A(net44),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 _5855_ (.A(net45),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_4 _5856_ (.A(net46),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 _5857_ (.A(net48),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 _5858_ (.A(net49),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 _5859_ (.A(net50),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_4 _5860_ (.A(net51),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_4 _5861_ (.A(net52),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 _5862_ (.A(net53),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 _5863_ (.A(net54),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 _5864_ (.A(net55),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_4 _5865_ (.A(net56),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 _5866_ (.A(net57),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 _5867_ (.A(net59),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_4 _5868_ (.A(net60),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_4 _5869_ (.A(net61),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_4 _5870_ (.A(net62),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_4 _5871_ (.A(net63),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 _5872_ (.A(net64),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_4 _5873_ (.A(net65),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 _5874_ (.A(net66),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_4 _5875_ (.A(net67),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_4 _5876_ (.A(net68),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_4 _5877_ (.A(net70),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_4 _5878_ (.A(net71),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_4 _5879_ (.A(net72),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_4 _5880_ (.A(net73),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_4 _5881_ (.A(net74),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_4 _5882_ (.A(net75),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 _5883_ (.A(net76),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_4 _5884_ (.A(net77),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_4 _5885_ (.A(net78),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_4 _5886_ (.A(net79),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_4 _5887_ (.A(net81),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_4 _5888_ (.A(net82),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_4 _5889_ (.A(net83),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_4 _5890_ (.A(net84),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_4 _5891_ (.A(net85),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_4 _5892_ (.A(net86),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_4 _5893_ (.A(net87),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_4 _5894_ (.A(net88),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_4 _5895_ (.A(net89),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_4 _5896_ (.A(net90),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_4 _5897_ (.A(net92),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_4 _5898_ (.A(net93),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_4 _5899_ (.A(net94),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_4 _5900_ (.A(net95),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_4 _5901_ (.A(net96),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_4 _5902_ (.A(net97),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_4 _5903_ (.A(net98),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_4 _5904_ (.A(net99),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_4 _5905_ (.A(net100),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_4 _5906_ (.A(net101),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_4 _5907_ (.A(net103),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_4 _5908_ (.A(net104),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_4 _5909_ (.A(net105),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_4 _5910_ (.A(net106),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_4 _5911_ (.A(net107),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 _5912_ (.A(net108),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_4 _5913_ (.A(net109),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_4 _5914_ (.A(net110),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_4 _5915_ (.A(net111),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_4 _5916_ (.A(net112),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_4 _5917_ (.A(net114),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_4 _5918_ (.A(net115),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 _5919_ (.A(net116),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_4 _5920_ (.A(net117),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_4 _5921_ (.A(net118),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_4 _5922_ (.A(net119),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_4 _5923_ (.A(net120),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_4 _5924_ (.A(net121),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_4 _5925_ (.A(net122),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_4 _5926_ (.A(net123),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_4 _5927_ (.A(net125),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 _5928_ (.A(net126),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_4 _5929_ (.A(net127),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_4 _5930_ (.A(net128),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_4 _5931_ (.A(net129),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_4 _5932_ (.A(net130),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_4 _5933_ (.A(net131),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_4 _5934_ (.A(net132),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_4_0_0_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.A(clknet_4_4_0_wb_clk_i),
    .X(clknet_leaf_100_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.A(clknet_4_4_0_wb_clk_i),
    .X(clknet_leaf_101_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.A(clknet_4_6_0_wb_clk_i),
    .X(clknet_leaf_102_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.A(clknet_4_6_0_wb_clk_i),
    .X(clknet_leaf_103_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.A(clknet_4_6_0_wb_clk_i),
    .X(clknet_leaf_104_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.A(clknet_4_6_0_wb_clk_i),
    .X(clknet_leaf_105_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.A(clknet_4_3_0_wb_clk_i),
    .X(clknet_leaf_106_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.A(clknet_4_3_0_wb_clk_i),
    .X(clknet_leaf_108_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.A(clknet_4_3_0_wb_clk_i),
    .X(clknet_leaf_109_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_4_2_0_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.A(clknet_4_3_0_wb_clk_i),
    .X(clknet_leaf_110_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.A(clknet_4_1_0_wb_clk_i),
    .X(clknet_leaf_111_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.A(clknet_4_1_0_wb_clk_i),
    .X(clknet_leaf_112_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.A(clknet_4_1_0_wb_clk_i),
    .X(clknet_leaf_113_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.A(clknet_4_1_0_wb_clk_i),
    .X(clknet_leaf_114_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.A(clknet_4_1_0_wb_clk_i),
    .X(clknet_leaf_115_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.A(clknet_4_1_0_wb_clk_i),
    .X(clknet_leaf_116_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.A(clknet_4_1_0_wb_clk_i),
    .X(clknet_leaf_117_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.A(clknet_4_0_0_wb_clk_i),
    .X(clknet_leaf_118_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.A(clknet_4_0_0_wb_clk_i),
    .X(clknet_leaf_119_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_4_3_0_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.A(clknet_4_0_0_wb_clk_i),
    .X(clknet_leaf_120_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.A(clknet_4_0_0_wb_clk_i),
    .X(clknet_leaf_121_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.A(clknet_4_0_0_wb_clk_i),
    .X(clknet_leaf_122_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_4_9_0_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_4_9_0_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_4_9_0_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_4_9_0_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_4_8_0_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_4_8_0_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_4_8_0_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_4_8_0_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_4_0_0_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_4_8_0_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_4_8_0_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_4_8_0_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_4_8_0_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_4_10_0_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_4_10_0_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_4_10_0_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_4_10_0_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_4_10_0_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_4_10_0_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_4_2_0_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_4_10_0_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_4_10_0_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_4_10_0_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_4_11_0_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_4_11_0_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_4_11_0_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_4_11_0_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_4_14_0_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_4_14_0_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_4_14_0_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_4_2_0_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_4_11_0_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_4_11_0_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_4_9_0_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_4_9_0_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_4_12_0_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_4_12_0_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_4_12_0_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_4_12_0_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_4_12_0_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_4_2_0_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_4_14_0_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.A(clknet_4_14_0_wb_clk_i),
    .X(clknet_leaf_51_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.A(clknet_4_14_0_wb_clk_i),
    .X(clknet_leaf_52_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.A(clknet_4_14_0_wb_clk_i),
    .X(clknet_leaf_53_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.A(clknet_4_14_0_wb_clk_i),
    .X(clknet_leaf_54_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.A(clknet_4_15_0_wb_clk_i),
    .X(clknet_leaf_55_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.A(clknet_4_15_0_wb_clk_i),
    .X(clknet_leaf_56_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.A(clknet_4_15_0_wb_clk_i),
    .X(clknet_leaf_57_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.A(clknet_4_15_0_wb_clk_i),
    .X(clknet_leaf_58_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.A(clknet_4_15_0_wb_clk_i),
    .X(clknet_leaf_59_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_4_2_0_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.A(clknet_4_15_0_wb_clk_i),
    .X(clknet_leaf_60_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.A(clknet_4_15_0_wb_clk_i),
    .X(clknet_leaf_61_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.A(clknet_4_15_0_wb_clk_i),
    .X(clknet_leaf_63_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.A(clknet_4_13_0_wb_clk_i),
    .X(clknet_leaf_64_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.A(clknet_4_13_0_wb_clk_i),
    .X(clknet_leaf_65_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.A(clknet_4_13_0_wb_clk_i),
    .X(clknet_leaf_66_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.A(clknet_4_13_0_wb_clk_i),
    .X(clknet_leaf_67_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.A(clknet_4_13_0_wb_clk_i),
    .X(clknet_leaf_68_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.A(clknet_4_13_0_wb_clk_i),
    .X(clknet_leaf_69_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_4_2_0_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.A(clknet_4_13_0_wb_clk_i),
    .X(clknet_leaf_70_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.A(clknet_4_13_0_wb_clk_i),
    .X(clknet_leaf_71_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.A(clknet_4_12_0_wb_clk_i),
    .X(clknet_leaf_72_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.A(clknet_4_6_0_wb_clk_i),
    .X(clknet_leaf_73_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.A(clknet_4_6_0_wb_clk_i),
    .X(clknet_leaf_74_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.A(clknet_4_6_0_wb_clk_i),
    .X(clknet_leaf_75_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.A(clknet_4_6_0_wb_clk_i),
    .X(clknet_leaf_76_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.A(clknet_4_7_0_wb_clk_i),
    .X(clknet_leaf_77_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.A(clknet_4_7_0_wb_clk_i),
    .X(clknet_leaf_78_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.A(clknet_4_7_0_wb_clk_i),
    .X(clknet_leaf_79_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_4_2_0_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.A(clknet_4_7_0_wb_clk_i),
    .X(clknet_leaf_80_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.A(clknet_4_7_0_wb_clk_i),
    .X(clknet_leaf_81_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.A(clknet_4_7_0_wb_clk_i),
    .X(clknet_leaf_83_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.A(clknet_4_7_0_wb_clk_i),
    .X(clknet_leaf_84_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.A(clknet_4_7_0_wb_clk_i),
    .X(clknet_leaf_85_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.A(clknet_4_5_0_wb_clk_i),
    .X(clknet_leaf_86_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.A(clknet_4_5_0_wb_clk_i),
    .X(clknet_leaf_87_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.A(clknet_4_5_0_wb_clk_i),
    .X(clknet_leaf_88_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.A(clknet_4_5_0_wb_clk_i),
    .X(clknet_leaf_89_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_4_2_0_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.A(clknet_4_5_0_wb_clk_i),
    .X(clknet_leaf_90_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.A(clknet_4_5_0_wb_clk_i),
    .X(clknet_leaf_91_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.A(clknet_4_5_0_wb_clk_i),
    .X(clknet_leaf_92_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.A(clknet_4_5_0_wb_clk_i),
    .X(clknet_leaf_93_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.A(clknet_4_4_0_wb_clk_i),
    .X(clknet_leaf_94_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.A(clknet_4_4_0_wb_clk_i),
    .X(clknet_leaf_95_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.A(clknet_4_4_0_wb_clk_i),
    .X(clknet_leaf_96_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.A(clknet_4_4_0_wb_clk_i),
    .X(clknet_leaf_97_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.A(clknet_4_4_0_wb_clk_i),
    .X(clknet_leaf_98_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.A(clknet_4_4_0_wb_clk_i),
    .X(clknet_leaf_99_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_4_2_0_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__buf_4 fanout406 (.A(_2363_),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_4 fanout407 (.A(_2363_),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_4 fanout408 (.A(_2298_),
    .X(net408));
 sky130_fd_sc_hd__buf_4 fanout409 (.A(_2295_),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_2 fanout410 (.A(_2295_),
    .X(net410));
 sky130_fd_sc_hd__buf_6 fanout411 (.A(_2104_),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_4 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__buf_4 fanout413 (.A(_1724_),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_4 fanout414 (.A(net415),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_4 fanout415 (.A(net235),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_4 fanout416 (.A(net235),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_2 fanout417 (.A(net235),
    .X(net417));
 sky130_fd_sc_hd__buf_6 fanout418 (.A(_1723_),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_4 fanout419 (.A(net1787),
    .X(net419));
 sky130_fd_sc_hd__buf_4 fanout420 (.A(net1764),
    .X(net420));
 sky130_fd_sc_hd__buf_4 fanout421 (.A(net1763),
    .X(net421));
 sky130_fd_sc_hd__buf_8 fanout422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__buf_6 fanout423 (.A(net1602),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_16 fanout424 (.A(net1598),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_8 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_6 fanout426 (.A(_2057_),
    .X(net426));
 sky130_fd_sc_hd__buf_4 fanout427 (.A(net1984),
    .X(net427));
 sky130_fd_sc_hd__buf_6 fanout428 (.A(net1982),
    .X(net428));
 sky130_fd_sc_hd__buf_4 fanout429 (.A(net2022),
    .X(net429));
 sky130_fd_sc_hd__buf_8 fanout430 (.A(_2021_),
    .X(net430));
 sky130_fd_sc_hd__buf_4 fanout431 (.A(_1977_),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_2 fanout432 (.A(_1977_),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_4 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__buf_4 fanout434 (.A(_1977_),
    .X(net434));
 sky130_fd_sc_hd__buf_4 fanout435 (.A(_1497_),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_4 fanout436 (.A(_1497_),
    .X(net436));
 sky130_fd_sc_hd__buf_4 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_6 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__buf_6 fanout439 (.A(_1442_),
    .X(net439));
 sky130_fd_sc_hd__buf_4 fanout440 (.A(net442),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_2 fanout441 (.A(net1284),
    .X(net441));
 sky130_fd_sc_hd__buf_6 fanout442 (.A(_1419_),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_4 fanout443 (.A(_2423_),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_4 fanout444 (.A(_2413_),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_2 fanout445 (.A(_2413_),
    .X(net445));
 sky130_fd_sc_hd__buf_8 fanout446 (.A(_1975_),
    .X(net446));
 sky130_fd_sc_hd__buf_6 fanout447 (.A(_1975_),
    .X(net447));
 sky130_fd_sc_hd__buf_6 fanout448 (.A(_1975_),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_4 fanout449 (.A(_1975_),
    .X(net449));
 sky130_fd_sc_hd__buf_6 fanout450 (.A(_1739_),
    .X(net450));
 sky130_fd_sc_hd__buf_4 fanout451 (.A(_1739_),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_8 fanout452 (.A(_1738_),
    .X(net452));
 sky130_fd_sc_hd__buf_2 fanout453 (.A(_1738_),
    .X(net453));
 sky130_fd_sc_hd__buf_8 fanout454 (.A(_1509_),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_4 fanout455 (.A(_1509_),
    .X(net455));
 sky130_fd_sc_hd__buf_6 fanout456 (.A(_1508_),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_4 fanout457 (.A(_1508_),
    .X(net457));
 sky130_fd_sc_hd__buf_6 fanout461 (.A(net464),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_8 fanout462 (.A(net464),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_4 fanout463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__buf_4 fanout464 (.A(_1731_),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_8 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_4 fanout466 (.A(_1730_),
    .X(net466));
 sky130_fd_sc_hd__buf_6 fanout467 (.A(_1730_),
    .X(net467));
 sky130_fd_sc_hd__buf_4 fanout468 (.A(_1730_),
    .X(net468));
 sky130_fd_sc_hd__buf_4 fanout469 (.A(net472),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_8 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_6 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_6 fanout472 (.A(_1727_),
    .X(net472));
 sky130_fd_sc_hd__buf_6 fanout473 (.A(net475),
    .X(net473));
 sky130_fd_sc_hd__buf_6 fanout474 (.A(net475),
    .X(net474));
 sky130_fd_sc_hd__buf_6 fanout475 (.A(_1504_),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_8 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_4 fanout477 (.A(net479),
    .X(net477));
 sky130_fd_sc_hd__buf_6 fanout478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_8 fanout479 (.A(_1503_),
    .X(net479));
 sky130_fd_sc_hd__buf_6 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_6 fanout481 (.A(net483),
    .X(net481));
 sky130_fd_sc_hd__buf_6 fanout482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__buf_4 fanout483 (.A(_1500_),
    .X(net483));
 sky130_fd_sc_hd__buf_6 fanout484 (.A(net486),
    .X(net484));
 sky130_fd_sc_hd__buf_4 fanout485 (.A(net1282),
    .X(net485));
 sky130_fd_sc_hd__buf_8 fanout486 (.A(_1404_),
    .X(net486));
 sky130_fd_sc_hd__buf_6 fanout487 (.A(_1404_),
    .X(net487));
 sky130_fd_sc_hd__buf_2 fanout488 (.A(_1404_),
    .X(net488));
 sky130_fd_sc_hd__buf_8 fanout489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_8 fanout490 (.A(net1629),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_8 fanout491 (.A(net1629),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_4 fanout492 (.A(net1645),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_8 fanout493 (.A(net496),
    .X(net493));
 sky130_fd_sc_hd__buf_6 fanout494 (.A(net495),
    .X(net494));
 sky130_fd_sc_hd__buf_6 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__buf_6 fanout496 (.A(_1726_),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_8 fanout497 (.A(_1502_),
    .X(net497));
 sky130_fd_sc_hd__buf_6 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_6 fanout499 (.A(net501),
    .X(net499));
 sky130_fd_sc_hd__buf_6 fanout500 (.A(net501),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_8 fanout501 (.A(_1499_),
    .X(net501));
 sky130_fd_sc_hd__buf_8 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__buf_12 fanout503 (.A(net506),
    .X(net503));
 sky130_fd_sc_hd__buf_8 fanout504 (.A(net506),
    .X(net504));
 sky130_fd_sc_hd__buf_6 fanout505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__buf_12 fanout506 (.A(_1403_),
    .X(net506));
 sky130_fd_sc_hd__buf_4 fanout507 (.A(_1397_),
    .X(net507));
 sky130_fd_sc_hd__buf_6 fanout508 (.A(_1396_),
    .X(net508));
 sky130_fd_sc_hd__buf_4 fanout509 (.A(_1396_),
    .X(net509));
 sky130_fd_sc_hd__buf_8 fanout510 (.A(_1371_),
    .X(net510));
 sky130_fd_sc_hd__buf_6 fanout511 (.A(\device.rxBuffer.endPointer[3] ),
    .X(net511));
 sky130_fd_sc_hd__buf_12 fanout512 (.A(\device.rxBuffer.endPointer[2] ),
    .X(net512));
 sky130_fd_sc_hd__buf_8 fanout513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__buf_8 fanout514 (.A(\device.rxBuffer.startPointer[2] ),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_16 fanout515 (.A(net517),
    .X(net515));
 sky130_fd_sc_hd__buf_4 fanout516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__buf_12 fanout517 (.A(\device.rxBuffer.startPointer[1] ),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_16 fanout518 (.A(\device.rxBuffer.startPointer[1] ),
    .X(net518));
 sky130_fd_sc_hd__buf_4 fanout519 (.A(\device.rxBuffer.startPointer[1] ),
    .X(net519));
 sky130_fd_sc_hd__buf_6 fanout520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__buf_6 fanout521 (.A(net524),
    .X(net521));
 sky130_fd_sc_hd__buf_6 fanout522 (.A(net524),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_16 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_8 fanout524 (.A(\device.rxBuffer.startPointer[0] ),
    .X(net524));
 sky130_fd_sc_hd__buf_6 fanout525 (.A(net528),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_16 fanout526 (.A(net528),
    .X(net526));
 sky130_fd_sc_hd__buf_6 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__buf_6 fanout528 (.A(\device.rxBuffer.startPointer[0] ),
    .X(net528));
 sky130_fd_sc_hd__buf_6 fanout529 (.A(\device.txBuffer.endPointer[2] ),
    .X(net529));
 sky130_fd_sc_hd__buf_6 fanout530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__buf_8 fanout531 (.A(\device.txBuffer.startPointer[2] ),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_16 fanout532 (.A(net533),
    .X(net532));
 sky130_fd_sc_hd__buf_4 fanout533 (.A(net537),
    .X(net533));
 sky130_fd_sc_hd__buf_8 fanout534 (.A(net537),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_4 fanout535 (.A(net537),
    .X(net535));
 sky130_fd_sc_hd__buf_8 fanout536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__buf_6 fanout537 (.A(\device.txBuffer.startPointer[1] ),
    .X(net537));
 sky130_fd_sc_hd__buf_6 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_6 fanout539 (.A(net540),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_16 fanout540 (.A(\device.txBuffer.startPointer[0] ),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_16 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__buf_6 fanout542 (.A(net547),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_16 fanout543 (.A(net547),
    .X(net543));
 sky130_fd_sc_hd__buf_4 fanout544 (.A(net547),
    .X(net544));
 sky130_fd_sc_hd__buf_8 fanout545 (.A(net547),
    .X(net545));
 sky130_fd_sc_hd__buf_4 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__buf_6 fanout547 (.A(\device.txBuffer.startPointer[0] ),
    .X(net547));
 sky130_fd_sc_hd__buf_4 fanout548 (.A(_2367_),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_4 fanout549 (.A(_2367_),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_8 fanout550 (.A(_2214_),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_4 fanout551 (.A(_2214_),
    .X(net551));
 sky130_fd_sc_hd__buf_6 fanout552 (.A(_2133_),
    .X(net552));
 sky130_fd_sc_hd__buf_6 fanout553 (.A(net557),
    .X(net553));
 sky130_fd_sc_hd__buf_4 fanout554 (.A(net557),
    .X(net554));
 sky130_fd_sc_hd__buf_6 fanout555 (.A(net557),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_4 fanout556 (.A(net557),
    .X(net556));
 sky130_fd_sc_hd__buf_8 fanout557 (.A(_2034_),
    .X(net557));
 sky130_fd_sc_hd__buf_4 fanout558 (.A(net559),
    .X(net558));
 sky130_fd_sc_hd__buf_6 fanout559 (.A(_1407_),
    .X(net559));
 sky130_fd_sc_hd__buf_4 fanout560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_4 fanout561 (.A(\device.txBuffer.dataIn_buffered[7] ),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_8 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__buf_4 fanout563 (.A(\device.txBuffer.dataIn_buffered[7] ),
    .X(net563));
 sky130_fd_sc_hd__buf_4 fanout564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_4 fanout565 (.A(\device.txBuffer.dataIn_buffered[6] ),
    .X(net565));
 sky130_fd_sc_hd__buf_6 fanout566 (.A(\device.txBuffer.dataIn_buffered[6] ),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_4 fanout567 (.A(\device.txBuffer.dataIn_buffered[6] ),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_8 fanout568 (.A(net571),
    .X(net568));
 sky130_fd_sc_hd__buf_4 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__buf_8 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__buf_6 fanout571 (.A(\device.txBuffer.dataIn_buffered[5] ),
    .X(net571));
 sky130_fd_sc_hd__buf_4 fanout572 (.A(\device.txBuffer.dataIn_buffered[4] ),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_8 fanout573 (.A(net575),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_2 fanout574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__buf_4 fanout575 (.A(\device.txBuffer.dataIn_buffered[4] ),
    .X(net575));
 sky130_fd_sc_hd__buf_4 fanout576 (.A(net579),
    .X(net576));
 sky130_fd_sc_hd__buf_4 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__buf_4 fanout578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__buf_6 fanout579 (.A(\device.txBuffer.dataIn_buffered[3] ),
    .X(net579));
 sky130_fd_sc_hd__buf_4 fanout580 (.A(\device.txBuffer.dataIn_buffered[2] ),
    .X(net580));
 sky130_fd_sc_hd__buf_4 fanout581 (.A(net583),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 fanout582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_4 fanout583 (.A(\device.txBuffer.dataIn_buffered[2] ),
    .X(net583));
 sky130_fd_sc_hd__buf_6 fanout584 (.A(\device.txBuffer.dataIn_buffered[1] ),
    .X(net584));
 sky130_fd_sc_hd__buf_4 fanout585 (.A(net587),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 fanout586 (.A(net587),
    .X(net586));
 sky130_fd_sc_hd__buf_4 fanout587 (.A(\device.txBuffer.dataIn_buffered[1] ),
    .X(net587));
 sky130_fd_sc_hd__buf_4 fanout588 (.A(\device.txBuffer.dataIn_buffered[0] ),
    .X(net588));
 sky130_fd_sc_hd__buf_4 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_4 fanout590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__buf_4 fanout591 (.A(\device.txBuffer.dataIn_buffered[0] ),
    .X(net591));
 sky130_fd_sc_hd__buf_4 fanout592 (.A(net596),
    .X(net592));
 sky130_fd_sc_hd__buf_2 fanout593 (.A(net596),
    .X(net593));
 sky130_fd_sc_hd__buf_4 fanout594 (.A(net596),
    .X(net594));
 sky130_fd_sc_hd__buf_2 fanout595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__buf_6 fanout596 (.A(\device.rxBuffer.dataIn_buffered[7] ),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_4 fanout597 (.A(net601),
    .X(net597));
 sky130_fd_sc_hd__buf_2 fanout598 (.A(net601),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_8 fanout599 (.A(net601),
    .X(net599));
 sky130_fd_sc_hd__buf_2 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__buf_6 fanout601 (.A(\device.rxBuffer.dataIn_buffered[6] ),
    .X(net601));
 sky130_fd_sc_hd__buf_4 fanout602 (.A(\device.rxBuffer.dataIn_buffered[5] ),
    .X(net602));
 sky130_fd_sc_hd__buf_2 fanout603 (.A(\device.rxBuffer.dataIn_buffered[5] ),
    .X(net603));
 sky130_fd_sc_hd__buf_4 fanout604 (.A(net605),
    .X(net604));
 sky130_fd_sc_hd__buf_2 fanout605 (.A(\device.rxBuffer.dataIn_buffered[5] ),
    .X(net605));
 sky130_fd_sc_hd__buf_4 fanout606 (.A(net609),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_2 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__buf_6 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__buf_8 fanout609 (.A(\device.rxBuffer.dataIn_buffered[4] ),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_4 fanout610 (.A(\device.rxBuffer.dataIn_buffered[3] ),
    .X(net610));
 sky130_fd_sc_hd__buf_2 fanout611 (.A(\device.rxBuffer.dataIn_buffered[3] ),
    .X(net611));
 sky130_fd_sc_hd__buf_4 fanout612 (.A(\device.rxBuffer.dataIn_buffered[3] ),
    .X(net612));
 sky130_fd_sc_hd__buf_2 fanout613 (.A(\device.rxBuffer.dataIn_buffered[3] ),
    .X(net613));
 sky130_fd_sc_hd__buf_4 fanout614 (.A(\device.rxBuffer.dataIn_buffered[2] ),
    .X(net614));
 sky130_fd_sc_hd__buf_2 fanout615 (.A(\device.rxBuffer.dataIn_buffered[2] ),
    .X(net615));
 sky130_fd_sc_hd__buf_4 fanout616 (.A(\device.rxBuffer.dataIn_buffered[2] ),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_2 fanout617 (.A(\device.rxBuffer.dataIn_buffered[2] ),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_4 fanout618 (.A(\device.rxBuffer.dataIn_buffered[1] ),
    .X(net618));
 sky130_fd_sc_hd__buf_2 fanout619 (.A(\device.rxBuffer.dataIn_buffered[1] ),
    .X(net619));
 sky130_fd_sc_hd__buf_4 fanout620 (.A(\device.rxBuffer.dataIn_buffered[1] ),
    .X(net620));
 sky130_fd_sc_hd__buf_2 fanout621 (.A(\device.rxBuffer.dataIn_buffered[1] ),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_4 fanout622 (.A(net624),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_4 fanout623 (.A(net624),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_4 fanout624 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__buf_4 fanout625 (.A(\device.rxBuffer.dataIn_buffered[0] ),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_8 fanout626 (.A(\wbPeripheralBusInterface.currentByteSelect[1] ),
    .X(net626));
 sky130_fd_sc_hd__buf_4 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__buf_6 fanout628 (.A(\wbPeripheralBusInterface.currentByteSelect[0] ),
    .X(net628));
 sky130_fd_sc_hd__buf_4 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__buf_6 fanout630 (.A(\wbPeripheralBusInterface.state[1] ),
    .X(net630));
 sky130_fd_sc_hd__buf_6 fanout631 (.A(\wbPeripheralBusInterface.state[0] ),
    .X(net631));
 sky130_fd_sc_hd__buf_4 fanout632 (.A(net1954),
    .X(net632));
 sky130_fd_sc_hd__buf_4 fanout633 (.A(net1990),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_8 fanout634 (.A(net1990),
    .X(net634));
 sky130_fd_sc_hd__buf_6 fanout635 (.A(net637),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_4 fanout636 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__buf_12 fanout637 (.A(_1373_),
    .X(net637));
 sky130_fd_sc_hd__buf_4 fanout638 (.A(net2924),
    .X(net638));
 sky130_fd_sc_hd__buf_6 fanout639 (.A(net141),
    .X(net639));
 sky130_fd_sc_hd__buf_6 fanout640 (.A(net141),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_8 fanout641 (.A(net141),
    .X(net641));
 sky130_fd_sc_hd__buf_12 fanout642 (.A(net1418),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_4 fanout643 (.A(net1418),
    .X(net643));
 sky130_fd_sc_hd__buf_8 fanout644 (.A(net1466),
    .X(net644));
 sky130_fd_sc_hd__buf_6 fanout645 (.A(net1483),
    .X(net645));
 sky130_fd_sc_hd__buf_2 fanout646 (.A(net1483),
    .X(net646));
 sky130_fd_sc_hd__buf_6 fanout647 (.A(net1466),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_8 fanout648 (.A(net1466),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_4 fanout649 (.A(net1466),
    .X(net649));
 sky130_fd_sc_hd__buf_12 fanout650 (.A(net134),
    .X(net650));
 sky130_fd_sc_hd__buf_2 hold10 (.A(net1374),
    .X(net1291));
 sky130_fd_sc_hd__buf_2 hold100 (.A(net1354),
    .X(net1381));
 sky130_fd_sc_hd__buf_2 hold1000 (.A(net2835),
    .X(net2281));
 sky130_fd_sc_hd__buf_2 hold1001 (.A(net2837),
    .X(net2282));
 sky130_fd_sc_hd__buf_2 hold1002 (.A(net2839),
    .X(net2283));
 sky130_fd_sc_hd__buf_2 hold1003 (.A(net3691),
    .X(net2284));
 sky130_fd_sc_hd__buf_2 hold1004 (.A(net3695),
    .X(net2285));
 sky130_fd_sc_hd__buf_2 hold1005 (.A(net3699),
    .X(net2286));
 sky130_fd_sc_hd__buf_2 hold1006 (.A(net2847),
    .X(net2287));
 sky130_fd_sc_hd__buf_2 hold1007 (.A(net2849),
    .X(net2288));
 sky130_fd_sc_hd__buf_2 hold1008 (.A(net2851),
    .X(net2289));
 sky130_fd_sc_hd__buf_2 hold1009 (.A(net3711),
    .X(net2290));
 sky130_fd_sc_hd__buf_2 hold101 (.A(net1355),
    .X(net1382));
 sky130_fd_sc_hd__buf_2 hold1010 (.A(net3715),
    .X(net2291));
 sky130_fd_sc_hd__buf_2 hold1011 (.A(net3719),
    .X(net2292));
 sky130_fd_sc_hd__buf_2 hold1012 (.A(net2859),
    .X(net2293));
 sky130_fd_sc_hd__buf_2 hold1013 (.A(net2861),
    .X(net2294));
 sky130_fd_sc_hd__buf_2 hold1014 (.A(net2863),
    .X(net2295));
 sky130_fd_sc_hd__buf_2 hold1015 (.A(net3739),
    .X(net2296));
 sky130_fd_sc_hd__buf_2 hold1016 (.A(net3743),
    .X(net2297));
 sky130_fd_sc_hd__buf_2 hold1017 (.A(net2881),
    .X(net2298));
 sky130_fd_sc_hd__buf_2 hold1018 (.A(net2883),
    .X(net2299));
 sky130_fd_sc_hd__buf_2 hold1019 (.A(net2885),
    .X(net2300));
 sky130_fd_sc_hd__buf_2 hold1020 (.A(net2887),
    .X(net2301));
 sky130_fd_sc_hd__buf_2 hold1021 (.A(net3721),
    .X(net2302));
 sky130_fd_sc_hd__buf_2 hold1022 (.A(net3725),
    .X(net2303));
 sky130_fd_sc_hd__buf_2 hold1023 (.A(net2869),
    .X(net2304));
 sky130_fd_sc_hd__buf_2 hold1024 (.A(net2871),
    .X(net2305));
 sky130_fd_sc_hd__buf_2 hold1025 (.A(net2873),
    .X(net2306));
 sky130_fd_sc_hd__buf_2 hold1026 (.A(net2875),
    .X(net2307));
 sky130_fd_sc_hd__buf_2 hold1027 (.A(net3730),
    .X(net2308));
 sky130_fd_sc_hd__buf_2 hold1028 (.A(net3734),
    .X(net2309));
 sky130_fd_sc_hd__buf_2 hold1029 (.A(net2893),
    .X(net2310));
 sky130_fd_sc_hd__buf_2 hold103 (.A(net1420),
    .X(net1384));
 sky130_fd_sc_hd__buf_2 hold1030 (.A(net2895),
    .X(net2311));
 sky130_fd_sc_hd__buf_2 hold1031 (.A(net2897),
    .X(net2312));
 sky130_fd_sc_hd__buf_2 hold1032 (.A(net2899),
    .X(net2313));
 sky130_fd_sc_hd__buf_2 hold1035 (.A(net4071),
    .X(net2316));
 sky130_fd_sc_hd__buf_2 hold1036 (.A(net1956),
    .X(net2317));
 sky130_fd_sc_hd__buf_2 hold1037 (.A(net3872),
    .X(net2318));
 sky130_fd_sc_hd__buf_2 hold1038 (.A(net3876),
    .X(net2319));
 sky130_fd_sc_hd__buf_2 hold1039 (.A(net2929),
    .X(net2320));
 sky130_fd_sc_hd__buf_2 hold104 (.A(net1422),
    .X(net1385));
 sky130_fd_sc_hd__buf_2 hold1040 (.A(net2931),
    .X(net2321));
 sky130_fd_sc_hd__buf_2 hold1041 (.A(net3139),
    .X(net2322));
 sky130_fd_sc_hd__buf_2 hold1042 (.A(net3141),
    .X(net2323));
 sky130_fd_sc_hd__buf_2 hold1043 (.A(net3143),
    .X(net2324));
 sky130_fd_sc_hd__buf_2 hold1044 (.A(net1476),
    .X(net2325));
 sky130_fd_sc_hd__buf_2 hold1045 (.A(net205),
    .X(net2326));
 sky130_fd_sc_hd__buf_2 hold1046 (.A(net1477),
    .X(net2327));
 sky130_fd_sc_hd__buf_2 hold1047 (.A(net1430),
    .X(net2328));
 sky130_fd_sc_hd__buf_2 hold1048 (.A(net1478),
    .X(net2329));
 sky130_fd_sc_hd__buf_2 hold1049 (.A(_2042_),
    .X(net2330));
 sky130_fd_sc_hd__buf_2 hold105 (.A(net1404),
    .X(net1386));
 sky130_fd_sc_hd__buf_2 hold1050 (.A(net1431),
    .X(net2331));
 sky130_fd_sc_hd__buf_2 hold1051 (.A(net3117),
    .X(net2332));
 sky130_fd_sc_hd__buf_2 hold1052 (.A(net3119),
    .X(net2333));
 sky130_fd_sc_hd__buf_2 hold1057 (.A(net2400),
    .X(net2338));
 sky130_fd_sc_hd__buf_2 hold1058 (.A(net2402),
    .X(net2339));
 sky130_fd_sc_hd__buf_2 hold1059 (.A(_2122_),
    .X(net2340));
 sky130_fd_sc_hd__buf_2 hold106 (.A(net1408),
    .X(net1387));
 sky130_fd_sc_hd__buf_2 hold1060 (.A(net3245),
    .X(net2341));
 sky130_fd_sc_hd__buf_2 hold1061 (.A(net3247),
    .X(net2342));
 sky130_fd_sc_hd__buf_2 hold1065 (.A(net3484),
    .X(net2346));
 sky130_fd_sc_hd__buf_2 hold1066 (.A(net3488),
    .X(net2347));
 sky130_fd_sc_hd__buf_2 hold1068 (.A(net4080),
    .X(net2349));
 sky130_fd_sc_hd__buf_2 hold1069 (.A(net3468),
    .X(net2350));
 sky130_fd_sc_hd__buf_2 hold107 (.A(net1412),
    .X(net1388));
 sky130_fd_sc_hd__buf_2 hold1072 (.A(net4021),
    .X(net2353));
 sky130_fd_sc_hd__buf_2 hold1073 (.A(net3113),
    .X(net2354));
 sky130_fd_sc_hd__buf_2 hold1074 (.A(net3115),
    .X(net2355));
 sky130_fd_sc_hd__buf_2 hold1075 (.A(net3145),
    .X(net2356));
 sky130_fd_sc_hd__buf_2 hold1076 (.A(net3147),
    .X(net2357));
 sky130_fd_sc_hd__buf_2 hold1078 (.A(net4087),
    .X(net2359));
 sky130_fd_sc_hd__buf_2 hold1079 (.A(net3477),
    .X(net2360));
 sky130_fd_sc_hd__buf_2 hold108 (.A(net1398),
    .X(net1389));
 sky130_fd_sc_hd__buf_2 hold1085 (.A(net3585),
    .X(net2366));
 sky130_fd_sc_hd__buf_2 hold1086 (.A(net3589),
    .X(net2367));
 sky130_fd_sc_hd__buf_2 hold109 (.A(net1416),
    .X(net1390));
 sky130_fd_sc_hd__buf_2 hold1092 (.A(net3598),
    .X(net2373));
 sky130_fd_sc_hd__buf_2 hold1093 (.A(net3602),
    .X(net2374));
 sky130_fd_sc_hd__buf_2 hold1099 (.A(net3647),
    .X(net2380));
 sky130_fd_sc_hd__buf_2 hold11 (.A(_1278_),
    .X(net1292));
 sky130_fd_sc_hd__buf_2 hold110 (.A(_1240_),
    .X(net1391));
 sky130_fd_sc_hd__buf_2 hold1100 (.A(net3651),
    .X(net2381));
 sky130_fd_sc_hd__buf_2 hold1106 (.A(net3621),
    .X(net2387));
 sky130_fd_sc_hd__buf_2 hold1107 (.A(net3625),
    .X(net2388));
 sky130_fd_sc_hd__buf_2 hold111 (.A(net1403),
    .X(net1392));
 sky130_fd_sc_hd__buf_2 hold1113 (.A(net3634),
    .X(net2394));
 sky130_fd_sc_hd__buf_2 hold1114 (.A(net3638),
    .X(net2395));
 sky130_fd_sc_hd__buf_2 hold1119 (.A(net4059),
    .X(net2400));
 sky130_fd_sc_hd__buf_2 hold112 (.A(net1405),
    .X(net1393));
 sky130_fd_sc_hd__buf_2 hold1120 (.A(net2338),
    .X(net2401));
 sky130_fd_sc_hd__buf_2 hold1121 (.A(net1479),
    .X(net2402));
 sky130_fd_sc_hd__buf_2 hold1122 (.A(net2339),
    .X(net2403));
 sky130_fd_sc_hd__buf_2 hold1123 (.A(_2125_),
    .X(net2404));
 sky130_fd_sc_hd__buf_2 hold1124 (.A(net1480),
    .X(net2405));
 sky130_fd_sc_hd__buf_2 hold1125 (.A(net3331),
    .X(net2406));
 sky130_fd_sc_hd__buf_2 hold1126 (.A(net3333),
    .X(net2407));
 sky130_fd_sc_hd__buf_2 hold113 (.A(net1407),
    .X(net1394));
 sky130_fd_sc_hd__buf_2 hold1132 (.A(net3660),
    .X(net2413));
 sky130_fd_sc_hd__buf_2 hold1133 (.A(net3664),
    .X(net2414));
 sky130_fd_sc_hd__buf_2 hold1139 (.A(net3683),
    .X(net2420));
 sky130_fd_sc_hd__buf_2 hold114 (.A(net1409),
    .X(net1395));
 sky130_fd_sc_hd__buf_2 hold1140 (.A(net3687),
    .X(net2421));
 sky130_fd_sc_hd__buf_2 hold115 (.A(net1411),
    .X(net1396));
 sky130_fd_sc_hd__buf_2 hold1151 (.A(net3496),
    .X(net2432));
 sky130_fd_sc_hd__buf_2 hold1152 (.A(net3500),
    .X(net2433));
 sky130_fd_sc_hd__buf_2 hold1157 (.A(net3508),
    .X(net2438));
 sky130_fd_sc_hd__buf_2 hold1158 (.A(net3512),
    .X(net2439));
 sky130_fd_sc_hd__buf_2 hold116 (.A(net1413),
    .X(net1397));
 sky130_fd_sc_hd__buf_2 hold1162 (.A(net4012),
    .X(net2443));
 sky130_fd_sc_hd__buf_2 hold1163 (.A(net3103),
    .X(net2444));
 sky130_fd_sc_hd__buf_2 hold1164 (.A(net3105),
    .X(net2445));
 sky130_fd_sc_hd__buf_2 hold1165 (.A(net3107),
    .X(net2446));
 sky130_fd_sc_hd__buf_2 hold1169 (.A(net4017),
    .X(net2450));
 sky130_fd_sc_hd__buf_2 hold117 (.A(net1333),
    .X(net1398));
 sky130_fd_sc_hd__buf_2 hold1170 (.A(net3126),
    .X(net2451));
 sky130_fd_sc_hd__buf_2 hold1171 (.A(net3128),
    .X(net2452));
 sky130_fd_sc_hd__buf_2 hold1172 (.A(net3130),
    .X(net2453));
 sky130_fd_sc_hd__buf_2 hold1176 (.A(net3152),
    .X(net2457));
 sky130_fd_sc_hd__buf_2 hold1177 (.A(net3154),
    .X(net2458));
 sky130_fd_sc_hd__buf_2 hold1178 (.A(net3156),
    .X(net2459));
 sky130_fd_sc_hd__buf_2 hold1179 (.A(net3158),
    .X(net2460));
 sky130_fd_sc_hd__buf_2 hold118 (.A(net1389),
    .X(net1399));
 sky130_fd_sc_hd__buf_2 hold1185 (.A(net3831),
    .X(net2466));
 sky130_fd_sc_hd__buf_2 hold1186 (.A(net3835),
    .X(net2467));
 sky130_fd_sc_hd__buf_2 hold119 (.A(net1415),
    .X(net1400));
 sky130_fd_sc_hd__buf_2 hold1192 (.A(net3844),
    .X(net2473));
 sky130_fd_sc_hd__buf_2 hold1193 (.A(net3848),
    .X(net2474));
 sky130_fd_sc_hd__buf_2 hold1197 (.A(net3185),
    .X(net2478));
 sky130_fd_sc_hd__buf_2 hold1198 (.A(net3187),
    .X(net2479));
 sky130_fd_sc_hd__buf_2 hold1199 (.A(net3189),
    .X(net2480));
 sky130_fd_sc_hd__buf_2 hold12 (.A(net3518),
    .X(net1293));
 sky130_fd_sc_hd__buf_2 hold120 (.A(net1390),
    .X(net1401));
 sky130_fd_sc_hd__buf_2 hold1200 (.A(net3191),
    .X(net2481));
 sky130_fd_sc_hd__buf_2 hold1204 (.A(net3174),
    .X(net2485));
 sky130_fd_sc_hd__buf_2 hold1205 (.A(net3176),
    .X(net2486));
 sky130_fd_sc_hd__buf_2 hold1206 (.A(net3178),
    .X(net2487));
 sky130_fd_sc_hd__buf_2 hold1207 (.A(net3180),
    .X(net2488));
 sky130_fd_sc_hd__buf_2 hold121 (.A(_1239_),
    .X(net1402));
 sky130_fd_sc_hd__buf_2 hold1211 (.A(net3196),
    .X(net2492));
 sky130_fd_sc_hd__buf_2 hold1212 (.A(net3198),
    .X(net2493));
 sky130_fd_sc_hd__buf_2 hold1213 (.A(net3200),
    .X(net2494));
 sky130_fd_sc_hd__buf_2 hold1214 (.A(net3202),
    .X(net2495));
 sky130_fd_sc_hd__buf_2 hold1218 (.A(net3163),
    .X(net2499));
 sky130_fd_sc_hd__buf_2 hold1219 (.A(net3165),
    .X(net2500));
 sky130_fd_sc_hd__buf_2 hold122 (.A(wbs_sel_i[2]),
    .X(net1403));
 sky130_fd_sc_hd__buf_2 hold1220 (.A(net3167),
    .X(net2501));
 sky130_fd_sc_hd__buf_2 hold1221 (.A(net3169),
    .X(net2502));
 sky130_fd_sc_hd__buf_2 hold1225 (.A(net3207),
    .X(net2506));
 sky130_fd_sc_hd__buf_2 hold1226 (.A(net3209),
    .X(net2507));
 sky130_fd_sc_hd__buf_2 hold1227 (.A(net3211),
    .X(net2508));
 sky130_fd_sc_hd__buf_2 hold1228 (.A(net3213),
    .X(net2509));
 sky130_fd_sc_hd__buf_2 hold123 (.A(net1392),
    .X(net1404));
 sky130_fd_sc_hd__buf_2 hold1232 (.A(net3218),
    .X(net2513));
 sky130_fd_sc_hd__buf_2 hold1233 (.A(net3220),
    .X(net2514));
 sky130_fd_sc_hd__buf_2 hold1234 (.A(net3222),
    .X(net2515));
 sky130_fd_sc_hd__buf_2 hold1235 (.A(net3224),
    .X(net2516));
 sky130_fd_sc_hd__buf_2 hold1239 (.A(net3229),
    .X(net2520));
 sky130_fd_sc_hd__buf_2 hold124 (.A(net1386),
    .X(net1405));
 sky130_fd_sc_hd__buf_2 hold1240 (.A(net3231),
    .X(net2521));
 sky130_fd_sc_hd__buf_2 hold1241 (.A(net3233),
    .X(net2522));
 sky130_fd_sc_hd__buf_2 hold1242 (.A(net3235),
    .X(net2523));
 sky130_fd_sc_hd__buf_2 hold1247 (.A(net3562),
    .X(net2528));
 sky130_fd_sc_hd__buf_2 hold1248 (.A(net3566),
    .X(net2529));
 sky130_fd_sc_hd__buf_2 hold125 (.A(net1393),
    .X(net1406));
 sky130_fd_sc_hd__buf_2 hold1254 (.A(net3753),
    .X(net2535));
 sky130_fd_sc_hd__buf_2 hold1255 (.A(net3757),
    .X(net2536));
 sky130_fd_sc_hd__buf_2 hold126 (.A(net1332),
    .X(net1407));
 sky130_fd_sc_hd__buf_2 hold1261 (.A(net3766),
    .X(net2542));
 sky130_fd_sc_hd__buf_2 hold1262 (.A(net3770),
    .X(net2543));
 sky130_fd_sc_hd__buf_2 hold1268 (.A(net3779),
    .X(net2549));
 sky130_fd_sc_hd__buf_2 hold1269 (.A(net3783),
    .X(net2550));
 sky130_fd_sc_hd__buf_2 hold127 (.A(net1394),
    .X(net1408));
 sky130_fd_sc_hd__buf_2 hold1275 (.A(net3805),
    .X(net2556));
 sky130_fd_sc_hd__buf_2 hold1276 (.A(net3809),
    .X(net2557));
 sky130_fd_sc_hd__buf_2 hold128 (.A(net1387),
    .X(net1409));
 sky130_fd_sc_hd__buf_2 hold1282 (.A(net3792),
    .X(net2563));
 sky130_fd_sc_hd__buf_2 hold1283 (.A(net3796),
    .X(net2564));
 sky130_fd_sc_hd__buf_2 hold1289 (.A(net3818),
    .X(net2570));
 sky130_fd_sc_hd__buf_2 hold129 (.A(net1395),
    .X(net1410));
 sky130_fd_sc_hd__buf_2 hold1290 (.A(net3822),
    .X(net2571));
 sky130_fd_sc_hd__buf_2 hold1293 (.A(net3854),
    .X(net2574));
 sky130_fd_sc_hd__buf_2 hold1294 (.A(net3858),
    .X(net2575));
 sky130_fd_sc_hd__buf_2 hold1298 (.A(net3865),
    .X(net2579));
 sky130_fd_sc_hd__buf_2 hold1299 (.A(net3869),
    .X(net2580));
 sky130_fd_sc_hd__buf_2 hold13 (.A(net2750),
    .X(net1294));
 sky130_fd_sc_hd__buf_2 hold130 (.A(net202),
    .X(net1411));
 sky130_fd_sc_hd__buf_2 hold1303 (.A(_2418_),
    .X(net2584));
 sky130_fd_sc_hd__buf_2 hold1304 (.A(net1739),
    .X(net2585));
 sky130_fd_sc_hd__buf_2 hold1305 (.A(net3907),
    .X(net2586));
 sky130_fd_sc_hd__buf_2 hold1306 (.A(net3911),
    .X(net2587));
 sky130_fd_sc_hd__buf_2 hold131 (.A(net1396),
    .X(net1412));
 sky130_fd_sc_hd__buf_2 hold1314 (.A(net3886),
    .X(net2595));
 sky130_fd_sc_hd__buf_2 hold1315 (.A(net3890),
    .X(net2596));
 sky130_fd_sc_hd__buf_2 hold132 (.A(net1388),
    .X(net1413));
 sky130_fd_sc_hd__buf_2 hold1323 (.A(net3899),
    .X(net2604));
 sky130_fd_sc_hd__buf_2 hold1324 (.A(net3903),
    .X(net2605));
 sky130_fd_sc_hd__buf_2 hold1327 (.A(net3915),
    .X(net2608));
 sky130_fd_sc_hd__buf_2 hold1328 (.A(net3919),
    .X(net2609));
 sky130_fd_sc_hd__buf_2 hold133 (.A(net1397),
    .X(net1414));
 sky130_fd_sc_hd__buf_2 hold1331 (.A(net3923),
    .X(net2612));
 sky130_fd_sc_hd__buf_2 hold1332 (.A(net3927),
    .X(net2613));
 sky130_fd_sc_hd__buf_2 hold1335 (.A(net3944),
    .X(net2616));
 sky130_fd_sc_hd__buf_2 hold1336 (.A(net3948),
    .X(net2617));
 sky130_fd_sc_hd__buf_2 hold1339 (.A(net3952),
    .X(net2620));
 sky130_fd_sc_hd__buf_2 hold134 (.A(_2127_),
    .X(net1415));
 sky130_fd_sc_hd__buf_2 hold1340 (.A(net3956),
    .X(net2621));
 sky130_fd_sc_hd__buf_2 hold1343 (.A(net3960),
    .X(net2624));
 sky130_fd_sc_hd__buf_2 hold1344 (.A(net3964),
    .X(net2625));
 sky130_fd_sc_hd__buf_2 hold135 (.A(net1400),
    .X(net1416));
 sky130_fd_sc_hd__buf_2 hold1352 (.A(net3936),
    .X(net2633));
 sky130_fd_sc_hd__buf_2 hold1353 (.A(net3940),
    .X(net2634));
 sky130_fd_sc_hd__buf_2 hold1356 (.A(net3968),
    .X(net2637));
 sky130_fd_sc_hd__buf_2 hold1357 (.A(net3972),
    .X(net2638));
 sky130_fd_sc_hd__buf_2 hold136 (.A(net1381),
    .X(net1417));
 sky130_fd_sc_hd__buf_2 hold1360 (.A(net3976),
    .X(net2641));
 sky130_fd_sc_hd__buf_2 hold1361 (.A(net3339),
    .X(net2642));
 sky130_fd_sc_hd__buf_2 hold1365 (.A(net3397),
    .X(net2646));
 sky130_fd_sc_hd__buf_2 hold1366 (.A(net3399),
    .X(net2647));
 sky130_fd_sc_hd__buf_2 hold1367 (.A(net3401),
    .X(net2648));
 sky130_fd_sc_hd__buf_2 hold1368 (.A(net1770),
    .X(net2649));
 sky130_fd_sc_hd__buf_2 hold137 (.A(net1382),
    .X(net1418));
 sky130_fd_sc_hd__buf_2 hold1372 (.A(net3406),
    .X(net2653));
 sky130_fd_sc_hd__buf_2 hold1373 (.A(net3408),
    .X(net2654));
 sky130_fd_sc_hd__buf_2 hold1374 (.A(net3410),
    .X(net2655));
 sky130_fd_sc_hd__buf_2 hold1375 (.A(net1775),
    .X(net2656));
 sky130_fd_sc_hd__buf_2 hold1379 (.A(net3415),
    .X(net2660));
 sky130_fd_sc_hd__buf_2 hold1380 (.A(net3417),
    .X(net2661));
 sky130_fd_sc_hd__buf_2 hold1381 (.A(net3419),
    .X(net2662));
 sky130_fd_sc_hd__buf_2 hold1382 (.A(net1803),
    .X(net2663));
 sky130_fd_sc_hd__buf_2 hold1386 (.A(net3424),
    .X(net2667));
 sky130_fd_sc_hd__buf_2 hold1387 (.A(net3426),
    .X(net2668));
 sky130_fd_sc_hd__buf_2 hold1388 (.A(net3428),
    .X(net2669));
 sky130_fd_sc_hd__buf_2 hold1389 (.A(net1823),
    .X(net2670));
 sky130_fd_sc_hd__buf_2 hold139 (.A(_2036_),
    .X(net1420));
 sky130_fd_sc_hd__buf_2 hold1393 (.A(net3433),
    .X(net2674));
 sky130_fd_sc_hd__buf_2 hold1394 (.A(net3435),
    .X(net2675));
 sky130_fd_sc_hd__buf_2 hold1395 (.A(net3437),
    .X(net2676));
 sky130_fd_sc_hd__buf_2 hold1396 (.A(net1842),
    .X(net2677));
 sky130_fd_sc_hd__buf_2 hold14 (.A(net2754),
    .X(net1295));
 sky130_fd_sc_hd__buf_2 hold140 (.A(net1384),
    .X(net1421));
 sky130_fd_sc_hd__buf_2 hold1402 (.A(net3444),
    .X(net2683));
 sky130_fd_sc_hd__buf_2 hold1403 (.A(net3446),
    .X(net2684));
 sky130_fd_sc_hd__buf_2 hold1404 (.A(net3448),
    .X(net2685));
 sky130_fd_sc_hd__buf_2 hold1405 (.A(net2235),
    .X(net2686));
 sky130_fd_sc_hd__buf_2 hold141 (.A(net1357),
    .X(net1422));
 sky130_fd_sc_hd__buf_2 hold1413 (.A(net3988),
    .X(net2694));
 sky130_fd_sc_hd__buf_2 hold1414 (.A(net3350),
    .X(net2695));
 sky130_fd_sc_hd__buf_2 hold1418 (.A(net3995),
    .X(net2699));
 sky130_fd_sc_hd__buf_2 hold1419 (.A(net3357),
    .X(net2700));
 sky130_fd_sc_hd__buf_2 hold142 (.A(net1445),
    .X(net1423));
 sky130_fd_sc_hd__buf_2 hold1423 (.A(net3362),
    .X(net2704));
 sky130_fd_sc_hd__buf_2 hold1424 (.A(net3364),
    .X(net2705));
 sky130_fd_sc_hd__buf_2 hold1428 (.A(net3369),
    .X(net2709));
 sky130_fd_sc_hd__buf_2 hold1429 (.A(net3371),
    .X(net2710));
 sky130_fd_sc_hd__buf_2 hold143 (.A(net1449),
    .X(net1424));
 sky130_fd_sc_hd__buf_2 hold1433 (.A(net3376),
    .X(net2714));
 sky130_fd_sc_hd__buf_2 hold1434 (.A(net3378),
    .X(net2715));
 sky130_fd_sc_hd__buf_2 hold1438 (.A(net3383),
    .X(net2719));
 sky130_fd_sc_hd__buf_2 hold1439 (.A(net3385),
    .X(net2720));
 sky130_fd_sc_hd__buf_2 hold144 (.A(net1453),
    .X(net1425));
 sky130_fd_sc_hd__buf_2 hold1443 (.A(net3390),
    .X(net2724));
 sky130_fd_sc_hd__buf_2 hold1444 (.A(net3392),
    .X(net2725));
 sky130_fd_sc_hd__buf_2 hold1447 (.A(net2736),
    .X(net2728));
 sky130_fd_sc_hd__buf_2 hold1448 (.A(net1733),
    .X(net2729));
 sky130_fd_sc_hd__buf_2 hold1449 (.A(net1696),
    .X(net2730));
 sky130_fd_sc_hd__buf_2 hold145 (.A(net1457),
    .X(net1426));
 sky130_fd_sc_hd__buf_2 hold1450 (.A(net1734),
    .X(net2731));
 sky130_fd_sc_hd__buf_2 hold1451 (.A(_1101_),
    .X(net2732));
 sky130_fd_sc_hd__buf_2 hold1452 (.A(net1697),
    .X(net2733));
 sky130_fd_sc_hd__buf_2 hold1455 (.A(net2740),
    .X(net2736));
 sky130_fd_sc_hd__buf_2 hold1456 (.A(net2728),
    .X(net2737));
 sky130_fd_sc_hd__buf_2 hold1459 (.A(net643),
    .X(net2740));
 sky130_fd_sc_hd__buf_2 hold146 (.A(net1441),
    .X(net1427));
 sky130_fd_sc_hd__buf_2 hold1462 (.A(net4168),
    .X(net2743));
 sky130_fd_sc_hd__buf_2 hold1463 (.A(net4073),
    .X(net2744));
 sky130_fd_sc_hd__buf_2 hold1464 (.A(net3515),
    .X(net2745));
 sky130_fd_sc_hd__buf_2 hold1465 (.A(net3517),
    .X(net2746));
 sky130_fd_sc_hd__buf_2 hold1466 (.A(net3519),
    .X(net2747));
 sky130_fd_sc_hd__buf_2 hold1467 (.A(net3521),
    .X(net2748));
 sky130_fd_sc_hd__buf_2 hold1468 (.A(net3523),
    .X(net2749));
 sky130_fd_sc_hd__buf_2 hold1469 (.A(net3525),
    .X(net2750));
 sky130_fd_sc_hd__buf_2 hold147 (.A(_1236_),
    .X(net1428));
 sky130_fd_sc_hd__buf_2 hold1470 (.A(net1294),
    .X(net2751));
 sky130_fd_sc_hd__buf_2 hold1471 (.A(net2239),
    .X(net2752));
 sky130_fd_sc_hd__buf_2 hold1472 (.A(_1079_),
    .X(net2753));
 sky130_fd_sc_hd__buf_2 hold1473 (.A(net2240),
    .X(net2754));
 sky130_fd_sc_hd__buf_2 hold1474 (.A(net1295),
    .X(net2755));
 sky130_fd_sc_hd__buf_2 hold1475 (.A(net2241),
    .X(net2756));
 sky130_fd_sc_hd__buf_2 hold1476 (.A(net3526),
    .X(net2757));
 sky130_fd_sc_hd__buf_2 hold1477 (.A(net3528),
    .X(net2758));
 sky130_fd_sc_hd__buf_2 hold1478 (.A(net3530),
    .X(net2759));
 sky130_fd_sc_hd__buf_2 hold1479 (.A(net3532),
    .X(net2760));
 sky130_fd_sc_hd__buf_2 hold148 (.A(net3142),
    .X(net1429));
 sky130_fd_sc_hd__buf_2 hold1480 (.A(net3534),
    .X(net2761));
 sky130_fd_sc_hd__buf_2 hold1481 (.A(net3536),
    .X(net2762));
 sky130_fd_sc_hd__buf_2 hold1482 (.A(net1300),
    .X(net2763));
 sky130_fd_sc_hd__buf_2 hold1483 (.A(net2245),
    .X(net2764));
 sky130_fd_sc_hd__buf_2 hold1484 (.A(_1080_),
    .X(net2765));
 sky130_fd_sc_hd__buf_2 hold1485 (.A(net2246),
    .X(net2766));
 sky130_fd_sc_hd__buf_2 hold1486 (.A(net1301),
    .X(net2767));
 sky130_fd_sc_hd__buf_2 hold1487 (.A(net2247),
    .X(net2768));
 sky130_fd_sc_hd__buf_2 hold1488 (.A(net3537),
    .X(net2769));
 sky130_fd_sc_hd__buf_2 hold1489 (.A(net3539),
    .X(net2770));
 sky130_fd_sc_hd__buf_2 hold149 (.A(net2327),
    .X(net1430));
 sky130_fd_sc_hd__buf_2 hold1490 (.A(net3541),
    .X(net2771));
 sky130_fd_sc_hd__buf_2 hold1491 (.A(net3543),
    .X(net2772));
 sky130_fd_sc_hd__buf_2 hold1492 (.A(net3545),
    .X(net2773));
 sky130_fd_sc_hd__buf_2 hold1493 (.A(net2250),
    .X(net2774));
 sky130_fd_sc_hd__buf_2 hold1494 (.A(net1306),
    .X(net2775));
 sky130_fd_sc_hd__buf_2 hold1495 (.A(net2251),
    .X(net2776));
 sky130_fd_sc_hd__buf_2 hold1496 (.A(_1081_),
    .X(net2777));
 sky130_fd_sc_hd__buf_2 hold1497 (.A(net2252),
    .X(net2778));
 sky130_fd_sc_hd__buf_2 hold1498 (.A(net1307),
    .X(net2779));
 sky130_fd_sc_hd__buf_2 hold1499 (.A(net2253),
    .X(net2780));
 sky130_fd_sc_hd__buf_2 hold15 (.A(net3703),
    .X(net1296));
 sky130_fd_sc_hd__buf_2 hold150 (.A(net2330),
    .X(net1431));
 sky130_fd_sc_hd__buf_2 hold1500 (.A(net3547),
    .X(net2781));
 sky130_fd_sc_hd__buf_2 hold1501 (.A(net3549),
    .X(net2782));
 sky130_fd_sc_hd__buf_2 hold1502 (.A(net3551),
    .X(net2783));
 sky130_fd_sc_hd__buf_2 hold1503 (.A(net3553),
    .X(net2784));
 sky130_fd_sc_hd__buf_2 hold1504 (.A(net3555),
    .X(net2785));
 sky130_fd_sc_hd__buf_2 hold1505 (.A(net2256),
    .X(net2786));
 sky130_fd_sc_hd__buf_2 hold1506 (.A(net1312),
    .X(net2787));
 sky130_fd_sc_hd__buf_2 hold1507 (.A(net2257),
    .X(net2788));
 sky130_fd_sc_hd__buf_2 hold1508 (.A(_1082_),
    .X(net2789));
 sky130_fd_sc_hd__buf_2 hold1509 (.A(net2258),
    .X(net2790));
 sky130_fd_sc_hd__buf_2 hold151 (.A(net3118),
    .X(net1432));
 sky130_fd_sc_hd__buf_2 hold1510 (.A(net1313),
    .X(net2791));
 sky130_fd_sc_hd__buf_2 hold1511 (.A(net2259),
    .X(net2792));
 sky130_fd_sc_hd__buf_2 hold1512 (.A(net3569),
    .X(net2793));
 sky130_fd_sc_hd__buf_2 hold1513 (.A(net3571),
    .X(net2794));
 sky130_fd_sc_hd__buf_2 hold1514 (.A(net3573),
    .X(net2795));
 sky130_fd_sc_hd__buf_2 hold1515 (.A(net3575),
    .X(net2796));
 sky130_fd_sc_hd__buf_2 hold1516 (.A(net3577),
    .X(net2797));
 sky130_fd_sc_hd__buf_2 hold1517 (.A(net2262),
    .X(net2798));
 sky130_fd_sc_hd__buf_2 hold1518 (.A(net1309),
    .X(net2799));
 sky130_fd_sc_hd__buf_2 hold1519 (.A(net2263),
    .X(net2800));
 sky130_fd_sc_hd__buf_2 hold152 (.A(net1444),
    .X(net1433));
 sky130_fd_sc_hd__buf_2 hold1520 (.A(_1083_),
    .X(net2801));
 sky130_fd_sc_hd__buf_2 hold1521 (.A(net2264),
    .X(net2802));
 sky130_fd_sc_hd__buf_2 hold1522 (.A(net1310),
    .X(net2803));
 sky130_fd_sc_hd__buf_2 hold1523 (.A(net2265),
    .X(net2804));
 sky130_fd_sc_hd__buf_2 hold1524 (.A(net3605),
    .X(net2805));
 sky130_fd_sc_hd__buf_2 hold1525 (.A(net3607),
    .X(net2806));
 sky130_fd_sc_hd__buf_2 hold1526 (.A(net3609),
    .X(net2807));
 sky130_fd_sc_hd__buf_2 hold1527 (.A(net3611),
    .X(net2808));
 sky130_fd_sc_hd__buf_2 hold1528 (.A(net3613),
    .X(net2809));
 sky130_fd_sc_hd__buf_2 hold1529 (.A(net2274),
    .X(net2810));
 sky130_fd_sc_hd__buf_2 hold153 (.A(net1446),
    .X(net1434));
 sky130_fd_sc_hd__buf_2 hold1530 (.A(net1318),
    .X(net2811));
 sky130_fd_sc_hd__buf_2 hold1531 (.A(net2275),
    .X(net2812));
 sky130_fd_sc_hd__buf_2 hold1532 (.A(_1084_),
    .X(net2813));
 sky130_fd_sc_hd__buf_2 hold1533 (.A(net2276),
    .X(net2814));
 sky130_fd_sc_hd__buf_2 hold1534 (.A(net1319),
    .X(net2815));
 sky130_fd_sc_hd__buf_2 hold1535 (.A(net2277),
    .X(net2816));
 sky130_fd_sc_hd__buf_2 hold1536 (.A(net3667),
    .X(net2817));
 sky130_fd_sc_hd__buf_2 hold1537 (.A(net3669),
    .X(net2818));
 sky130_fd_sc_hd__buf_2 hold1538 (.A(net3671),
    .X(net2819));
 sky130_fd_sc_hd__buf_2 hold1539 (.A(net3673),
    .X(net2820));
 sky130_fd_sc_hd__buf_2 hold154 (.A(net1448),
    .X(net1435));
 sky130_fd_sc_hd__buf_2 hold1540 (.A(net3675),
    .X(net2821));
 sky130_fd_sc_hd__buf_2 hold1541 (.A(net2268),
    .X(net2822));
 sky130_fd_sc_hd__buf_2 hold1542 (.A(net1288),
    .X(net2823));
 sky130_fd_sc_hd__buf_2 hold1543 (.A(net2269),
    .X(net2824));
 sky130_fd_sc_hd__buf_2 hold1544 (.A(_1085_),
    .X(net2825));
 sky130_fd_sc_hd__buf_2 hold1545 (.A(net2270),
    .X(net2826));
 sky130_fd_sc_hd__buf_2 hold1546 (.A(net1289),
    .X(net2827));
 sky130_fd_sc_hd__buf_2 hold1547 (.A(net2271),
    .X(net2828));
 sky130_fd_sc_hd__buf_2 hold1548 (.A(net3700),
    .X(net2829));
 sky130_fd_sc_hd__buf_2 hold1549 (.A(net3702),
    .X(net2830));
 sky130_fd_sc_hd__buf_2 hold155 (.A(net1450),
    .X(net1436));
 sky130_fd_sc_hd__buf_2 hold1550 (.A(net3704),
    .X(net2831));
 sky130_fd_sc_hd__buf_2 hold1551 (.A(net3706),
    .X(net2832));
 sky130_fd_sc_hd__buf_2 hold1552 (.A(net3708),
    .X(net2833));
 sky130_fd_sc_hd__buf_2 hold1553 (.A(net2280),
    .X(net2834));
 sky130_fd_sc_hd__buf_2 hold1554 (.A(net1297),
    .X(net2835));
 sky130_fd_sc_hd__buf_2 hold1555 (.A(net2281),
    .X(net2836));
 sky130_fd_sc_hd__buf_2 hold1556 (.A(_1086_),
    .X(net2837));
 sky130_fd_sc_hd__buf_2 hold1557 (.A(net2282),
    .X(net2838));
 sky130_fd_sc_hd__buf_2 hold1558 (.A(net1298),
    .X(net2839));
 sky130_fd_sc_hd__buf_2 hold1559 (.A(net2283),
    .X(net2840));
 sky130_fd_sc_hd__buf_2 hold156 (.A(net1452),
    .X(net1437));
 sky130_fd_sc_hd__buf_2 hold1560 (.A(net3690),
    .X(net2841));
 sky130_fd_sc_hd__buf_2 hold1561 (.A(net3692),
    .X(net2842));
 sky130_fd_sc_hd__buf_2 hold1562 (.A(net3694),
    .X(net2843));
 sky130_fd_sc_hd__buf_2 hold1563 (.A(net3696),
    .X(net2844));
 sky130_fd_sc_hd__buf_2 hold1564 (.A(net3698),
    .X(net2845));
 sky130_fd_sc_hd__buf_2 hold1565 (.A(net2286),
    .X(net2846));
 sky130_fd_sc_hd__buf_2 hold1566 (.A(net1303),
    .X(net2847));
 sky130_fd_sc_hd__buf_2 hold1567 (.A(net2287),
    .X(net2848));
 sky130_fd_sc_hd__buf_2 hold1568 (.A(_1077_),
    .X(net2849));
 sky130_fd_sc_hd__buf_2 hold1569 (.A(net2288),
    .X(net2850));
 sky130_fd_sc_hd__buf_2 hold157 (.A(net1454),
    .X(net1438));
 sky130_fd_sc_hd__buf_2 hold1570 (.A(net1304),
    .X(net2851));
 sky130_fd_sc_hd__buf_2 hold1571 (.A(net2289),
    .X(net2852));
 sky130_fd_sc_hd__buf_2 hold1572 (.A(net3710),
    .X(net2853));
 sky130_fd_sc_hd__buf_2 hold1573 (.A(net3712),
    .X(net2854));
 sky130_fd_sc_hd__buf_2 hold1574 (.A(net3714),
    .X(net2855));
 sky130_fd_sc_hd__buf_2 hold1575 (.A(net3716),
    .X(net2856));
 sky130_fd_sc_hd__buf_2 hold1576 (.A(net3718),
    .X(net2857));
 sky130_fd_sc_hd__buf_2 hold1577 (.A(net2292),
    .X(net2858));
 sky130_fd_sc_hd__buf_2 hold1578 (.A(net1321),
    .X(net2859));
 sky130_fd_sc_hd__buf_2 hold1579 (.A(net2293),
    .X(net2860));
 sky130_fd_sc_hd__buf_2 hold158 (.A(net1456),
    .X(net1439));
 sky130_fd_sc_hd__buf_2 hold1580 (.A(_1078_),
    .X(net2861));
 sky130_fd_sc_hd__buf_2 hold1581 (.A(net2294),
    .X(net2862));
 sky130_fd_sc_hd__buf_2 hold1582 (.A(net1322),
    .X(net2863));
 sky130_fd_sc_hd__buf_2 hold1583 (.A(net2295),
    .X(net2864));
 sky130_fd_sc_hd__buf_2 hold1584 (.A(net3720),
    .X(net2865));
 sky130_fd_sc_hd__buf_2 hold1585 (.A(net3722),
    .X(net2866));
 sky130_fd_sc_hd__buf_2 hold1586 (.A(net3724),
    .X(net2867));
 sky130_fd_sc_hd__buf_2 hold1587 (.A(net3726),
    .X(net2868));
 sky130_fd_sc_hd__buf_2 hold1588 (.A(net3728),
    .X(net2869));
 sky130_fd_sc_hd__buf_2 hold1589 (.A(net2304),
    .X(net2870));
 sky130_fd_sc_hd__buf_2 hold159 (.A(net1458),
    .X(net1440));
 sky130_fd_sc_hd__buf_2 hold1590 (.A(net1327),
    .X(net2871));
 sky130_fd_sc_hd__buf_2 hold1591 (.A(net2305),
    .X(net2872));
 sky130_fd_sc_hd__buf_2 hold1592 (.A(_1087_),
    .X(net2873));
 sky130_fd_sc_hd__buf_2 hold1593 (.A(net2306),
    .X(net2874));
 sky130_fd_sc_hd__buf_2 hold1594 (.A(net1328),
    .X(net2875));
 sky130_fd_sc_hd__buf_2 hold1595 (.A(net2307),
    .X(net2876));
 sky130_fd_sc_hd__buf_2 hold1596 (.A(net3738),
    .X(net2877));
 sky130_fd_sc_hd__buf_2 hold1597 (.A(net3740),
    .X(net2878));
 sky130_fd_sc_hd__buf_2 hold1598 (.A(net3742),
    .X(net2879));
 sky130_fd_sc_hd__buf_2 hold1599 (.A(net3744),
    .X(net2880));
 sky130_fd_sc_hd__buf_2 hold16 (.A(net2834),
    .X(net1297));
 sky130_fd_sc_hd__buf_2 hold160 (.A(_2126_),
    .X(net1441));
 sky130_fd_sc_hd__buf_2 hold1600 (.A(net3746),
    .X(net2881));
 sky130_fd_sc_hd__buf_2 hold1601 (.A(net2298),
    .X(net2882));
 sky130_fd_sc_hd__buf_2 hold1602 (.A(net1324),
    .X(net2883));
 sky130_fd_sc_hd__buf_2 hold1603 (.A(net2299),
    .X(net2884));
 sky130_fd_sc_hd__buf_2 hold1604 (.A(_1089_),
    .X(net2885));
 sky130_fd_sc_hd__buf_2 hold1605 (.A(net2300),
    .X(net2886));
 sky130_fd_sc_hd__buf_2 hold1606 (.A(net1325),
    .X(net2887));
 sky130_fd_sc_hd__buf_2 hold1607 (.A(net2301),
    .X(net2888));
 sky130_fd_sc_hd__buf_2 hold1608 (.A(net3729),
    .X(net2889));
 sky130_fd_sc_hd__buf_2 hold1609 (.A(net3731),
    .X(net2890));
 sky130_fd_sc_hd__buf_2 hold161 (.A(net1427),
    .X(net1442));
 sky130_fd_sc_hd__buf_2 hold1610 (.A(net3733),
    .X(net2891));
 sky130_fd_sc_hd__buf_2 hold1611 (.A(net3735),
    .X(net2892));
 sky130_fd_sc_hd__buf_2 hold1612 (.A(net3737),
    .X(net2893));
 sky130_fd_sc_hd__buf_2 hold1613 (.A(net2310),
    .X(net2894));
 sky130_fd_sc_hd__buf_2 hold1614 (.A(net1330),
    .X(net2895));
 sky130_fd_sc_hd__buf_2 hold1615 (.A(net2311),
    .X(net2896));
 sky130_fd_sc_hd__buf_2 hold1616 (.A(_1088_),
    .X(net2897));
 sky130_fd_sc_hd__buf_2 hold1617 (.A(net2312),
    .X(net2898));
 sky130_fd_sc_hd__buf_2 hold1618 (.A(net1331),
    .X(net2899));
 sky130_fd_sc_hd__buf_2 hold1619 (.A(net2313),
    .X(net2900));
 sky130_fd_sc_hd__buf_2 hold162 (.A(_1234_),
    .X(net1443));
 sky130_fd_sc_hd__buf_2 hold1621 (.A(net4078),
    .X(net2902));
 sky130_fd_sc_hd__buf_2 hold1622 (.A(net4082),
    .X(net2903));
 sky130_fd_sc_hd__buf_2 hold1623 (.A(net3467),
    .X(net2904));
 sky130_fd_sc_hd__buf_2 hold1624 (.A(net3469),
    .X(net2905));
 sky130_fd_sc_hd__buf_2 hold1628 (.A(net4107),
    .X(net2909));
 sky130_fd_sc_hd__buf_2 hold1629 (.A(net3485),
    .X(net2910));
 sky130_fd_sc_hd__buf_2 hold163 (.A(wbs_sel_i[1]),
    .X(net1444));
 sky130_fd_sc_hd__buf_2 hold1630 (.A(net3487),
    .X(net2911));
 sky130_fd_sc_hd__buf_2 hold1631 (.A(net3489),
    .X(net2912));
 sky130_fd_sc_hd__buf_2 hold1639 (.A(net4085),
    .X(net2920));
 sky130_fd_sc_hd__buf_2 hold164 (.A(net1433),
    .X(net1445));
 sky130_fd_sc_hd__buf_2 hold1640 (.A(net3474),
    .X(net2921));
 sky130_fd_sc_hd__buf_2 hold1641 (.A(net3476),
    .X(net2922));
 sky130_fd_sc_hd__buf_2 hold1642 (.A(net3478),
    .X(net2923));
 sky130_fd_sc_hd__buf_2 hold1643 (.A(net2317),
    .X(net2924));
 sky130_fd_sc_hd__buf_2 hold1644 (.A(net3871),
    .X(net2925));
 sky130_fd_sc_hd__buf_2 hold1645 (.A(net3873),
    .X(net2926));
 sky130_fd_sc_hd__buf_2 hold1646 (.A(net3875),
    .X(net2927));
 sky130_fd_sc_hd__buf_2 hold1647 (.A(net3877),
    .X(net2928));
 sky130_fd_sc_hd__buf_2 hold1648 (.A(_0952_),
    .X(net2929));
 sky130_fd_sc_hd__buf_2 hold1649 (.A(net2320),
    .X(net2930));
 sky130_fd_sc_hd__buf_2 hold165 (.A(net1423),
    .X(net1446));
 sky130_fd_sc_hd__buf_2 hold1650 (.A(net1487),
    .X(net2931));
 sky130_fd_sc_hd__buf_2 hold1651 (.A(net2321),
    .X(net2932));
 sky130_fd_sc_hd__buf_2 hold1657 (.A(net3584),
    .X(net2938));
 sky130_fd_sc_hd__buf_2 hold1658 (.A(net3586),
    .X(net2939));
 sky130_fd_sc_hd__buf_2 hold1659 (.A(net3588),
    .X(net2940));
 sky130_fd_sc_hd__buf_2 hold166 (.A(net1434),
    .X(net1447));
 sky130_fd_sc_hd__buf_2 hold1660 (.A(net3590),
    .X(net2941));
 sky130_fd_sc_hd__buf_2 hold1666 (.A(net3597),
    .X(net2947));
 sky130_fd_sc_hd__buf_2 hold1667 (.A(net3599),
    .X(net2948));
 sky130_fd_sc_hd__buf_2 hold1668 (.A(net3601),
    .X(net2949));
 sky130_fd_sc_hd__buf_2 hold1669 (.A(net3603),
    .X(net2950));
 sky130_fd_sc_hd__buf_2 hold167 (.A(net1314),
    .X(net1448));
 sky130_fd_sc_hd__buf_2 hold1675 (.A(net3633),
    .X(net2956));
 sky130_fd_sc_hd__buf_2 hold1676 (.A(net3635),
    .X(net2957));
 sky130_fd_sc_hd__buf_2 hold1677 (.A(net3637),
    .X(net2958));
 sky130_fd_sc_hd__buf_2 hold1678 (.A(net3639),
    .X(net2959));
 sky130_fd_sc_hd__buf_2 hold168 (.A(net1435),
    .X(net1449));
 sky130_fd_sc_hd__buf_2 hold1683 (.A(net4101),
    .X(net2964));
 sky130_fd_sc_hd__buf_2 hold1684 (.A(net3497),
    .X(net2965));
 sky130_fd_sc_hd__buf_2 hold1685 (.A(net3499),
    .X(net2966));
 sky130_fd_sc_hd__buf_2 hold1686 (.A(net3501),
    .X(net2967));
 sky130_fd_sc_hd__buf_2 hold169 (.A(net1424),
    .X(net1450));
 sky130_fd_sc_hd__buf_2 hold1692 (.A(net3620),
    .X(net2973));
 sky130_fd_sc_hd__buf_2 hold1693 (.A(net3622),
    .X(net2974));
 sky130_fd_sc_hd__buf_2 hold1694 (.A(net3624),
    .X(net2975));
 sky130_fd_sc_hd__buf_2 hold1695 (.A(net3626),
    .X(net2976));
 sky130_fd_sc_hd__buf_2 hold17 (.A(net2838),
    .X(net1298));
 sky130_fd_sc_hd__buf_2 hold170 (.A(net1436),
    .X(net1451));
 sky130_fd_sc_hd__buf_2 hold1701 (.A(net3646),
    .X(net2982));
 sky130_fd_sc_hd__buf_2 hold1702 (.A(net3648),
    .X(net2983));
 sky130_fd_sc_hd__buf_2 hold1703 (.A(net3650),
    .X(net2984));
 sky130_fd_sc_hd__buf_2 hold1704 (.A(net3652),
    .X(net2985));
 sky130_fd_sc_hd__buf_2 hold1709 (.A(net4094),
    .X(net2990));
 sky130_fd_sc_hd__buf_2 hold171 (.A(net201),
    .X(net1452));
 sky130_fd_sc_hd__buf_2 hold1710 (.A(net3509),
    .X(net2991));
 sky130_fd_sc_hd__buf_2 hold1711 (.A(net3511),
    .X(net2992));
 sky130_fd_sc_hd__buf_2 hold1712 (.A(net3513),
    .X(net2993));
 sky130_fd_sc_hd__buf_2 hold1718 (.A(net3659),
    .X(net2999));
 sky130_fd_sc_hd__buf_2 hold1719 (.A(net3661),
    .X(net3000));
 sky130_fd_sc_hd__buf_2 hold172 (.A(net1437),
    .X(net1453));
 sky130_fd_sc_hd__buf_2 hold1720 (.A(net3663),
    .X(net3001));
 sky130_fd_sc_hd__buf_2 hold1721 (.A(net3665),
    .X(net3002));
 sky130_fd_sc_hd__buf_2 hold1727 (.A(net3682),
    .X(net3008));
 sky130_fd_sc_hd__buf_2 hold1728 (.A(net3684),
    .X(net3009));
 sky130_fd_sc_hd__buf_2 hold1729 (.A(net3686),
    .X(net3010));
 sky130_fd_sc_hd__buf_2 hold173 (.A(net1425),
    .X(net1454));
 sky130_fd_sc_hd__buf_2 hold1730 (.A(net3688),
    .X(net3011));
 sky130_fd_sc_hd__buf_2 hold1735 (.A(net4113),
    .X(net3016));
 sky130_fd_sc_hd__buf_2 hold1736 (.A(net3563),
    .X(net3017));
 sky130_fd_sc_hd__buf_2 hold1737 (.A(net3565),
    .X(net3018));
 sky130_fd_sc_hd__buf_2 hold1738 (.A(net3567),
    .X(net3019));
 sky130_fd_sc_hd__buf_2 hold174 (.A(net1438),
    .X(net1455));
 sky130_fd_sc_hd__buf_2 hold1744 (.A(net3830),
    .X(net3025));
 sky130_fd_sc_hd__buf_2 hold1745 (.A(net3832),
    .X(net3026));
 sky130_fd_sc_hd__buf_2 hold1746 (.A(net3834),
    .X(net3027));
 sky130_fd_sc_hd__buf_2 hold1747 (.A(net3836),
    .X(net3028));
 sky130_fd_sc_hd__buf_2 hold175 (.A(net1315),
    .X(net1456));
 sky130_fd_sc_hd__buf_2 hold1753 (.A(net3843),
    .X(net3034));
 sky130_fd_sc_hd__buf_2 hold1754 (.A(net3845),
    .X(net3035));
 sky130_fd_sc_hd__buf_2 hold1755 (.A(net3847),
    .X(net3036));
 sky130_fd_sc_hd__buf_2 hold1756 (.A(net3849),
    .X(net3037));
 sky130_fd_sc_hd__buf_2 hold176 (.A(net1439),
    .X(net1457));
 sky130_fd_sc_hd__buf_2 hold1762 (.A(net3752),
    .X(net3043));
 sky130_fd_sc_hd__buf_2 hold1763 (.A(net3754),
    .X(net3044));
 sky130_fd_sc_hd__buf_2 hold1764 (.A(net3756),
    .X(net3045));
 sky130_fd_sc_hd__buf_2 hold1765 (.A(net3758),
    .X(net3046));
 sky130_fd_sc_hd__buf_2 hold177 (.A(net1426),
    .X(net1458));
 sky130_fd_sc_hd__buf_2 hold1771 (.A(net3765),
    .X(net3052));
 sky130_fd_sc_hd__buf_2 hold1772 (.A(net3767),
    .X(net3053));
 sky130_fd_sc_hd__buf_2 hold1773 (.A(net3769),
    .X(net3054));
 sky130_fd_sc_hd__buf_2 hold1774 (.A(net3771),
    .X(net3055));
 sky130_fd_sc_hd__buf_2 hold178 (.A(net3327),
    .X(net1459));
 sky130_fd_sc_hd__buf_2 hold1780 (.A(net3778),
    .X(net3061));
 sky130_fd_sc_hd__buf_2 hold1781 (.A(net3780),
    .X(net3062));
 sky130_fd_sc_hd__buf_2 hold1782 (.A(net3782),
    .X(net3063));
 sky130_fd_sc_hd__buf_2 hold1783 (.A(net3784),
    .X(net3064));
 sky130_fd_sc_hd__buf_2 hold1789 (.A(net3804),
    .X(net3070));
 sky130_fd_sc_hd__buf_2 hold179 (.A(net1578),
    .X(net1460));
 sky130_fd_sc_hd__buf_2 hold1790 (.A(net3806),
    .X(net3071));
 sky130_fd_sc_hd__buf_2 hold1791 (.A(net3808),
    .X(net3072));
 sky130_fd_sc_hd__buf_2 hold1792 (.A(net3810),
    .X(net3073));
 sky130_fd_sc_hd__buf_2 hold1798 (.A(net3791),
    .X(net3079));
 sky130_fd_sc_hd__buf_2 hold1799 (.A(net3793),
    .X(net3080));
 sky130_fd_sc_hd__buf_2 hold18 (.A(net3529),
    .X(net1299));
 sky130_fd_sc_hd__buf_2 hold180 (.A(net3329),
    .X(net1461));
 sky130_fd_sc_hd__buf_2 hold1800 (.A(net3795),
    .X(net3081));
 sky130_fd_sc_hd__buf_2 hold1801 (.A(net3797),
    .X(net3082));
 sky130_fd_sc_hd__buf_2 hold1807 (.A(net3817),
    .X(net3088));
 sky130_fd_sc_hd__buf_2 hold1808 (.A(net3819),
    .X(net3089));
 sky130_fd_sc_hd__buf_2 hold1809 (.A(net3821),
    .X(net3090));
 sky130_fd_sc_hd__buf_2 hold181 (.A(net3243),
    .X(net1462));
 sky130_fd_sc_hd__buf_2 hold1810 (.A(net3823),
    .X(net3091));
 sky130_fd_sc_hd__buf_2 hold1813 (.A(net3853),
    .X(net3094));
 sky130_fd_sc_hd__buf_2 hold1814 (.A(net3855),
    .X(net3095));
 sky130_fd_sc_hd__buf_2 hold1815 (.A(net3857),
    .X(net3096));
 sky130_fd_sc_hd__buf_2 hold1816 (.A(net3859),
    .X(net3097));
 sky130_fd_sc_hd__buf_2 hold182 (.A(net3246),
    .X(net1463));
 sky130_fd_sc_hd__buf_2 hold1820 (.A(net4011),
    .X(net3101));
 sky130_fd_sc_hd__buf_2 hold1821 (.A(net2443),
    .X(net3102));
 sky130_fd_sc_hd__buf_2 hold1822 (.A(net2008),
    .X(net3103));
 sky130_fd_sc_hd__buf_2 hold1823 (.A(net2444),
    .X(net3104));
 sky130_fd_sc_hd__buf_2 hold1824 (.A(_0933_),
    .X(net3105));
 sky130_fd_sc_hd__buf_2 hold1825 (.A(net2445),
    .X(net3106));
 sky130_fd_sc_hd__buf_2 hold1826 (.A(net2009),
    .X(net3107));
 sky130_fd_sc_hd__buf_2 hold1827 (.A(net2446),
    .X(net3108));
 sky130_fd_sc_hd__buf_2 hold183 (.A(net639),
    .X(net1464));
 sky130_fd_sc_hd__buf_2 hold1830 (.A(net4020),
    .X(net3111));
 sky130_fd_sc_hd__buf_2 hold1831 (.A(net2353),
    .X(net3112));
 sky130_fd_sc_hd__buf_2 hold1832 (.A(_2040_),
    .X(net3113));
 sky130_fd_sc_hd__buf_2 hold1833 (.A(net2354),
    .X(net3114));
 sky130_fd_sc_hd__buf_2 hold1834 (.A(net1473),
    .X(net3115));
 sky130_fd_sc_hd__buf_2 hold1835 (.A(net2355),
    .X(net3116));
 sky130_fd_sc_hd__buf_2 hold1836 (.A(_1011_),
    .X(net3117));
 sky130_fd_sc_hd__buf_2 hold1837 (.A(net2332),
    .X(net3118));
 sky130_fd_sc_hd__buf_2 hold1838 (.A(net1432),
    .X(net3119));
 sky130_fd_sc_hd__buf_2 hold1839 (.A(net2333),
    .X(net3120));
 sky130_fd_sc_hd__buf_2 hold184 (.A(net4164),
    .X(net1465));
 sky130_fd_sc_hd__buf_2 hold1843 (.A(net4016),
    .X(net3124));
 sky130_fd_sc_hd__buf_2 hold1844 (.A(net2450),
    .X(net3125));
 sky130_fd_sc_hd__buf_2 hold1845 (.A(net2067),
    .X(net3126));
 sky130_fd_sc_hd__buf_2 hold1846 (.A(net2451),
    .X(net3127));
 sky130_fd_sc_hd__buf_2 hold1847 (.A(_0936_),
    .X(net3128));
 sky130_fd_sc_hd__buf_2 hold1848 (.A(net2452),
    .X(net3129));
 sky130_fd_sc_hd__buf_2 hold1849 (.A(net2068),
    .X(net3130));
 sky130_fd_sc_hd__buf_2 hold185 (.A(net1417),
    .X(net1466));
 sky130_fd_sc_hd__buf_2 hold1850 (.A(net2453),
    .X(net3131));
 sky130_fd_sc_hd__buf_2 hold1854 (.A(net3864),
    .X(net3135));
 sky130_fd_sc_hd__buf_2 hold1855 (.A(net3866),
    .X(net3136));
 sky130_fd_sc_hd__buf_2 hold1856 (.A(net3868),
    .X(net3137));
 sky130_fd_sc_hd__buf_2 hold1857 (.A(net2580),
    .X(net3138));
 sky130_fd_sc_hd__buf_2 hold1858 (.A(wbs_we_i),
    .X(net3139));
 sky130_fd_sc_hd__buf_2 hold1859 (.A(net2322),
    .X(net3140));
 sky130_fd_sc_hd__buf_2 hold186 (.A(net3475),
    .X(net1467));
 sky130_fd_sc_hd__buf_2 hold1860 (.A(net1475),
    .X(net3141));
 sky130_fd_sc_hd__buf_2 hold1861 (.A(net2323),
    .X(net3142));
 sky130_fd_sc_hd__buf_2 hold1862 (.A(net1429),
    .X(net3143));
 sky130_fd_sc_hd__buf_2 hold1863 (.A(net2324),
    .X(net3144));
 sky130_fd_sc_hd__buf_2 hold1864 (.A(_1012_),
    .X(net3145));
 sky130_fd_sc_hd__buf_2 hold1865 (.A(net2356),
    .X(net3146));
 sky130_fd_sc_hd__buf_2 hold1866 (.A(net1474),
    .X(net3147));
 sky130_fd_sc_hd__buf_2 hold1867 (.A(net2357),
    .X(net3148));
 sky130_fd_sc_hd__buf_2 hold187 (.A(net3325),
    .X(net1468));
 sky130_fd_sc_hd__buf_2 hold1871 (.A(net4025),
    .X(net3152));
 sky130_fd_sc_hd__buf_2 hold1872 (.A(net2457),
    .X(net3153));
 sky130_fd_sc_hd__buf_2 hold1873 (.A(net1865),
    .X(net3154));
 sky130_fd_sc_hd__buf_2 hold1874 (.A(net2458),
    .X(net3155));
 sky130_fd_sc_hd__buf_2 hold1875 (.A(_0937_),
    .X(net3156));
 sky130_fd_sc_hd__buf_2 hold1876 (.A(net2459),
    .X(net3157));
 sky130_fd_sc_hd__buf_2 hold1877 (.A(net1866),
    .X(net3158));
 sky130_fd_sc_hd__buf_2 hold1878 (.A(net2460),
    .X(net3159));
 sky130_fd_sc_hd__buf_2 hold188 (.A(net1575),
    .X(net1469));
 sky130_fd_sc_hd__buf_2 hold1882 (.A(net4029),
    .X(net3163));
 sky130_fd_sc_hd__buf_2 hold1883 (.A(net2499),
    .X(net3164));
 sky130_fd_sc_hd__buf_2 hold1884 (.A(net2148),
    .X(net3165));
 sky130_fd_sc_hd__buf_2 hold1885 (.A(net2500),
    .X(net3166));
 sky130_fd_sc_hd__buf_2 hold1886 (.A(_0943_),
    .X(net3167));
 sky130_fd_sc_hd__buf_2 hold1887 (.A(net2501),
    .X(net3168));
 sky130_fd_sc_hd__buf_2 hold1888 (.A(net2149),
    .X(net3169));
 sky130_fd_sc_hd__buf_2 hold1889 (.A(net2502),
    .X(net3170));
 sky130_fd_sc_hd__buf_2 hold189 (.A(net1577),
    .X(net1470));
 sky130_fd_sc_hd__buf_2 hold1893 (.A(net4033),
    .X(net3174));
 sky130_fd_sc_hd__buf_2 hold1894 (.A(net2485),
    .X(net3175));
 sky130_fd_sc_hd__buf_2 hold1895 (.A(net2122),
    .X(net3176));
 sky130_fd_sc_hd__buf_2 hold1896 (.A(net2486),
    .X(net3177));
 sky130_fd_sc_hd__buf_2 hold1897 (.A(_0940_),
    .X(net3178));
 sky130_fd_sc_hd__buf_2 hold1898 (.A(net2487),
    .X(net3179));
 sky130_fd_sc_hd__buf_2 hold1899 (.A(net2123),
    .X(net3180));
 sky130_fd_sc_hd__buf_2 hold19 (.A(net2762),
    .X(net1300));
 sky130_fd_sc_hd__buf_2 hold190 (.A(net1579),
    .X(net1471));
 sky130_fd_sc_hd__buf_2 hold1900 (.A(net2488),
    .X(net3181));
 sky130_fd_sc_hd__buf_2 hold1904 (.A(net4037),
    .X(net3185));
 sky130_fd_sc_hd__buf_2 hold1905 (.A(net2478),
    .X(net3186));
 sky130_fd_sc_hd__buf_2 hold1906 (.A(net2138),
    .X(net3187));
 sky130_fd_sc_hd__buf_2 hold1907 (.A(net2479),
    .X(net3188));
 sky130_fd_sc_hd__buf_2 hold1908 (.A(_0942_),
    .X(net3189));
 sky130_fd_sc_hd__buf_2 hold1909 (.A(net2480),
    .X(net3190));
 sky130_fd_sc_hd__buf_2 hold191 (.A(_2039_),
    .X(net1472));
 sky130_fd_sc_hd__buf_2 hold1910 (.A(net2139),
    .X(net3191));
 sky130_fd_sc_hd__buf_2 hold1911 (.A(net2481),
    .X(net3192));
 sky130_fd_sc_hd__buf_2 hold1915 (.A(net4041),
    .X(net3196));
 sky130_fd_sc_hd__buf_2 hold1916 (.A(net2492),
    .X(net3197));
 sky130_fd_sc_hd__buf_2 hold1917 (.A(net2133),
    .X(net3198));
 sky130_fd_sc_hd__buf_2 hold1918 (.A(net2493),
    .X(net3199));
 sky130_fd_sc_hd__buf_2 hold1919 (.A(_0939_),
    .X(net3200));
 sky130_fd_sc_hd__buf_2 hold192 (.A(net3114),
    .X(net1473));
 sky130_fd_sc_hd__buf_2 hold1920 (.A(net2494),
    .X(net3201));
 sky130_fd_sc_hd__buf_2 hold1921 (.A(net2134),
    .X(net3202));
 sky130_fd_sc_hd__buf_2 hold1922 (.A(net2495),
    .X(net3203));
 sky130_fd_sc_hd__buf_2 hold1926 (.A(net4049),
    .X(net3207));
 sky130_fd_sc_hd__buf_2 hold1927 (.A(net2506),
    .X(net3208));
 sky130_fd_sc_hd__buf_2 hold1928 (.A(net1870),
    .X(net3209));
 sky130_fd_sc_hd__buf_2 hold1929 (.A(net2507),
    .X(net3210));
 sky130_fd_sc_hd__buf_2 hold193 (.A(net3146),
    .X(net1474));
 sky130_fd_sc_hd__buf_2 hold1930 (.A(_0935_),
    .X(net3211));
 sky130_fd_sc_hd__buf_2 hold1931 (.A(net2508),
    .X(net3212));
 sky130_fd_sc_hd__buf_2 hold1932 (.A(net1871),
    .X(net3213));
 sky130_fd_sc_hd__buf_2 hold1933 (.A(net2509),
    .X(net3214));
 sky130_fd_sc_hd__buf_2 hold1937 (.A(net4053),
    .X(net3218));
 sky130_fd_sc_hd__buf_2 hold1938 (.A(net2513),
    .X(net3219));
 sky130_fd_sc_hd__buf_2 hold1939 (.A(net2143),
    .X(net3220));
 sky130_fd_sc_hd__buf_2 hold194 (.A(net3140),
    .X(net1475));
 sky130_fd_sc_hd__buf_2 hold1940 (.A(net2514),
    .X(net3221));
 sky130_fd_sc_hd__buf_2 hold1941 (.A(_0938_),
    .X(net3222));
 sky130_fd_sc_hd__buf_2 hold1942 (.A(net2515),
    .X(net3223));
 sky130_fd_sc_hd__buf_2 hold1943 (.A(net2144),
    .X(net3224));
 sky130_fd_sc_hd__buf_2 hold1944 (.A(net2516),
    .X(net3225));
 sky130_fd_sc_hd__buf_2 hold1948 (.A(net4045),
    .X(net3229));
 sky130_fd_sc_hd__buf_2 hold1949 (.A(net2520),
    .X(net3230));
 sky130_fd_sc_hd__buf_2 hold195 (.A(net3144),
    .X(net1476));
 sky130_fd_sc_hd__buf_2 hold1950 (.A(net2084),
    .X(net3231));
 sky130_fd_sc_hd__buf_2 hold1951 (.A(net2521),
    .X(net3232));
 sky130_fd_sc_hd__buf_2 hold1952 (.A(_0934_),
    .X(net3233));
 sky130_fd_sc_hd__buf_2 hold1953 (.A(net2522),
    .X(net3234));
 sky130_fd_sc_hd__buf_2 hold1954 (.A(net2085),
    .X(net3235));
 sky130_fd_sc_hd__buf_2 hold1955 (.A(net2523),
    .X(net3236));
 sky130_fd_sc_hd__buf_2 hold196 (.A(net2326),
    .X(net1477));
 sky130_fd_sc_hd__buf_2 hold1960 (.A(net3328),
    .X(net3241));
 sky130_fd_sc_hd__buf_2 hold1961 (.A(net3330),
    .X(net3242));
 sky130_fd_sc_hd__buf_2 hold1962 (.A(_2124_),
    .X(net3243));
 sky130_fd_sc_hd__buf_2 hold1963 (.A(net1462),
    .X(net3244));
 sky130_fd_sc_hd__buf_2 hold1964 (.A(_1099_),
    .X(net3245));
 sky130_fd_sc_hd__buf_2 hold1965 (.A(net2341),
    .X(net3246));
 sky130_fd_sc_hd__buf_2 hold1966 (.A(net1463),
    .X(net3247));
 sky130_fd_sc_hd__buf_2 hold1967 (.A(net2342),
    .X(net3248));
 sky130_fd_sc_hd__buf_2 hold197 (.A(net2328),
    .X(net1478));
 sky130_fd_sc_hd__buf_2 hold1975 (.A(net3885),
    .X(net3256));
 sky130_fd_sc_hd__buf_2 hold1976 (.A(net3887),
    .X(net3257));
 sky130_fd_sc_hd__buf_2 hold1977 (.A(net3889),
    .X(net3258));
 sky130_fd_sc_hd__buf_2 hold1978 (.A(net2596),
    .X(net3259));
 sky130_fd_sc_hd__buf_2 hold198 (.A(net2401),
    .X(net1479));
 sky130_fd_sc_hd__buf_2 hold1986 (.A(net3898),
    .X(net3267));
 sky130_fd_sc_hd__buf_2 hold1987 (.A(net3900),
    .X(net3268));
 sky130_fd_sc_hd__buf_2 hold1988 (.A(net3902),
    .X(net3269));
 sky130_fd_sc_hd__buf_2 hold1989 (.A(net2605),
    .X(net3270));
 sky130_fd_sc_hd__buf_2 hold199 (.A(net2404),
    .X(net1480));
 sky130_fd_sc_hd__buf_2 hold1992 (.A(net3906),
    .X(net3273));
 sky130_fd_sc_hd__buf_2 hold1993 (.A(net3908),
    .X(net3274));
 sky130_fd_sc_hd__buf_2 hold1994 (.A(net3910),
    .X(net3275));
 sky130_fd_sc_hd__buf_2 hold1995 (.A(net2587),
    .X(net3276));
 sky130_fd_sc_hd__buf_2 hold1998 (.A(net3914),
    .X(net3279));
 sky130_fd_sc_hd__buf_2 hold1999 (.A(net3916),
    .X(net3280));
 sky130_fd_sc_hd__buf_2 hold20 (.A(net2766),
    .X(net1301));
 sky130_fd_sc_hd__buf_2 hold200 (.A(net3332),
    .X(net1481));
 sky130_fd_sc_hd__buf_2 hold2000 (.A(net3918),
    .X(net3281));
 sky130_fd_sc_hd__buf_2 hold2001 (.A(net2609),
    .X(net3282));
 sky130_fd_sc_hd__buf_2 hold2004 (.A(net3922),
    .X(net3285));
 sky130_fd_sc_hd__buf_2 hold2005 (.A(net3924),
    .X(net3286));
 sky130_fd_sc_hd__buf_2 hold2006 (.A(net3926),
    .X(net3287));
 sky130_fd_sc_hd__buf_2 hold2007 (.A(net2613),
    .X(net3288));
 sky130_fd_sc_hd__buf_2 hold2010 (.A(net3943),
    .X(net3291));
 sky130_fd_sc_hd__buf_2 hold2011 (.A(net3945),
    .X(net3292));
 sky130_fd_sc_hd__buf_2 hold2012 (.A(net3947),
    .X(net3293));
 sky130_fd_sc_hd__buf_2 hold2013 (.A(net2617),
    .X(net3294));
 sky130_fd_sc_hd__buf_2 hold202 (.A(net647),
    .X(net1483));
 sky130_fd_sc_hd__buf_2 hold2021 (.A(net3935),
    .X(net3302));
 sky130_fd_sc_hd__buf_2 hold2022 (.A(net3937),
    .X(net3303));
 sky130_fd_sc_hd__buf_2 hold2023 (.A(net3939),
    .X(net3304));
 sky130_fd_sc_hd__buf_2 hold2024 (.A(net2634),
    .X(net3305));
 sky130_fd_sc_hd__buf_2 hold2027 (.A(net3951),
    .X(net3308));
 sky130_fd_sc_hd__buf_2 hold2028 (.A(net3953),
    .X(net3309));
 sky130_fd_sc_hd__buf_2 hold2029 (.A(net3955),
    .X(net3310));
 sky130_fd_sc_hd__buf_2 hold203 (.A(net3856),
    .X(net1484));
 sky130_fd_sc_hd__buf_2 hold2030 (.A(net2621),
    .X(net3311));
 sky130_fd_sc_hd__buf_2 hold2033 (.A(net3959),
    .X(net3314));
 sky130_fd_sc_hd__buf_2 hold2034 (.A(net3961),
    .X(net3315));
 sky130_fd_sc_hd__buf_2 hold2035 (.A(net3963),
    .X(net3316));
 sky130_fd_sc_hd__buf_2 hold2036 (.A(net2625),
    .X(net3317));
 sky130_fd_sc_hd__buf_2 hold2039 (.A(net3967),
    .X(net3320));
 sky130_fd_sc_hd__buf_2 hold204 (.A(net1464),
    .X(net1485));
 sky130_fd_sc_hd__buf_2 hold2040 (.A(net3969),
    .X(net3321));
 sky130_fd_sc_hd__buf_2 hold2041 (.A(net3971),
    .X(net3322));
 sky130_fd_sc_hd__buf_2 hold2042 (.A(net2638),
    .X(net3323));
 sky130_fd_sc_hd__buf_2 hold2043 (.A(wbs_stb_i),
    .X(net3324));
 sky130_fd_sc_hd__buf_2 hold2044 (.A(net1573),
    .X(net3325));
 sky130_fd_sc_hd__buf_2 hold2045 (.A(net1468),
    .X(net3326));
 sky130_fd_sc_hd__buf_2 hold2046 (.A(net1574),
    .X(net3327));
 sky130_fd_sc_hd__buf_2 hold2047 (.A(_2123_),
    .X(net3328));
 sky130_fd_sc_hd__buf_2 hold2048 (.A(net3241),
    .X(net3329));
 sky130_fd_sc_hd__buf_2 hold2049 (.A(net1461),
    .X(net3330));
 sky130_fd_sc_hd__buf_2 hold205 (.A(net3874),
    .X(net1486));
 sky130_fd_sc_hd__buf_2 hold2050 (.A(_1100_),
    .X(net3331));
 sky130_fd_sc_hd__buf_2 hold2051 (.A(net2406),
    .X(net3332));
 sky130_fd_sc_hd__buf_2 hold2052 (.A(net1481),
    .X(net3333));
 sky130_fd_sc_hd__buf_2 hold2053 (.A(net2407),
    .X(net3334));
 sky130_fd_sc_hd__buf_2 hold2056 (.A(net3975),
    .X(net3337));
 sky130_fd_sc_hd__buf_2 hold2057 (.A(net3977),
    .X(net3338));
 sky130_fd_sc_hd__buf_2 hold2058 (.A(net3979),
    .X(net3339));
 sky130_fd_sc_hd__buf_2 hold2059 (.A(net2642),
    .X(net3340));
 sky130_fd_sc_hd__buf_2 hold206 (.A(net2930),
    .X(net1487));
 sky130_fd_sc_hd__buf_2 hold2067 (.A(net3987),
    .X(net3348));
 sky130_fd_sc_hd__buf_2 hold2068 (.A(net3989),
    .X(net3349));
 sky130_fd_sc_hd__buf_2 hold2069 (.A(net2210),
    .X(net3350));
 sky130_fd_sc_hd__buf_2 hold2070 (.A(net2695),
    .X(net3351));
 sky130_fd_sc_hd__buf_2 hold2074 (.A(net3994),
    .X(net3355));
 sky130_fd_sc_hd__buf_2 hold2075 (.A(net2699),
    .X(net3356));
 sky130_fd_sc_hd__buf_2 hold2076 (.A(net1718),
    .X(net3357));
 sky130_fd_sc_hd__buf_2 hold2077 (.A(net2700),
    .X(net3358));
 sky130_fd_sc_hd__buf_2 hold2081 (.A(_0974_),
    .X(net3362));
 sky130_fd_sc_hd__buf_2 hold2082 (.A(net2704),
    .X(net3363));
 sky130_fd_sc_hd__buf_2 hold2083 (.A(net1726),
    .X(net3364));
 sky130_fd_sc_hd__buf_2 hold2084 (.A(net2705),
    .X(net3365));
 sky130_fd_sc_hd__buf_2 hold2088 (.A(_0977_),
    .X(net3369));
 sky130_fd_sc_hd__buf_2 hold2089 (.A(net2709),
    .X(net3370));
 sky130_fd_sc_hd__buf_2 hold209 (.A(net1682),
    .X(net1490));
 sky130_fd_sc_hd__buf_2 hold2090 (.A(net1722),
    .X(net3371));
 sky130_fd_sc_hd__buf_2 hold2091 (.A(net2710),
    .X(net3372));
 sky130_fd_sc_hd__buf_2 hold2095 (.A(_0976_),
    .X(net3376));
 sky130_fd_sc_hd__buf_2 hold2096 (.A(net2714),
    .X(net3377));
 sky130_fd_sc_hd__buf_2 hold2097 (.A(net1730),
    .X(net3378));
 sky130_fd_sc_hd__buf_2 hold2098 (.A(net2715),
    .X(net3379));
 sky130_fd_sc_hd__buf_2 hold21 (.A(net3693),
    .X(net1302));
 sky130_fd_sc_hd__buf_2 hold210 (.A(net1518),
    .X(net1491));
 sky130_fd_sc_hd__buf_2 hold2102 (.A(_0971_),
    .X(net3383));
 sky130_fd_sc_hd__buf_2 hold2103 (.A(net2719),
    .X(net3384));
 sky130_fd_sc_hd__buf_2 hold2104 (.A(net1744),
    .X(net3385));
 sky130_fd_sc_hd__buf_2 hold2105 (.A(net2720),
    .X(net3386));
 sky130_fd_sc_hd__buf_2 hold2109 (.A(_0972_),
    .X(net3390));
 sky130_fd_sc_hd__buf_2 hold211 (.A(net1507),
    .X(net1492));
 sky130_fd_sc_hd__buf_2 hold2110 (.A(net2724),
    .X(net3391));
 sky130_fd_sc_hd__buf_2 hold2111 (.A(net1755),
    .X(net3392));
 sky130_fd_sc_hd__buf_2 hold2112 (.A(net2725),
    .X(net3393));
 sky130_fd_sc_hd__buf_2 hold2116 (.A(_2079_),
    .X(net3397));
 sky130_fd_sc_hd__buf_2 hold2117 (.A(net2646),
    .X(net3398));
 sky130_fd_sc_hd__buf_2 hold2118 (.A(net1769),
    .X(net3399));
 sky130_fd_sc_hd__buf_2 hold2119 (.A(net2647),
    .X(net3400));
 sky130_fd_sc_hd__buf_2 hold212 (.A(net1511),
    .X(net1493));
 sky130_fd_sc_hd__buf_2 hold2120 (.A(_1056_),
    .X(net3401));
 sky130_fd_sc_hd__buf_2 hold2121 (.A(net2648),
    .X(net3402));
 sky130_fd_sc_hd__buf_2 hold2125 (.A(_2075_),
    .X(net3406));
 sky130_fd_sc_hd__buf_2 hold2126 (.A(net2653),
    .X(net3407));
 sky130_fd_sc_hd__buf_2 hold2127 (.A(net1774),
    .X(net3408));
 sky130_fd_sc_hd__buf_2 hold2128 (.A(net2654),
    .X(net3409));
 sky130_fd_sc_hd__buf_2 hold2129 (.A(_1055_),
    .X(net3410));
 sky130_fd_sc_hd__buf_2 hold213 (.A(_1248_),
    .X(net1494));
 sky130_fd_sc_hd__buf_2 hold2130 (.A(net2655),
    .X(net3411));
 sky130_fd_sc_hd__buf_2 hold2134 (.A(_2083_),
    .X(net3415));
 sky130_fd_sc_hd__buf_2 hold2135 (.A(net2660),
    .X(net3416));
 sky130_fd_sc_hd__buf_2 hold2136 (.A(net1802),
    .X(net3417));
 sky130_fd_sc_hd__buf_2 hold2137 (.A(net2661),
    .X(net3418));
 sky130_fd_sc_hd__buf_2 hold2138 (.A(_1057_),
    .X(net3419));
 sky130_fd_sc_hd__buf_2 hold2139 (.A(net2662),
    .X(net3420));
 sky130_fd_sc_hd__buf_2 hold214 (.A(net1516),
    .X(net1495));
 sky130_fd_sc_hd__buf_2 hold2143 (.A(_2091_),
    .X(net3424));
 sky130_fd_sc_hd__buf_2 hold2144 (.A(net2667),
    .X(net3425));
 sky130_fd_sc_hd__buf_2 hold2145 (.A(net1822),
    .X(net3426));
 sky130_fd_sc_hd__buf_2 hold2146 (.A(net2668),
    .X(net3427));
 sky130_fd_sc_hd__buf_2 hold2147 (.A(_1059_),
    .X(net3428));
 sky130_fd_sc_hd__buf_2 hold2148 (.A(net2669),
    .X(net3429));
 sky130_fd_sc_hd__buf_2 hold215 (.A(net1504),
    .X(net1496));
 sky130_fd_sc_hd__buf_2 hold2152 (.A(_2071_),
    .X(net3433));
 sky130_fd_sc_hd__buf_2 hold2153 (.A(net2674),
    .X(net3434));
 sky130_fd_sc_hd__buf_2 hold2154 (.A(net1841),
    .X(net3435));
 sky130_fd_sc_hd__buf_2 hold2155 (.A(net2675),
    .X(net3436));
 sky130_fd_sc_hd__buf_2 hold2156 (.A(_1054_),
    .X(net3437));
 sky130_fd_sc_hd__buf_2 hold2157 (.A(net2676),
    .X(net3438));
 sky130_fd_sc_hd__buf_2 hold216 (.A(net1506),
    .X(net1497));
 sky130_fd_sc_hd__buf_2 hold2163 (.A(net437),
    .X(net3444));
 sky130_fd_sc_hd__buf_2 hold2164 (.A(net2683),
    .X(net3445));
 sky130_fd_sc_hd__buf_2 hold2165 (.A(net2234),
    .X(net3446));
 sky130_fd_sc_hd__buf_2 hold2166 (.A(net2684),
    .X(net3447));
 sky130_fd_sc_hd__buf_2 hold2167 (.A(_0582_),
    .X(net3448));
 sky130_fd_sc_hd__buf_2 hold2168 (.A(net2685),
    .X(net3449));
 sky130_fd_sc_hd__buf_2 hold217 (.A(net1508),
    .X(net1498));
 sky130_fd_sc_hd__buf_2 hold2171 (.A(net4166),
    .X(net3452));
 sky130_fd_sc_hd__buf_2 hold2172 (.A(net4070),
    .X(net3453));
 sky130_fd_sc_hd__buf_2 hold2173 (.A(net4072),
    .X(net3454));
 sky130_fd_sc_hd__buf_2 hold2174 (.A(net4074),
    .X(net3455));
 sky130_fd_sc_hd__buf_2 hold218 (.A(net1510),
    .X(net1499));
 sky130_fd_sc_hd__buf_2 hold2182 (.A(net4077),
    .X(net3463));
 sky130_fd_sc_hd__buf_2 hold2183 (.A(net4079),
    .X(net3464));
 sky130_fd_sc_hd__buf_2 hold2184 (.A(net4081),
    .X(net3465));
 sky130_fd_sc_hd__buf_2 hold2185 (.A(net2903),
    .X(net3466));
 sky130_fd_sc_hd__buf_2 hold2186 (.A(net1342),
    .X(net3467));
 sky130_fd_sc_hd__buf_2 hold2187 (.A(net2904),
    .X(net3468));
 sky130_fd_sc_hd__buf_2 hold2188 (.A(net2350),
    .X(net3469));
 sky130_fd_sc_hd__buf_2 hold2189 (.A(net2905),
    .X(net3470));
 sky130_fd_sc_hd__buf_2 hold219 (.A(net1512),
    .X(net1500));
 sky130_fd_sc_hd__buf_2 hold2191 (.A(net4084),
    .X(net3472));
 sky130_fd_sc_hd__buf_2 hold2192 (.A(net4086),
    .X(net3473));
 sky130_fd_sc_hd__buf_2 hold2193 (.A(net4088),
    .X(net3474));
 sky130_fd_sc_hd__buf_2 hold2194 (.A(net2921),
    .X(net3475));
 sky130_fd_sc_hd__buf_2 hold2195 (.A(net1467),
    .X(net3476));
 sky130_fd_sc_hd__buf_2 hold2196 (.A(net2922),
    .X(net3477));
 sky130_fd_sc_hd__buf_2 hold2197 (.A(net2360),
    .X(net3478));
 sky130_fd_sc_hd__buf_2 hold2198 (.A(net2923),
    .X(net3479));
 sky130_fd_sc_hd__buf_2 hold22 (.A(net2846),
    .X(net1303));
 sky130_fd_sc_hd__buf_2 hold220 (.A(_1249_),
    .X(net1501));
 sky130_fd_sc_hd__buf_2 hold2202 (.A(net4106),
    .X(net3483));
 sky130_fd_sc_hd__buf_2 hold2203 (.A(net2909),
    .X(net3484));
 sky130_fd_sc_hd__buf_2 hold2204 (.A(net2346),
    .X(net3485));
 sky130_fd_sc_hd__buf_2 hold2205 (.A(net2910),
    .X(net3486));
 sky130_fd_sc_hd__buf_2 hold2206 (.A(net1977),
    .X(net3487));
 sky130_fd_sc_hd__buf_2 hold2207 (.A(net2911),
    .X(net3488));
 sky130_fd_sc_hd__buf_2 hold2208 (.A(net2347),
    .X(net3489));
 sky130_fd_sc_hd__buf_2 hold2209 (.A(net2912),
    .X(net3490));
 sky130_fd_sc_hd__buf_2 hold221 (.A(net1515),
    .X(net1502));
 sky130_fd_sc_hd__buf_2 hold2214 (.A(net4100),
    .X(net3495));
 sky130_fd_sc_hd__buf_2 hold2215 (.A(net4102),
    .X(net3496));
 sky130_fd_sc_hd__buf_2 hold2216 (.A(net2432),
    .X(net3497));
 sky130_fd_sc_hd__buf_2 hold2217 (.A(net2965),
    .X(net3498));
 sky130_fd_sc_hd__buf_2 hold2218 (.A(net1909),
    .X(net3499));
 sky130_fd_sc_hd__buf_2 hold2219 (.A(net2966),
    .X(net3500));
 sky130_fd_sc_hd__buf_2 hold222 (.A(net1517),
    .X(net1503));
 sky130_fd_sc_hd__buf_2 hold2220 (.A(net2433),
    .X(net3501));
 sky130_fd_sc_hd__buf_2 hold2221 (.A(net2967),
    .X(net3502));
 sky130_fd_sc_hd__buf_2 hold2226 (.A(net4093),
    .X(net3507));
 sky130_fd_sc_hd__buf_2 hold2227 (.A(net4095),
    .X(net3508));
 sky130_fd_sc_hd__buf_2 hold2228 (.A(net2438),
    .X(net3509));
 sky130_fd_sc_hd__buf_2 hold2229 (.A(net2991),
    .X(net3510));
 sky130_fd_sc_hd__buf_2 hold223 (.A(net1491),
    .X(net1504));
 sky130_fd_sc_hd__buf_2 hold2230 (.A(net1922),
    .X(net3511));
 sky130_fd_sc_hd__buf_2 hold2231 (.A(net2992),
    .X(net3512));
 sky130_fd_sc_hd__buf_2 hold2232 (.A(net2439),
    .X(net3513));
 sky130_fd_sc_hd__buf_2 hold2233 (.A(net2993),
    .X(net3514));
 sky130_fd_sc_hd__buf_2 hold2234 (.A(wbs_adr_i[4]),
    .X(net3515));
 sky130_fd_sc_hd__buf_2 hold2235 (.A(net2745),
    .X(net3516));
 sky130_fd_sc_hd__buf_2 hold2236 (.A(net2236),
    .X(net3517));
 sky130_fd_sc_hd__buf_2 hold2237 (.A(net2746),
    .X(net3518));
 sky130_fd_sc_hd__buf_2 hold2238 (.A(net1293),
    .X(net3519));
 sky130_fd_sc_hd__buf_2 hold2239 (.A(net2747),
    .X(net3520));
 sky130_fd_sc_hd__buf_2 hold224 (.A(net1496),
    .X(net1505));
 sky130_fd_sc_hd__buf_2 hold2240 (.A(net2237),
    .X(net3521));
 sky130_fd_sc_hd__buf_2 hold2241 (.A(net2748),
    .X(net3522));
 sky130_fd_sc_hd__buf_2 hold2242 (.A(net161),
    .X(net3523));
 sky130_fd_sc_hd__buf_2 hold2243 (.A(net2749),
    .X(net3524));
 sky130_fd_sc_hd__buf_2 hold2244 (.A(net2238),
    .X(net3525));
 sky130_fd_sc_hd__buf_2 hold2245 (.A(wbs_adr_i[5]),
    .X(net3526));
 sky130_fd_sc_hd__buf_2 hold2246 (.A(net2757),
    .X(net3527));
 sky130_fd_sc_hd__buf_2 hold2247 (.A(net2242),
    .X(net3528));
 sky130_fd_sc_hd__buf_2 hold2248 (.A(net2758),
    .X(net3529));
 sky130_fd_sc_hd__buf_2 hold2249 (.A(net1299),
    .X(net3530));
 sky130_fd_sc_hd__buf_2 hold225 (.A(net203),
    .X(net1506));
 sky130_fd_sc_hd__buf_2 hold2250 (.A(net2759),
    .X(net3531));
 sky130_fd_sc_hd__buf_2 hold2251 (.A(net2243),
    .X(net3532));
 sky130_fd_sc_hd__buf_2 hold2252 (.A(net2760),
    .X(net3533));
 sky130_fd_sc_hd__buf_2 hold2253 (.A(net162),
    .X(net3534));
 sky130_fd_sc_hd__buf_2 hold2254 (.A(net2761),
    .X(net3535));
 sky130_fd_sc_hd__buf_2 hold2255 (.A(net2244),
    .X(net3536));
 sky130_fd_sc_hd__buf_2 hold2256 (.A(wbs_adr_i[6]),
    .X(net3537));
 sky130_fd_sc_hd__buf_2 hold2257 (.A(net2769),
    .X(net3538));
 sky130_fd_sc_hd__buf_2 hold2258 (.A(net2248),
    .X(net3539));
 sky130_fd_sc_hd__buf_2 hold2259 (.A(net2770),
    .X(net3540));
 sky130_fd_sc_hd__buf_2 hold226 (.A(net1497),
    .X(net1507));
 sky130_fd_sc_hd__buf_2 hold2260 (.A(net1305),
    .X(net3541));
 sky130_fd_sc_hd__buf_2 hold2261 (.A(net2771),
    .X(net3542));
 sky130_fd_sc_hd__buf_2 hold2262 (.A(net2249),
    .X(net3543));
 sky130_fd_sc_hd__buf_2 hold2263 (.A(net2772),
    .X(net3544));
 sky130_fd_sc_hd__buf_2 hold2264 (.A(net163),
    .X(net3545));
 sky130_fd_sc_hd__buf_2 hold2265 (.A(net2773),
    .X(net3546));
 sky130_fd_sc_hd__buf_2 hold2266 (.A(wbs_adr_i[7]),
    .X(net3547));
 sky130_fd_sc_hd__buf_2 hold2267 (.A(net2781),
    .X(net3548));
 sky130_fd_sc_hd__buf_2 hold2268 (.A(net2254),
    .X(net3549));
 sky130_fd_sc_hd__buf_2 hold2269 (.A(net2782),
    .X(net3550));
 sky130_fd_sc_hd__buf_2 hold227 (.A(net1492),
    .X(net1508));
 sky130_fd_sc_hd__buf_2 hold2270 (.A(net1311),
    .X(net3551));
 sky130_fd_sc_hd__buf_2 hold2271 (.A(net2783),
    .X(net3552));
 sky130_fd_sc_hd__buf_2 hold2272 (.A(net2255),
    .X(net3553));
 sky130_fd_sc_hd__buf_2 hold2273 (.A(net2784),
    .X(net3554));
 sky130_fd_sc_hd__buf_2 hold2274 (.A(net164),
    .X(net3555));
 sky130_fd_sc_hd__buf_2 hold2275 (.A(net2785),
    .X(net3556));
 sky130_fd_sc_hd__buf_2 hold228 (.A(net1498),
    .X(net1509));
 sky130_fd_sc_hd__buf_2 hold2280 (.A(net4112),
    .X(net3561));
 sky130_fd_sc_hd__buf_2 hold2281 (.A(net3016),
    .X(net3562));
 sky130_fd_sc_hd__buf_2 hold2282 (.A(net2528),
    .X(net3563));
 sky130_fd_sc_hd__buf_2 hold2283 (.A(net3017),
    .X(net3564));
 sky130_fd_sc_hd__buf_2 hold2284 (.A(net1943),
    .X(net3565));
 sky130_fd_sc_hd__buf_2 hold2285 (.A(net3018),
    .X(net3566));
 sky130_fd_sc_hd__buf_2 hold2286 (.A(net2529),
    .X(net3567));
 sky130_fd_sc_hd__buf_2 hold2287 (.A(net3019),
    .X(net3568));
 sky130_fd_sc_hd__buf_2 hold2288 (.A(wbs_adr_i[8]),
    .X(net3569));
 sky130_fd_sc_hd__buf_2 hold2289 (.A(net2793),
    .X(net3570));
 sky130_fd_sc_hd__buf_2 hold229 (.A(_2128_),
    .X(net1510));
 sky130_fd_sc_hd__buf_2 hold2290 (.A(net2260),
    .X(net3571));
 sky130_fd_sc_hd__buf_2 hold2291 (.A(net2794),
    .X(net3572));
 sky130_fd_sc_hd__buf_2 hold2292 (.A(net1308),
    .X(net3573));
 sky130_fd_sc_hd__buf_2 hold2293 (.A(net2795),
    .X(net3574));
 sky130_fd_sc_hd__buf_2 hold2294 (.A(net2261),
    .X(net3575));
 sky130_fd_sc_hd__buf_2 hold2295 (.A(net2796),
    .X(net3576));
 sky130_fd_sc_hd__buf_2 hold2296 (.A(net165),
    .X(net3577));
 sky130_fd_sc_hd__buf_2 hold2297 (.A(net2797),
    .X(net3578));
 sky130_fd_sc_hd__buf_2 hold23 (.A(net2850),
    .X(net1304));
 sky130_fd_sc_hd__buf_2 hold230 (.A(net1499),
    .X(net1511));
 sky130_fd_sc_hd__buf_2 hold2303 (.A(_0895_),
    .X(net3584));
 sky130_fd_sc_hd__buf_2 hold2304 (.A(net2938),
    .X(net3585));
 sky130_fd_sc_hd__buf_2 hold2305 (.A(net2366),
    .X(net3586));
 sky130_fd_sc_hd__buf_2 hold2306 (.A(net2939),
    .X(net3587));
 sky130_fd_sc_hd__buf_2 hold2307 (.A(net1998),
    .X(net3588));
 sky130_fd_sc_hd__buf_2 hold2308 (.A(net2940),
    .X(net3589));
 sky130_fd_sc_hd__buf_2 hold2309 (.A(net2367),
    .X(net3590));
 sky130_fd_sc_hd__buf_2 hold231 (.A(net1493),
    .X(net1512));
 sky130_fd_sc_hd__buf_2 hold2310 (.A(net2941),
    .X(net3591));
 sky130_fd_sc_hd__buf_2 hold2316 (.A(_0893_),
    .X(net3597));
 sky130_fd_sc_hd__buf_2 hold2317 (.A(net2947),
    .X(net3598));
 sky130_fd_sc_hd__buf_2 hold2318 (.A(net2373),
    .X(net3599));
 sky130_fd_sc_hd__buf_2 hold2319 (.A(net2948),
    .X(net3600));
 sky130_fd_sc_hd__buf_2 hold232 (.A(net1500),
    .X(net1513));
 sky130_fd_sc_hd__buf_2 hold2320 (.A(net2004),
    .X(net3601));
 sky130_fd_sc_hd__buf_2 hold2321 (.A(net2949),
    .X(net3602));
 sky130_fd_sc_hd__buf_2 hold2322 (.A(net2374),
    .X(net3603));
 sky130_fd_sc_hd__buf_2 hold2323 (.A(net2950),
    .X(net3604));
 sky130_fd_sc_hd__buf_2 hold2324 (.A(wbs_adr_i[9]),
    .X(net3605));
 sky130_fd_sc_hd__buf_2 hold2325 (.A(net2805),
    .X(net3606));
 sky130_fd_sc_hd__buf_2 hold2326 (.A(net2272),
    .X(net3607));
 sky130_fd_sc_hd__buf_2 hold2327 (.A(net2806),
    .X(net3608));
 sky130_fd_sc_hd__buf_2 hold2328 (.A(net1317),
    .X(net3609));
 sky130_fd_sc_hd__buf_2 hold2329 (.A(net2807),
    .X(net3610));
 sky130_fd_sc_hd__buf_2 hold233 (.A(_1247_),
    .X(net1514));
 sky130_fd_sc_hd__buf_2 hold2330 (.A(net2273),
    .X(net3611));
 sky130_fd_sc_hd__buf_2 hold2331 (.A(net2808),
    .X(net3612));
 sky130_fd_sc_hd__buf_2 hold2332 (.A(net166),
    .X(net3613));
 sky130_fd_sc_hd__buf_2 hold2333 (.A(net2809),
    .X(net3614));
 sky130_fd_sc_hd__buf_2 hold2339 (.A(_0894_),
    .X(net3620));
 sky130_fd_sc_hd__buf_2 hold234 (.A(wbs_sel_i[3]),
    .X(net1515));
 sky130_fd_sc_hd__buf_2 hold2340 (.A(net2973),
    .X(net3621));
 sky130_fd_sc_hd__buf_2 hold2341 (.A(net2387),
    .X(net3622));
 sky130_fd_sc_hd__buf_2 hold2342 (.A(net2974),
    .X(net3623));
 sky130_fd_sc_hd__buf_2 hold2343 (.A(net2029),
    .X(net3624));
 sky130_fd_sc_hd__buf_2 hold2344 (.A(net2975),
    .X(net3625));
 sky130_fd_sc_hd__buf_2 hold2345 (.A(net2388),
    .X(net3626));
 sky130_fd_sc_hd__buf_2 hold2346 (.A(net2976),
    .X(net3627));
 sky130_fd_sc_hd__buf_2 hold235 (.A(net1502),
    .X(net1516));
 sky130_fd_sc_hd__buf_2 hold2352 (.A(_0892_),
    .X(net3633));
 sky130_fd_sc_hd__buf_2 hold2353 (.A(net2956),
    .X(net3634));
 sky130_fd_sc_hd__buf_2 hold2354 (.A(net2394),
    .X(net3635));
 sky130_fd_sc_hd__buf_2 hold2355 (.A(net2957),
    .X(net3636));
 sky130_fd_sc_hd__buf_2 hold2356 (.A(net2047),
    .X(net3637));
 sky130_fd_sc_hd__buf_2 hold2357 (.A(net2958),
    .X(net3638));
 sky130_fd_sc_hd__buf_2 hold2358 (.A(net2395),
    .X(net3639));
 sky130_fd_sc_hd__buf_2 hold2359 (.A(net2959),
    .X(net3640));
 sky130_fd_sc_hd__buf_2 hold236 (.A(net1495),
    .X(net1517));
 sky130_fd_sc_hd__buf_2 hold2365 (.A(_0890_),
    .X(net3646));
 sky130_fd_sc_hd__buf_2 hold2366 (.A(net2982),
    .X(net3647));
 sky130_fd_sc_hd__buf_2 hold2367 (.A(net2380),
    .X(net3648));
 sky130_fd_sc_hd__buf_2 hold2368 (.A(net2983),
    .X(net3649));
 sky130_fd_sc_hd__buf_2 hold2369 (.A(net2035),
    .X(net3650));
 sky130_fd_sc_hd__buf_2 hold237 (.A(net1503),
    .X(net1518));
 sky130_fd_sc_hd__buf_2 hold2370 (.A(net2984),
    .X(net3651));
 sky130_fd_sc_hd__buf_2 hold2371 (.A(net2381),
    .X(net3652));
 sky130_fd_sc_hd__buf_2 hold2372 (.A(net2985),
    .X(net3653));
 sky130_fd_sc_hd__buf_2 hold2378 (.A(_0948_),
    .X(net3659));
 sky130_fd_sc_hd__buf_2 hold2379 (.A(net2999),
    .X(net3660));
 sky130_fd_sc_hd__buf_2 hold2380 (.A(net2413),
    .X(net3661));
 sky130_fd_sc_hd__buf_2 hold2381 (.A(net3000),
    .X(net3662));
 sky130_fd_sc_hd__buf_2 hold2382 (.A(net2190),
    .X(net3663));
 sky130_fd_sc_hd__buf_2 hold2383 (.A(net3001),
    .X(net3664));
 sky130_fd_sc_hd__buf_2 hold2384 (.A(net2414),
    .X(net3665));
 sky130_fd_sc_hd__buf_2 hold2385 (.A(net3002),
    .X(net3666));
 sky130_fd_sc_hd__buf_2 hold2386 (.A(wbs_adr_i[10]),
    .X(net3667));
 sky130_fd_sc_hd__buf_2 hold2387 (.A(net2817),
    .X(net3668));
 sky130_fd_sc_hd__buf_2 hold2388 (.A(net2266),
    .X(net3669));
 sky130_fd_sc_hd__buf_2 hold2389 (.A(net2818),
    .X(net3670));
 sky130_fd_sc_hd__buf_2 hold2390 (.A(net1287),
    .X(net3671));
 sky130_fd_sc_hd__buf_2 hold2391 (.A(net2819),
    .X(net3672));
 sky130_fd_sc_hd__buf_2 hold2392 (.A(net2267),
    .X(net3673));
 sky130_fd_sc_hd__buf_2 hold2393 (.A(net2820),
    .X(net3674));
 sky130_fd_sc_hd__buf_2 hold2394 (.A(net136),
    .X(net3675));
 sky130_fd_sc_hd__buf_2 hold2395 (.A(net2821),
    .X(net3676));
 sky130_fd_sc_hd__buf_2 hold24 (.A(net3540),
    .X(net1305));
 sky130_fd_sc_hd__buf_2 hold240 (.A(net3917),
    .X(net1521));
 sky130_fd_sc_hd__buf_2 hold2401 (.A(_0949_),
    .X(net3682));
 sky130_fd_sc_hd__buf_2 hold2402 (.A(net3008),
    .X(net3683));
 sky130_fd_sc_hd__buf_2 hold2403 (.A(net2420),
    .X(net3684));
 sky130_fd_sc_hd__buf_2 hold2404 (.A(net3009),
    .X(net3685));
 sky130_fd_sc_hd__buf_2 hold2405 (.A(net2184),
    .X(net3686));
 sky130_fd_sc_hd__buf_2 hold2406 (.A(net3010),
    .X(net3687));
 sky130_fd_sc_hd__buf_2 hold2407 (.A(net2421),
    .X(net3688));
 sky130_fd_sc_hd__buf_2 hold2408 (.A(net3011),
    .X(net3689));
 sky130_fd_sc_hd__buf_2 hold2409 (.A(wbs_adr_i[2]),
    .X(net3690));
 sky130_fd_sc_hd__buf_2 hold2410 (.A(net2841),
    .X(net3691));
 sky130_fd_sc_hd__buf_2 hold2411 (.A(net2284),
    .X(net3692));
 sky130_fd_sc_hd__buf_2 hold2412 (.A(net2842),
    .X(net3693));
 sky130_fd_sc_hd__buf_2 hold2413 (.A(net1302),
    .X(net3694));
 sky130_fd_sc_hd__buf_2 hold2414 (.A(net2843),
    .X(net3695));
 sky130_fd_sc_hd__buf_2 hold2415 (.A(net2285),
    .X(net3696));
 sky130_fd_sc_hd__buf_2 hold2416 (.A(net2844),
    .X(net3697));
 sky130_fd_sc_hd__buf_2 hold2417 (.A(net157),
    .X(net3698));
 sky130_fd_sc_hd__buf_2 hold2418 (.A(net2845),
    .X(net3699));
 sky130_fd_sc_hd__buf_2 hold2419 (.A(wbs_adr_i[11]),
    .X(net3700));
 sky130_fd_sc_hd__buf_2 hold2420 (.A(net2829),
    .X(net3701));
 sky130_fd_sc_hd__buf_2 hold2421 (.A(net2278),
    .X(net3702));
 sky130_fd_sc_hd__buf_2 hold2422 (.A(net2830),
    .X(net3703));
 sky130_fd_sc_hd__buf_2 hold2423 (.A(net1296),
    .X(net3704));
 sky130_fd_sc_hd__buf_2 hold2424 (.A(net2831),
    .X(net3705));
 sky130_fd_sc_hd__buf_2 hold2425 (.A(net2279),
    .X(net3706));
 sky130_fd_sc_hd__buf_2 hold2426 (.A(net2832),
    .X(net3707));
 sky130_fd_sc_hd__buf_2 hold2427 (.A(net137),
    .X(net3708));
 sky130_fd_sc_hd__buf_2 hold2428 (.A(net2833),
    .X(net3709));
 sky130_fd_sc_hd__buf_2 hold2429 (.A(wbs_adr_i[3]),
    .X(net3710));
 sky130_fd_sc_hd__buf_2 hold243 (.A(net3925),
    .X(net1524));
 sky130_fd_sc_hd__buf_2 hold2430 (.A(net2853),
    .X(net3711));
 sky130_fd_sc_hd__buf_2 hold2431 (.A(net2290),
    .X(net3712));
 sky130_fd_sc_hd__buf_2 hold2432 (.A(net2854),
    .X(net3713));
 sky130_fd_sc_hd__buf_2 hold2433 (.A(net1320),
    .X(net3714));
 sky130_fd_sc_hd__buf_2 hold2434 (.A(net2855),
    .X(net3715));
 sky130_fd_sc_hd__buf_2 hold2435 (.A(net2291),
    .X(net3716));
 sky130_fd_sc_hd__buf_2 hold2436 (.A(net2856),
    .X(net3717));
 sky130_fd_sc_hd__buf_2 hold2437 (.A(net160),
    .X(net3718));
 sky130_fd_sc_hd__buf_2 hold2438 (.A(net2857),
    .X(net3719));
 sky130_fd_sc_hd__buf_2 hold2439 (.A(wbs_adr_i[12]),
    .X(net3720));
 sky130_fd_sc_hd__buf_2 hold2440 (.A(net2865),
    .X(net3721));
 sky130_fd_sc_hd__buf_2 hold2441 (.A(net2302),
    .X(net3722));
 sky130_fd_sc_hd__buf_2 hold2442 (.A(net2866),
    .X(net3723));
 sky130_fd_sc_hd__buf_2 hold2443 (.A(net1326),
    .X(net3724));
 sky130_fd_sc_hd__buf_2 hold2444 (.A(net2867),
    .X(net3725));
 sky130_fd_sc_hd__buf_2 hold2445 (.A(net2303),
    .X(net3726));
 sky130_fd_sc_hd__buf_2 hold2446 (.A(net2868),
    .X(net3727));
 sky130_fd_sc_hd__buf_2 hold2447 (.A(net138),
    .X(net3728));
 sky130_fd_sc_hd__buf_2 hold2448 (.A(wbs_adr_i[13]),
    .X(net3729));
 sky130_fd_sc_hd__buf_2 hold2449 (.A(net2889),
    .X(net3730));
 sky130_fd_sc_hd__buf_2 hold245 (.A(net1554),
    .X(net1526));
 sky130_fd_sc_hd__buf_2 hold2450 (.A(net2308),
    .X(net3731));
 sky130_fd_sc_hd__buf_2 hold2451 (.A(net2890),
    .X(net3732));
 sky130_fd_sc_hd__buf_2 hold2452 (.A(net1329),
    .X(net3733));
 sky130_fd_sc_hd__buf_2 hold2453 (.A(net2891),
    .X(net3734));
 sky130_fd_sc_hd__buf_2 hold2454 (.A(net2309),
    .X(net3735));
 sky130_fd_sc_hd__buf_2 hold2455 (.A(net2892),
    .X(net3736));
 sky130_fd_sc_hd__buf_2 hold2456 (.A(net139),
    .X(net3737));
 sky130_fd_sc_hd__buf_2 hold2457 (.A(wbs_adr_i[14]),
    .X(net3738));
 sky130_fd_sc_hd__buf_2 hold2458 (.A(net2877),
    .X(net3739));
 sky130_fd_sc_hd__buf_2 hold2459 (.A(net2296),
    .X(net3740));
 sky130_fd_sc_hd__buf_2 hold246 (.A(_0994_),
    .X(net1527));
 sky130_fd_sc_hd__buf_2 hold2460 (.A(net2878),
    .X(net3741));
 sky130_fd_sc_hd__buf_2 hold2461 (.A(net1323),
    .X(net3742));
 sky130_fd_sc_hd__buf_2 hold2462 (.A(net2879),
    .X(net3743));
 sky130_fd_sc_hd__buf_2 hold2463 (.A(net2297),
    .X(net3744));
 sky130_fd_sc_hd__buf_2 hold2464 (.A(net2880),
    .X(net3745));
 sky130_fd_sc_hd__buf_2 hold2465 (.A(net140),
    .X(net3746));
 sky130_fd_sc_hd__buf_2 hold2471 (.A(net4125),
    .X(net3752));
 sky130_fd_sc_hd__buf_2 hold2472 (.A(net3043),
    .X(net3753));
 sky130_fd_sc_hd__buf_2 hold2473 (.A(net2535),
    .X(net3754));
 sky130_fd_sc_hd__buf_2 hold2474 (.A(net3044),
    .X(net3755));
 sky130_fd_sc_hd__buf_2 hold2475 (.A(net2091),
    .X(net3756));
 sky130_fd_sc_hd__buf_2 hold2476 (.A(net3045),
    .X(net3757));
 sky130_fd_sc_hd__buf_2 hold2477 (.A(net2536),
    .X(net3758));
 sky130_fd_sc_hd__buf_2 hold2478 (.A(net3046),
    .X(net3759));
 sky130_fd_sc_hd__buf_2 hold248 (.A(net1552),
    .X(net1529));
 sky130_fd_sc_hd__buf_2 hold2484 (.A(net4119),
    .X(net3765));
 sky130_fd_sc_hd__buf_2 hold2485 (.A(net3052),
    .X(net3766));
 sky130_fd_sc_hd__buf_2 hold2486 (.A(net2542),
    .X(net3767));
 sky130_fd_sc_hd__buf_2 hold2487 (.A(net3053),
    .X(net3768));
 sky130_fd_sc_hd__buf_2 hold2488 (.A(net2074),
    .X(net3769));
 sky130_fd_sc_hd__buf_2 hold2489 (.A(net3054),
    .X(net3770));
 sky130_fd_sc_hd__buf_2 hold249 (.A(net1556),
    .X(net1530));
 sky130_fd_sc_hd__buf_2 hold2490 (.A(net2543),
    .X(net3771));
 sky130_fd_sc_hd__buf_2 hold2491 (.A(net3055),
    .X(net3772));
 sky130_fd_sc_hd__buf_2 hold2497 (.A(net4131),
    .X(net3778));
 sky130_fd_sc_hd__buf_2 hold2498 (.A(net3061),
    .X(net3779));
 sky130_fd_sc_hd__buf_2 hold2499 (.A(net2549),
    .X(net3780));
 sky130_fd_sc_hd__buf_2 hold25 (.A(net2774),
    .X(net1306));
 sky130_fd_sc_hd__buf_2 hold250 (.A(_0993_),
    .X(net1531));
 sky130_fd_sc_hd__buf_2 hold2500 (.A(net3062),
    .X(net3781));
 sky130_fd_sc_hd__buf_2 hold2501 (.A(net2080),
    .X(net3782));
 sky130_fd_sc_hd__buf_2 hold2502 (.A(net3063),
    .X(net3783));
 sky130_fd_sc_hd__buf_2 hold2503 (.A(net2550),
    .X(net3784));
 sky130_fd_sc_hd__buf_2 hold2504 (.A(net3064),
    .X(net3785));
 sky130_fd_sc_hd__buf_2 hold2510 (.A(net4137),
    .X(net3791));
 sky130_fd_sc_hd__buf_2 hold2511 (.A(net3079),
    .X(net3792));
 sky130_fd_sc_hd__buf_2 hold2512 (.A(net2563),
    .X(net3793));
 sky130_fd_sc_hd__buf_2 hold2513 (.A(net3080),
    .X(net3794));
 sky130_fd_sc_hd__buf_2 hold2514 (.A(net2097),
    .X(net3795));
 sky130_fd_sc_hd__buf_2 hold2515 (.A(net3081),
    .X(net3796));
 sky130_fd_sc_hd__buf_2 hold2516 (.A(net2564),
    .X(net3797));
 sky130_fd_sc_hd__buf_2 hold2517 (.A(net3082),
    .X(net3798));
 sky130_fd_sc_hd__buf_2 hold2523 (.A(net4149),
    .X(net3804));
 sky130_fd_sc_hd__buf_2 hold2524 (.A(net3070),
    .X(net3805));
 sky130_fd_sc_hd__buf_2 hold2525 (.A(net2556),
    .X(net3806));
 sky130_fd_sc_hd__buf_2 hold2526 (.A(net3071),
    .X(net3807));
 sky130_fd_sc_hd__buf_2 hold2527 (.A(net2114),
    .X(net3808));
 sky130_fd_sc_hd__buf_2 hold2528 (.A(net3072),
    .X(net3809));
 sky130_fd_sc_hd__buf_2 hold2529 (.A(net2557),
    .X(net3810));
 sky130_fd_sc_hd__buf_2 hold253 (.A(net3946),
    .X(net1534));
 sky130_fd_sc_hd__buf_2 hold2530 (.A(net3073),
    .X(net3811));
 sky130_fd_sc_hd__buf_2 hold2536 (.A(net4143),
    .X(net3817));
 sky130_fd_sc_hd__buf_2 hold2537 (.A(net3088),
    .X(net3818));
 sky130_fd_sc_hd__buf_2 hold2538 (.A(net2570),
    .X(net3819));
 sky130_fd_sc_hd__buf_2 hold2539 (.A(net3089),
    .X(net3820));
 sky130_fd_sc_hd__buf_2 hold2540 (.A(net2129),
    .X(net3821));
 sky130_fd_sc_hd__buf_2 hold2541 (.A(net3090),
    .X(net3822));
 sky130_fd_sc_hd__buf_2 hold2542 (.A(net2571),
    .X(net3823));
 sky130_fd_sc_hd__buf_2 hold2543 (.A(net3091),
    .X(net3824));
 sky130_fd_sc_hd__buf_2 hold2549 (.A(net4156),
    .X(net3830));
 sky130_fd_sc_hd__buf_2 hold255 (.A(net1551),
    .X(net1536));
 sky130_fd_sc_hd__buf_2 hold2550 (.A(net3025),
    .X(net3831));
 sky130_fd_sc_hd__buf_2 hold2551 (.A(net2466),
    .X(net3832));
 sky130_fd_sc_hd__buf_2 hold2552 (.A(net3026),
    .X(net3833));
 sky130_fd_sc_hd__buf_2 hold2553 (.A(net1793),
    .X(net3834));
 sky130_fd_sc_hd__buf_2 hold2554 (.A(net3027),
    .X(net3835));
 sky130_fd_sc_hd__buf_2 hold2555 (.A(net2467),
    .X(net3836));
 sky130_fd_sc_hd__buf_2 hold2556 (.A(net3028),
    .X(net3837));
 sky130_fd_sc_hd__buf_2 hold256 (.A(net1553),
    .X(net1537));
 sky130_fd_sc_hd__buf_2 hold2562 (.A(_0951_),
    .X(net3843));
 sky130_fd_sc_hd__buf_2 hold2563 (.A(net3034),
    .X(net3844));
 sky130_fd_sc_hd__buf_2 hold2564 (.A(net2473),
    .X(net3845));
 sky130_fd_sc_hd__buf_2 hold2565 (.A(net3035),
    .X(net3846));
 sky130_fd_sc_hd__buf_2 hold2566 (.A(net1829),
    .X(net3847));
 sky130_fd_sc_hd__buf_2 hold2567 (.A(net3036),
    .X(net3848));
 sky130_fd_sc_hd__buf_2 hold2568 (.A(net2474),
    .X(net3849));
 sky130_fd_sc_hd__buf_2 hold2569 (.A(net3037),
    .X(net3850));
 sky130_fd_sc_hd__buf_2 hold257 (.A(net1555),
    .X(net1538));
 sky130_fd_sc_hd__buf_2 hold2572 (.A(_0922_),
    .X(net3853));
 sky130_fd_sc_hd__buf_2 hold2573 (.A(net3094),
    .X(net3854));
 sky130_fd_sc_hd__buf_2 hold2574 (.A(net2574),
    .X(net3855));
 sky130_fd_sc_hd__buf_2 hold2575 (.A(net3095),
    .X(net3856));
 sky130_fd_sc_hd__buf_2 hold2576 (.A(net1484),
    .X(net3857));
 sky130_fd_sc_hd__buf_2 hold2577 (.A(net3096),
    .X(net3858));
 sky130_fd_sc_hd__buf_2 hold2578 (.A(net2575),
    .X(net3859));
 sky130_fd_sc_hd__buf_2 hold2579 (.A(net3097),
    .X(net3860));
 sky130_fd_sc_hd__buf_2 hold258 (.A(net1557),
    .X(net1539));
 sky130_fd_sc_hd__buf_2 hold2582 (.A(net645),
    .X(net3863));
 sky130_fd_sc_hd__buf_2 hold2583 (.A(_0925_),
    .X(net3864));
 sky130_fd_sc_hd__buf_2 hold2584 (.A(net3135),
    .X(net3865));
 sky130_fd_sc_hd__buf_2 hold2585 (.A(net2579),
    .X(net3866));
 sky130_fd_sc_hd__buf_2 hold2586 (.A(net3136),
    .X(net3867));
 sky130_fd_sc_hd__buf_2 hold2587 (.A(net1664),
    .X(net3868));
 sky130_fd_sc_hd__buf_2 hold2588 (.A(net3137),
    .X(net3869));
 sky130_fd_sc_hd__buf_2 hold259 (.A(_0990_),
    .X(net1540));
 sky130_fd_sc_hd__buf_2 hold2590 (.A(_2431_),
    .X(net3871));
 sky130_fd_sc_hd__buf_2 hold2591 (.A(net2925),
    .X(net3872));
 sky130_fd_sc_hd__buf_2 hold2592 (.A(net2318),
    .X(net3873));
 sky130_fd_sc_hd__buf_2 hold2593 (.A(net2926),
    .X(net3874));
 sky130_fd_sc_hd__buf_2 hold2594 (.A(net1486),
    .X(net3875));
 sky130_fd_sc_hd__buf_2 hold2595 (.A(net2927),
    .X(net3876));
 sky130_fd_sc_hd__buf_2 hold2596 (.A(net2319),
    .X(net3877));
 sky130_fd_sc_hd__buf_2 hold26 (.A(net2778),
    .X(net1307));
 sky130_fd_sc_hd__buf_2 hold2604 (.A(_0897_),
    .X(net3885));
 sky130_fd_sc_hd__buf_2 hold2605 (.A(net3256),
    .X(net3886));
 sky130_fd_sc_hd__buf_2 hold2606 (.A(net2595),
    .X(net3887));
 sky130_fd_sc_hd__buf_2 hold2607 (.A(net3257),
    .X(net3888));
 sky130_fd_sc_hd__buf_2 hold2608 (.A(net2063),
    .X(net3889));
 sky130_fd_sc_hd__buf_2 hold2609 (.A(net3258),
    .X(net3890));
 sky130_fd_sc_hd__buf_2 hold2617 (.A(_0896_),
    .X(net3898));
 sky130_fd_sc_hd__buf_2 hold2618 (.A(net3267),
    .X(net3899));
 sky130_fd_sc_hd__buf_2 hold2619 (.A(net2604),
    .X(net3900));
 sky130_fd_sc_hd__buf_2 hold262 (.A(net3954),
    .X(net1543));
 sky130_fd_sc_hd__buf_2 hold2620 (.A(net3268),
    .X(net3901));
 sky130_fd_sc_hd__buf_2 hold2621 (.A(net2055),
    .X(net3902));
 sky130_fd_sc_hd__buf_2 hold2622 (.A(net3269),
    .X(net3903));
 sky130_fd_sc_hd__buf_2 hold2625 (.A(_0941_),
    .X(net3906));
 sky130_fd_sc_hd__buf_2 hold2626 (.A(net3273),
    .X(net3907));
 sky130_fd_sc_hd__buf_2 hold2627 (.A(net2586),
    .X(net3908));
 sky130_fd_sc_hd__buf_2 hold2628 (.A(net3274),
    .X(net3909));
 sky130_fd_sc_hd__buf_2 hold2629 (.A(net1740),
    .X(net3910));
 sky130_fd_sc_hd__buf_2 hold2630 (.A(net3275),
    .X(net3911));
 sky130_fd_sc_hd__buf_2 hold2633 (.A(_0981_),
    .X(net3914));
 sky130_fd_sc_hd__buf_2 hold2634 (.A(net3279),
    .X(net3915));
 sky130_fd_sc_hd__buf_2 hold2635 (.A(net2608),
    .X(net3916));
 sky130_fd_sc_hd__buf_2 hold2636 (.A(net3280),
    .X(net3917));
 sky130_fd_sc_hd__buf_2 hold2637 (.A(net1521),
    .X(net3918));
 sky130_fd_sc_hd__buf_2 hold2638 (.A(net3281),
    .X(net3919));
 sky130_fd_sc_hd__buf_2 hold2641 (.A(_0983_),
    .X(net3922));
 sky130_fd_sc_hd__buf_2 hold2642 (.A(net3285),
    .X(net3923));
 sky130_fd_sc_hd__buf_2 hold2643 (.A(net2612),
    .X(net3924));
 sky130_fd_sc_hd__buf_2 hold2644 (.A(net3286),
    .X(net3925));
 sky130_fd_sc_hd__buf_2 hold2645 (.A(net1524),
    .X(net3926));
 sky130_fd_sc_hd__buf_2 hold2646 (.A(net3287),
    .X(net3927));
 sky130_fd_sc_hd__buf_2 hold265 (.A(net3962),
    .X(net1546));
 sky130_fd_sc_hd__buf_2 hold2654 (.A(_1333_),
    .X(net3935));
 sky130_fd_sc_hd__buf_2 hold2655 (.A(net3302),
    .X(net3936));
 sky130_fd_sc_hd__buf_2 hold2656 (.A(net2633),
    .X(net3937));
 sky130_fd_sc_hd__buf_2 hold2657 (.A(net3303),
    .X(net3938));
 sky130_fd_sc_hd__buf_2 hold2658 (.A(net1963),
    .X(net3939));
 sky130_fd_sc_hd__buf_2 hold2659 (.A(net3304),
    .X(net3940));
 sky130_fd_sc_hd__buf_2 hold2662 (.A(_0982_),
    .X(net3943));
 sky130_fd_sc_hd__buf_2 hold2663 (.A(net3291),
    .X(net3944));
 sky130_fd_sc_hd__buf_2 hold2664 (.A(net2616),
    .X(net3945));
 sky130_fd_sc_hd__buf_2 hold2665 (.A(net3292),
    .X(net3946));
 sky130_fd_sc_hd__buf_2 hold2666 (.A(net1534),
    .X(net3947));
 sky130_fd_sc_hd__buf_2 hold2667 (.A(net3293),
    .X(net3948));
 sky130_fd_sc_hd__buf_2 hold267 (.A(net1635),
    .X(net1548));
 sky130_fd_sc_hd__buf_2 hold2670 (.A(_0978_),
    .X(net3951));
 sky130_fd_sc_hd__buf_2 hold2671 (.A(net3308),
    .X(net3952));
 sky130_fd_sc_hd__buf_2 hold2672 (.A(net2620),
    .X(net3953));
 sky130_fd_sc_hd__buf_2 hold2673 (.A(net3309),
    .X(net3954));
 sky130_fd_sc_hd__buf_2 hold2674 (.A(net1543),
    .X(net3955));
 sky130_fd_sc_hd__buf_2 hold2675 (.A(net3310),
    .X(net3956));
 sky130_fd_sc_hd__buf_2 hold2678 (.A(_0980_),
    .X(net3959));
 sky130_fd_sc_hd__buf_2 hold2679 (.A(net3314),
    .X(net3960));
 sky130_fd_sc_hd__buf_2 hold268 (.A(_0998_),
    .X(net1549));
 sky130_fd_sc_hd__buf_2 hold2680 (.A(net2624),
    .X(net3961));
 sky130_fd_sc_hd__buf_2 hold2681 (.A(net3315),
    .X(net3962));
 sky130_fd_sc_hd__buf_2 hold2682 (.A(net1546),
    .X(net3963));
 sky130_fd_sc_hd__buf_2 hold2683 (.A(net3316),
    .X(net3964));
 sky130_fd_sc_hd__buf_2 hold2686 (.A(_0979_),
    .X(net3967));
 sky130_fd_sc_hd__buf_2 hold2687 (.A(net3320),
    .X(net3968));
 sky130_fd_sc_hd__buf_2 hold2688 (.A(net2637),
    .X(net3969));
 sky130_fd_sc_hd__buf_2 hold2689 (.A(net3321),
    .X(net3970));
 sky130_fd_sc_hd__buf_2 hold2690 (.A(net1572),
    .X(net3971));
 sky130_fd_sc_hd__buf_2 hold2691 (.A(net3322),
    .X(net3972));
 sky130_fd_sc_hd__buf_2 hold2694 (.A(_0984_),
    .X(net3975));
 sky130_fd_sc_hd__buf_2 hold2695 (.A(net3337),
    .X(net3976));
 sky130_fd_sc_hd__buf_2 hold2696 (.A(net2641),
    .X(net3977));
 sky130_fd_sc_hd__buf_2 hold2697 (.A(net3338),
    .X(net3978));
 sky130_fd_sc_hd__buf_2 hold2698 (.A(net1658),
    .X(net3979));
 sky130_fd_sc_hd__buf_2 hold27 (.A(net3572),
    .X(net1308));
 sky130_fd_sc_hd__buf_2 hold270 (.A(net1648),
    .X(net1551));
 sky130_fd_sc_hd__buf_2 hold2706 (.A(_1334_),
    .X(net3987));
 sky130_fd_sc_hd__buf_2 hold2707 (.A(net3348),
    .X(net3988));
 sky130_fd_sc_hd__buf_2 hold2708 (.A(net2694),
    .X(net3989));
 sky130_fd_sc_hd__buf_2 hold2709 (.A(net3349),
    .X(net3990));
 sky130_fd_sc_hd__buf_2 hold271 (.A(net1536),
    .X(net1552));
 sky130_fd_sc_hd__buf_2 hold2712 (.A(net3998),
    .X(net3993));
 sky130_fd_sc_hd__buf_2 hold2713 (.A(_0975_),
    .X(net3994));
 sky130_fd_sc_hd__buf_2 hold2714 (.A(net3355),
    .X(net3995));
 sky130_fd_sc_hd__buf_2 hold2717 (.A(net4001),
    .X(net3998));
 sky130_fd_sc_hd__buf_2 hold272 (.A(net1529),
    .X(net1553));
 sky130_fd_sc_hd__buf_2 hold2720 (.A(net642),
    .X(net4001));
 sky130_fd_sc_hd__buf_2 hold273 (.A(net1537),
    .X(net1554));
 sky130_fd_sc_hd__buf_2 hold2730 (.A(_2408_),
    .X(net4011));
 sky130_fd_sc_hd__buf_2 hold2731 (.A(net3101),
    .X(net4012));
 sky130_fd_sc_hd__buf_2 hold2735 (.A(_2411_),
    .X(net4016));
 sky130_fd_sc_hd__buf_2 hold2736 (.A(net3124),
    .X(net4017));
 sky130_fd_sc_hd__buf_2 hold2739 (.A(net1472),
    .X(net4020));
 sky130_fd_sc_hd__buf_2 hold274 (.A(net1526),
    .X(net1555));
 sky130_fd_sc_hd__buf_2 hold2740 (.A(net3111),
    .X(net4021));
 sky130_fd_sc_hd__buf_2 hold2744 (.A(_2412_),
    .X(net4025));
 sky130_fd_sc_hd__buf_2 hold2748 (.A(_2420_),
    .X(net4029));
 sky130_fd_sc_hd__buf_2 hold275 (.A(net1538),
    .X(net1556));
 sky130_fd_sc_hd__buf_2 hold2752 (.A(_2416_),
    .X(net4033));
 sky130_fd_sc_hd__buf_2 hold2756 (.A(_2419_),
    .X(net4037));
 sky130_fd_sc_hd__buf_2 hold276 (.A(net1530),
    .X(net1557));
 sky130_fd_sc_hd__buf_2 hold2760 (.A(_2415_),
    .X(net4041));
 sky130_fd_sc_hd__buf_2 hold2764 (.A(_2409_),
    .X(net4045));
 sky130_fd_sc_hd__buf_2 hold2768 (.A(_2410_),
    .X(net4049));
 sky130_fd_sc_hd__buf_2 hold277 (.A(net1539),
    .X(net1558));
 sky130_fd_sc_hd__buf_2 hold2772 (.A(_2414_),
    .X(net4053));
 sky130_fd_sc_hd__buf_2 hold2778 (.A(_2121_),
    .X(net4059));
 sky130_fd_sc_hd__buf_2 hold278 (.A(_0995_),
    .X(net1559));
 sky130_fd_sc_hd__buf_2 hold2787 (.A(net4165),
    .X(net4068));
 sky130_fd_sc_hd__buf_2 hold2788 (.A(net4167),
    .X(net4069));
 sky130_fd_sc_hd__buf_2 hold2789 (.A(net4169),
    .X(net4070));
 sky130_fd_sc_hd__buf_2 hold2790 (.A(net3453),
    .X(net4071));
 sky130_fd_sc_hd__buf_2 hold2791 (.A(net2316),
    .X(net4072));
 sky130_fd_sc_hd__buf_2 hold2792 (.A(net3454),
    .X(net4073));
 sky130_fd_sc_hd__buf_2 hold2793 (.A(net2744),
    .X(net4074));
 sky130_fd_sc_hd__buf_2 hold2794 (.A(net3455),
    .X(net4075));
 sky130_fd_sc_hd__buf_2 hold2796 (.A(_0924_),
    .X(net4077));
 sky130_fd_sc_hd__buf_2 hold2797 (.A(net3463),
    .X(net4078));
 sky130_fd_sc_hd__buf_2 hold2798 (.A(net2902),
    .X(net4079));
 sky130_fd_sc_hd__buf_2 hold2799 (.A(net3464),
    .X(net4080));
 sky130_fd_sc_hd__buf_2 hold28 (.A(net2798),
    .X(net1309));
 sky130_fd_sc_hd__buf_2 hold280 (.A(net1633),
    .X(net1561));
 sky130_fd_sc_hd__buf_2 hold2800 (.A(net2349),
    .X(net4081));
 sky130_fd_sc_hd__buf_2 hold2801 (.A(net3465),
    .X(net4082));
 sky130_fd_sc_hd__buf_2 hold2803 (.A(_0985_),
    .X(net4084));
 sky130_fd_sc_hd__buf_2 hold2804 (.A(net3472),
    .X(net4085));
 sky130_fd_sc_hd__buf_2 hold2805 (.A(net2920),
    .X(net4086));
 sky130_fd_sc_hd__buf_2 hold2806 (.A(net3473),
    .X(net4087));
 sky130_fd_sc_hd__buf_2 hold2807 (.A(net2359),
    .X(net4088));
 sky130_fd_sc_hd__buf_2 hold281 (.A(net1637),
    .X(net1562));
 sky130_fd_sc_hd__buf_2 hold2812 (.A(_1313_),
    .X(net4093));
 sky130_fd_sc_hd__buf_2 hold2813 (.A(net3507),
    .X(net4094));
 sky130_fd_sc_hd__buf_2 hold2814 (.A(net2990),
    .X(net4095));
 sky130_fd_sc_hd__buf_2 hold2819 (.A(_1312_),
    .X(net4100));
 sky130_fd_sc_hd__buf_2 hold282 (.A(_0996_),
    .X(net1563));
 sky130_fd_sc_hd__buf_2 hold2820 (.A(net3495),
    .X(net4101));
 sky130_fd_sc_hd__buf_2 hold2821 (.A(net2964),
    .X(net4102));
 sky130_fd_sc_hd__buf_2 hold2825 (.A(_0954_),
    .X(net4106));
 sky130_fd_sc_hd__buf_2 hold2826 (.A(net3483),
    .X(net4107));
 sky130_fd_sc_hd__buf_2 hold2831 (.A(_0581_),
    .X(net4112));
 sky130_fd_sc_hd__buf_2 hold2832 (.A(net3561),
    .X(net4113));
 sky130_fd_sc_hd__buf_2 hold2838 (.A(_1307_),
    .X(net4119));
 sky130_fd_sc_hd__buf_2 hold284 (.A(net1632),
    .X(net1565));
 sky130_fd_sc_hd__buf_2 hold2844 (.A(_1306_),
    .X(net4125));
 sky130_fd_sc_hd__buf_2 hold285 (.A(net1634),
    .X(net1566));
 sky130_fd_sc_hd__buf_2 hold2850 (.A(_1308_),
    .X(net4131));
 sky130_fd_sc_hd__buf_2 hold2856 (.A(_1311_),
    .X(net4137));
 sky130_fd_sc_hd__buf_2 hold286 (.A(net1636),
    .X(net1567));
 sky130_fd_sc_hd__buf_2 hold2862 (.A(_1309_),
    .X(net4143));
 sky130_fd_sc_hd__buf_2 hold2868 (.A(_1310_),
    .X(net4149));
 sky130_fd_sc_hd__buf_2 hold2869 (.A(net1483),
    .X(net4150));
 sky130_fd_sc_hd__buf_2 hold287 (.A(net1638),
    .X(net1568));
 sky130_fd_sc_hd__buf_2 hold2875 (.A(_0953_),
    .X(net4156));
 sky130_fd_sc_hd__buf_2 hold288 (.A(_0997_),
    .X(net1569));
 sky130_fd_sc_hd__buf_2 hold2883 (.A(_0891_),
    .X(net4164));
 sky130_fd_sc_hd__buf_2 hold2884 (.A(net1465),
    .X(net4165));
 sky130_fd_sc_hd__buf_2 hold2885 (.A(net4068),
    .X(net4166));
 sky130_fd_sc_hd__buf_2 hold2886 (.A(net3452),
    .X(net4167));
 sky130_fd_sc_hd__buf_2 hold2887 (.A(net4069),
    .X(net4168));
 sky130_fd_sc_hd__buf_2 hold2888 (.A(net2743),
    .X(net4169));
 sky130_fd_sc_hd__buf_2 hold2889 (.A(_1405_),
    .X(net4170));
 sky130_fd_sc_hd__buf_2 hold2890 (.A(net4187),
    .X(net4171));
 sky130_fd_sc_hd__buf_2 hold2893 (.A(net4185),
    .X(net4174));
 sky130_fd_sc_hd__buf_2 hold2894 (.A(net4189),
    .X(net4175));
 sky130_fd_sc_hd__buf_2 hold2897 (.A(net4184),
    .X(net4178));
 sky130_fd_sc_hd__buf_2 hold2898 (.A(net4186),
    .X(net4179));
 sky130_fd_sc_hd__buf_2 hold2899 (.A(net4188),
    .X(net4180));
 sky130_fd_sc_hd__buf_2 hold29 (.A(net2802),
    .X(net1310));
 sky130_fd_sc_hd__buf_2 hold2900 (.A(net4175),
    .X(net4181));
 sky130_fd_sc_hd__buf_2 hold2903 (.A(_0950_),
    .X(net4184));
 sky130_fd_sc_hd__buf_2 hold2904 (.A(net4178),
    .X(net4185));
 sky130_fd_sc_hd__buf_2 hold2905 (.A(net4174),
    .X(net4186));
 sky130_fd_sc_hd__buf_2 hold2906 (.A(net4179),
    .X(net4187));
 sky130_fd_sc_hd__buf_2 hold2907 (.A(net4171),
    .X(net4188));
 sky130_fd_sc_hd__buf_2 hold2908 (.A(net4180),
    .X(net4189));
 sky130_fd_sc_hd__buf_2 hold291 (.A(net3970),
    .X(net1572));
 sky130_fd_sc_hd__buf_2 hold292 (.A(net3324),
    .X(net1573));
 sky130_fd_sc_hd__buf_2 hold293 (.A(net3326),
    .X(net1574));
 sky130_fd_sc_hd__buf_2 hold294 (.A(net1459),
    .X(net1575));
 sky130_fd_sc_hd__buf_2 hold295 (.A(net1469),
    .X(net1576));
 sky130_fd_sc_hd__buf_2 hold296 (.A(net204),
    .X(net1577));
 sky130_fd_sc_hd__buf_2 hold297 (.A(net1470),
    .X(net1578));
 sky130_fd_sc_hd__buf_2 hold298 (.A(net1460),
    .X(net1579));
 sky130_fd_sc_hd__buf_2 hold299 (.A(net1471),
    .X(net1580));
 sky130_fd_sc_hd__buf_2 hold30 (.A(net3550),
    .X(net1311));
 sky130_fd_sc_hd__buf_2 hold300 (.A(_2119_),
    .X(net1581));
 sky130_fd_sc_hd__buf_2 hold301 (.A(_2120_),
    .X(net1582));
 sky130_fd_sc_hd__buf_2 hold302 (.A(net1600),
    .X(net1583));
 sky130_fd_sc_hd__buf_2 hold303 (.A(_1091_),
    .X(net1584));
 sky130_fd_sc_hd__buf_2 hold308 (.A(net1609),
    .X(net1589));
 sky130_fd_sc_hd__buf_2 hold309 (.A(net1599),
    .X(net1590));
 sky130_fd_sc_hd__buf_2 hold31 (.A(net2786),
    .X(net1312));
 sky130_fd_sc_hd__buf_2 hold310 (.A(net1601),
    .X(net1591));
 sky130_fd_sc_hd__buf_2 hold311 (.A(_1093_),
    .X(net1592));
 sky130_fd_sc_hd__buf_2 hold316 (.A(net1608),
    .X(net1597));
 sky130_fd_sc_hd__buf_2 hold317 (.A(net1589),
    .X(net1598));
 sky130_fd_sc_hd__buf_2 hold318 (.A(net424),
    .X(net1599));
 sky130_fd_sc_hd__buf_2 hold319 (.A(net1590),
    .X(net1600));
 sky130_fd_sc_hd__buf_2 hold32 (.A(net2790),
    .X(net1313));
 sky130_fd_sc_hd__buf_2 hold320 (.A(net1583),
    .X(net1601));
 sky130_fd_sc_hd__buf_2 hold321 (.A(net1591),
    .X(net1602));
 sky130_fd_sc_hd__buf_2 hold322 (.A(_1095_),
    .X(net1603));
 sky130_fd_sc_hd__buf_2 hold327 (.A(net1582),
    .X(net1608));
 sky130_fd_sc_hd__buf_2 hold328 (.A(net1597),
    .X(net1609));
 sky130_fd_sc_hd__buf_2 hold33 (.A(net1447),
    .X(net1314));
 sky130_fd_sc_hd__buf_2 hold34 (.A(net1455),
    .X(net1315));
 sky130_fd_sc_hd__buf_2 hold348 (.A(net1653),
    .X(net1629));
 sky130_fd_sc_hd__buf_2 hold349 (.A(net491),
    .X(net1630));
 sky130_fd_sc_hd__buf_2 hold35 (.A(_1279_),
    .X(net1316));
 sky130_fd_sc_hd__buf_2 hold351 (.A(net1655),
    .X(net1632));
 sky130_fd_sc_hd__buf_2 hold352 (.A(net1565),
    .X(net1633));
 sky130_fd_sc_hd__buf_2 hold353 (.A(net1561),
    .X(net1634));
 sky130_fd_sc_hd__buf_2 hold354 (.A(net1566),
    .X(net1635));
 sky130_fd_sc_hd__buf_2 hold355 (.A(net1548),
    .X(net1636));
 sky130_fd_sc_hd__buf_2 hold356 (.A(net1567),
    .X(net1637));
 sky130_fd_sc_hd__buf_2 hold357 (.A(net1562),
    .X(net1638));
 sky130_fd_sc_hd__buf_2 hold358 (.A(net1568),
    .X(net1639));
 sky130_fd_sc_hd__buf_2 hold359 (.A(_1001_),
    .X(net1640));
 sky130_fd_sc_hd__buf_2 hold36 (.A(net3608),
    .X(net1317));
 sky130_fd_sc_hd__buf_2 hold363 (.A(net1652),
    .X(net1644));
 sky130_fd_sc_hd__buf_2 hold364 (.A(net1629),
    .X(net1645));
 sky130_fd_sc_hd__buf_2 hold365 (.A(_0999_),
    .X(net1646));
 sky130_fd_sc_hd__buf_2 hold367 (.A(net648),
    .X(net1648));
 sky130_fd_sc_hd__buf_2 hold37 (.A(net2810),
    .X(net1318));
 sky130_fd_sc_hd__buf_2 hold371 (.A(_2037_),
    .X(net1652));
 sky130_fd_sc_hd__buf_2 hold372 (.A(net1644),
    .X(net1653));
 sky130_fd_sc_hd__buf_2 hold374 (.A(net1660),
    .X(net1655));
 sky130_fd_sc_hd__buf_2 hold377 (.A(net3978),
    .X(net1658));
 sky130_fd_sc_hd__buf_2 hold379 (.A(net649),
    .X(net1660));
 sky130_fd_sc_hd__buf_2 hold38 (.A(net2814),
    .X(net1319));
 sky130_fd_sc_hd__buf_2 hold383 (.A(net3867),
    .X(net1664));
 sky130_fd_sc_hd__buf_2 hold386 (.A(net1680),
    .X(net1667));
 sky130_fd_sc_hd__buf_2 hold387 (.A(net1684),
    .X(net1668));
 sky130_fd_sc_hd__buf_2 hold388 (.A(_1192_),
    .X(net1669));
 sky130_fd_sc_hd__buf_2 hold39 (.A(net3713),
    .X(net1320));
 sky130_fd_sc_hd__buf_2 hold391 (.A(net1679),
    .X(net1672));
 sky130_fd_sc_hd__buf_2 hold392 (.A(net1681),
    .X(net1673));
 sky130_fd_sc_hd__buf_2 hold393 (.A(net1683),
    .X(net1674));
 sky130_fd_sc_hd__buf_2 hold394 (.A(net1685),
    .X(net1675));
 sky130_fd_sc_hd__buf_2 hold395 (.A(_1193_),
    .X(net1676));
 sky130_fd_sc_hd__buf_2 hold398 (.A(net1689),
    .X(net1679));
 sky130_fd_sc_hd__buf_2 hold399 (.A(net1672),
    .X(net1680));
 sky130_fd_sc_hd__buf_2 hold40 (.A(net2858),
    .X(net1321));
 sky130_fd_sc_hd__buf_2 hold400 (.A(net1667),
    .X(net1681));
 sky130_fd_sc_hd__buf_2 hold401 (.A(net1673),
    .X(net1682));
 sky130_fd_sc_hd__buf_2 hold402 (.A(net1490),
    .X(net1683));
 sky130_fd_sc_hd__buf_2 hold403 (.A(net1674),
    .X(net1684));
 sky130_fd_sc_hd__buf_2 hold404 (.A(net1668),
    .X(net1685));
 sky130_fd_sc_hd__buf_2 hold405 (.A(net1675),
    .X(net1686));
 sky130_fd_sc_hd__buf_2 hold408 (.A(_0561_),
    .X(net1689));
 sky130_fd_sc_hd__buf_2 hold41 (.A(net2862),
    .X(net1322));
 sky130_fd_sc_hd__buf_2 hold415 (.A(net2729),
    .X(net1696));
 sky130_fd_sc_hd__buf_2 hold416 (.A(net2732),
    .X(net1697));
 sky130_fd_sc_hd__buf_2 hold42 (.A(net3741),
    .X(net1323));
 sky130_fd_sc_hd__buf_2 hold425 (.A(net1783),
    .X(net1706));
 sky130_fd_sc_hd__buf_2 hold426 (.A(_0874_),
    .X(net1707));
 sky130_fd_sc_hd__buf_2 hold43 (.A(net2882),
    .X(net1324));
 sky130_fd_sc_hd__buf_2 hold431 (.A(net1781),
    .X(net1712));
 sky130_fd_sc_hd__buf_2 hold432 (.A(net1785),
    .X(net1713));
 sky130_fd_sc_hd__buf_2 hold433 (.A(_0875_),
    .X(net1714));
 sky130_fd_sc_hd__buf_2 hold437 (.A(net3356),
    .X(net1718));
 sky130_fd_sc_hd__buf_2 hold44 (.A(net2886),
    .X(net1325));
 sky130_fd_sc_hd__buf_2 hold441 (.A(net3370),
    .X(net1722));
 sky130_fd_sc_hd__buf_2 hold445 (.A(net3363),
    .X(net1726));
 sky130_fd_sc_hd__buf_2 hold449 (.A(net3377),
    .X(net1730));
 sky130_fd_sc_hd__buf_2 hold45 (.A(net3723),
    .X(net1326));
 sky130_fd_sc_hd__buf_2 hold452 (.A(net2737),
    .X(net1733));
 sky130_fd_sc_hd__buf_2 hold453 (.A(net2730),
    .X(net1734));
 sky130_fd_sc_hd__buf_2 hold454 (.A(_0973_),
    .X(net1735));
 sky130_fd_sc_hd__buf_2 hold458 (.A(net2584),
    .X(net1739));
 sky130_fd_sc_hd__buf_2 hold459 (.A(net3909),
    .X(net1740));
 sky130_fd_sc_hd__buf_2 hold46 (.A(net2870),
    .X(net1327));
 sky130_fd_sc_hd__buf_2 hold463 (.A(net3384),
    .X(net1744));
 sky130_fd_sc_hd__buf_2 hold468 (.A(net2105),
    .X(net1749));
 sky130_fd_sc_hd__buf_2 hold469 (.A(_2426_),
    .X(net1750));
 sky130_fd_sc_hd__buf_2 hold47 (.A(net2874),
    .X(net1328));
 sky130_fd_sc_hd__buf_2 hold470 (.A(_0947_),
    .X(net1751));
 sky130_fd_sc_hd__buf_2 hold474 (.A(net3391),
    .X(net1755));
 sky130_fd_sc_hd__buf_2 hold479 (.A(net1780),
    .X(net1760));
 sky130_fd_sc_hd__buf_2 hold48 (.A(net3732),
    .X(net1329));
 sky130_fd_sc_hd__buf_2 hold480 (.A(net1782),
    .X(net1761));
 sky130_fd_sc_hd__buf_2 hold481 (.A(net1784),
    .X(net1762));
 sky130_fd_sc_hd__buf_2 hold482 (.A(net1786),
    .X(net1763));
 sky130_fd_sc_hd__buf_2 hold483 (.A(net421),
    .X(net1764));
 sky130_fd_sc_hd__buf_2 hold484 (.A(_0878_),
    .X(net1765));
 sky130_fd_sc_hd__buf_2 hold488 (.A(net3398),
    .X(net1769));
 sky130_fd_sc_hd__buf_2 hold489 (.A(net3402),
    .X(net1770));
 sky130_fd_sc_hd__buf_2 hold49 (.A(net2894),
    .X(net1330));
 sky130_fd_sc_hd__buf_2 hold493 (.A(net3407),
    .X(net1774));
 sky130_fd_sc_hd__buf_2 hold494 (.A(net3411),
    .X(net1775));
 sky130_fd_sc_hd__buf_2 hold499 (.A(net1798),
    .X(net1780));
 sky130_fd_sc_hd__buf_2 hold50 (.A(net2898),
    .X(net1331));
 sky130_fd_sc_hd__buf_2 hold500 (.A(net1760),
    .X(net1781));
 sky130_fd_sc_hd__buf_2 hold501 (.A(net1712),
    .X(net1782));
 sky130_fd_sc_hd__buf_2 hold502 (.A(net1761),
    .X(net1783));
 sky130_fd_sc_hd__buf_2 hold503 (.A(net1706),
    .X(net1784));
 sky130_fd_sc_hd__buf_2 hold504 (.A(net1762),
    .X(net1785));
 sky130_fd_sc_hd__buf_2 hold505 (.A(net1713),
    .X(net1786));
 sky130_fd_sc_hd__buf_2 hold506 (.A(net1763),
    .X(net1787));
 sky130_fd_sc_hd__buf_2 hold51 (.A(net1406),
    .X(net1332));
 sky130_fd_sc_hd__buf_2 hold512 (.A(net3833),
    .X(net1793));
 sky130_fd_sc_hd__buf_2 hold517 (.A(_2129_),
    .X(net1798));
 sky130_fd_sc_hd__buf_2 hold52 (.A(net1414),
    .X(net1333));
 sky130_fd_sc_hd__buf_2 hold521 (.A(net3416),
    .X(net1802));
 sky130_fd_sc_hd__buf_2 hold522 (.A(net3420),
    .X(net1803));
 sky130_fd_sc_hd__buf_2 hold525 (.A(net1860),
    .X(net1806));
 sky130_fd_sc_hd__buf_2 hold526 (.A(_2087_),
    .X(net1807));
 sky130_fd_sc_hd__buf_2 hold527 (.A(_1058_),
    .X(net1808));
 sky130_fd_sc_hd__buf_2 hold53 (.A(_1280_),
    .X(net1334));
 sky130_fd_sc_hd__buf_2 hold534 (.A(net1858),
    .X(net1815));
 sky130_fd_sc_hd__buf_2 hold535 (.A(net1834),
    .X(net1816));
 sky130_fd_sc_hd__buf_2 hold536 (.A(_2096_),
    .X(net1817));
 sky130_fd_sc_hd__buf_2 hold537 (.A(_1060_),
    .X(net1818));
 sky130_fd_sc_hd__buf_2 hold54 (.A(net1364),
    .X(net1335));
 sky130_fd_sc_hd__buf_2 hold541 (.A(net3425),
    .X(net1822));
 sky130_fd_sc_hd__buf_2 hold542 (.A(net3429),
    .X(net1823));
 sky130_fd_sc_hd__buf_2 hold548 (.A(net3846),
    .X(net1829));
 sky130_fd_sc_hd__buf_2 hold55 (.A(net1368),
    .X(net1336));
 sky130_fd_sc_hd__buf_2 hold551 (.A(net1857),
    .X(net1832));
 sky130_fd_sc_hd__buf_2 hold552 (.A(net1859),
    .X(net1833));
 sky130_fd_sc_hd__buf_2 hold553 (.A(net1861),
    .X(net1834));
 sky130_fd_sc_hd__buf_2 hold554 (.A(net1816),
    .X(net1835));
 sky130_fd_sc_hd__buf_2 hold555 (.A(_2099_),
    .X(net1836));
 sky130_fd_sc_hd__buf_2 hold556 (.A(_1061_),
    .X(net1837));
 sky130_fd_sc_hd__buf_2 hold56 (.A(net1372),
    .X(net1337));
 sky130_fd_sc_hd__buf_2 hold560 (.A(net3434),
    .X(net1841));
 sky130_fd_sc_hd__buf_2 hold561 (.A(net3438),
    .X(net1842));
 sky130_fd_sc_hd__buf_2 hold57 (.A(net1376),
    .X(net1338));
 sky130_fd_sc_hd__buf_2 hold570 (.A(net2103),
    .X(net1851));
 sky130_fd_sc_hd__buf_2 hold571 (.A(net2107),
    .X(net1852));
 sky130_fd_sc_hd__buf_2 hold572 (.A(net2020),
    .X(net1853));
 sky130_fd_sc_hd__buf_2 hold573 (.A(_0762_),
    .X(net1854));
 sky130_fd_sc_hd__buf_2 hold576 (.A(net1880),
    .X(net1857));
 sky130_fd_sc_hd__buf_2 hold577 (.A(net1832),
    .X(net1858));
 sky130_fd_sc_hd__buf_2 hold578 (.A(net1815),
    .X(net1859));
 sky130_fd_sc_hd__buf_2 hold579 (.A(net1833),
    .X(net1860));
 sky130_fd_sc_hd__buf_2 hold58 (.A(net1359),
    .X(net1339));
 sky130_fd_sc_hd__buf_2 hold580 (.A(net1806),
    .X(net1861));
 sky130_fd_sc_hd__buf_2 hold584 (.A(net3153),
    .X(net1865));
 sky130_fd_sc_hd__buf_2 hold585 (.A(net3157),
    .X(net1866));
 sky130_fd_sc_hd__buf_2 hold589 (.A(net3208),
    .X(net1870));
 sky130_fd_sc_hd__buf_2 hold59 (.A(_1005_),
    .X(net1340));
 sky130_fd_sc_hd__buf_2 hold590 (.A(net3212),
    .X(net1871));
 sky130_fd_sc_hd__buf_2 hold594 (.A(net2040),
    .X(net1875));
 sky130_fd_sc_hd__buf_2 hold595 (.A(net2021),
    .X(net1876));
 sky130_fd_sc_hd__buf_2 hold596 (.A(_0763_),
    .X(net1877));
 sky130_fd_sc_hd__buf_2 hold599 (.A(net646),
    .X(net1880));
 sky130_fd_sc_hd__buf_2 hold6 (.A(net3670),
    .X(net1287));
 sky130_fd_sc_hd__buf_2 hold60 (.A(net650),
    .X(net1341));
 sky130_fd_sc_hd__buf_2 hold61 (.A(net3466),
    .X(net1342));
 sky130_fd_sc_hd__buf_2 hold62 (.A(net1363),
    .X(net1343));
 sky130_fd_sc_hd__buf_2 hold628 (.A(net3498),
    .X(net1909));
 sky130_fd_sc_hd__buf_2 hold63 (.A(net1365),
    .X(net1344));
 sky130_fd_sc_hd__buf_2 hold64 (.A(net1367),
    .X(net1345));
 sky130_fd_sc_hd__buf_2 hold641 (.A(net3510),
    .X(net1922));
 sky130_fd_sc_hd__buf_2 hold65 (.A(net1369),
    .X(net1346));
 sky130_fd_sc_hd__buf_2 hold66 (.A(net1371),
    .X(net1347));
 sky130_fd_sc_hd__buf_2 hold662 (.A(net3564),
    .X(net1943));
 sky130_fd_sc_hd__buf_2 hold666 (.A(net2014),
    .X(net1947));
 sky130_fd_sc_hd__buf_2 hold667 (.A(net1983),
    .X(net1948));
 sky130_fd_sc_hd__buf_2 hold668 (.A(_0739_),
    .X(net1949));
 sky130_fd_sc_hd__buf_2 hold67 (.A(net1373),
    .X(net1348));
 sky130_fd_sc_hd__buf_2 hold672 (.A(net2154),
    .X(net1953));
 sky130_fd_sc_hd__buf_2 hold673 (.A(net1991),
    .X(net1954));
 sky130_fd_sc_hd__buf_2 hold674 (.A(_1076_),
    .X(net1955));
 sky130_fd_sc_hd__buf_2 hold675 (.A(net1485),
    .X(net1956));
 sky130_fd_sc_hd__buf_2 hold68 (.A(net1375),
    .X(net1349));
 sky130_fd_sc_hd__buf_2 hold682 (.A(net3938),
    .X(net1963));
 sky130_fd_sc_hd__buf_2 hold687 (.A(net2102),
    .X(net1968));
 sky130_fd_sc_hd__buf_2 hold688 (.A(net2104),
    .X(net1969));
 sky130_fd_sc_hd__buf_2 hold689 (.A(net2106),
    .X(net1970));
 sky130_fd_sc_hd__buf_2 hold69 (.A(net1377),
    .X(net1350));
 sky130_fd_sc_hd__buf_2 hold690 (.A(net1852),
    .X(net1971));
 sky130_fd_sc_hd__buf_2 hold691 (.A(_2424_),
    .X(net1972));
 sky130_fd_sc_hd__buf_2 hold692 (.A(_0946_),
    .X(net1973));
 sky130_fd_sc_hd__buf_2 hold696 (.A(net3486),
    .X(net1977));
 sky130_fd_sc_hd__buf_2 hold7 (.A(net2822),
    .X(net1288));
 sky130_fd_sc_hd__buf_2 hold70 (.A(net1380),
    .X(net1351));
 sky130_fd_sc_hd__buf_2 hold700 (.A(net2013),
    .X(net1981));
 sky130_fd_sc_hd__buf_2 hold701 (.A(net2015),
    .X(net1982));
 sky130_fd_sc_hd__buf_2 hold702 (.A(net428),
    .X(net1983));
 sky130_fd_sc_hd__buf_2 hold703 (.A(net1948),
    .X(net1984));
 sky130_fd_sc_hd__buf_2 hold704 (.A(_0740_),
    .X(net1985));
 sky130_fd_sc_hd__buf_2 hold708 (.A(net2153),
    .X(net1989));
 sky130_fd_sc_hd__buf_2 hold709 (.A(net2155),
    .X(net1990));
 sky130_fd_sc_hd__buf_2 hold71 (.A(net1360),
    .X(net1352));
 sky130_fd_sc_hd__buf_2 hold710 (.A(net633),
    .X(net1991));
 sky130_fd_sc_hd__buf_2 hold711 (.A(net1954),
    .X(net1992));
 sky130_fd_sc_hd__buf_2 hold717 (.A(net3587),
    .X(net1998));
 sky130_fd_sc_hd__buf_2 hold72 (.A(_1006_),
    .X(net1353));
 sky130_fd_sc_hd__buf_2 hold723 (.A(net3600),
    .X(net2004));
 sky130_fd_sc_hd__buf_2 hold727 (.A(net3102),
    .X(net2008));
 sky130_fd_sc_hd__buf_2 hold728 (.A(net3106),
    .X(net2009));
 sky130_fd_sc_hd__buf_2 hold73 (.A(net1341),
    .X(net1354));
 sky130_fd_sc_hd__buf_2 hold732 (.A(_2045_),
    .X(net2013));
 sky130_fd_sc_hd__buf_2 hold733 (.A(net1981),
    .X(net2014));
 sky130_fd_sc_hd__buf_2 hold734 (.A(net1947),
    .X(net2015));
 sky130_fd_sc_hd__buf_2 hold738 (.A(net2039),
    .X(net2019));
 sky130_fd_sc_hd__buf_2 hold739 (.A(net2041),
    .X(net2020));
 sky130_fd_sc_hd__buf_2 hold74 (.A(net644),
    .X(net1355));
 sky130_fd_sc_hd__buf_2 hold740 (.A(net1853),
    .X(net2021));
 sky130_fd_sc_hd__buf_2 hold741 (.A(net1876),
    .X(net2022));
 sky130_fd_sc_hd__buf_2 hold742 (.A(net429),
    .X(net2023));
 sky130_fd_sc_hd__buf_2 hold748 (.A(net3623),
    .X(net2029));
 sky130_fd_sc_hd__buf_2 hold754 (.A(net3649),
    .X(net2035));
 sky130_fd_sc_hd__buf_2 hold758 (.A(_2044_),
    .X(net2039));
 sky130_fd_sc_hd__buf_2 hold759 (.A(net2019),
    .X(net2040));
 sky130_fd_sc_hd__buf_2 hold76 (.A(net1421),
    .X(net1357));
 sky130_fd_sc_hd__buf_2 hold760 (.A(net1875),
    .X(net2041));
 sky130_fd_sc_hd__buf_2 hold766 (.A(net3636),
    .X(net2047));
 sky130_fd_sc_hd__buf_2 hold77 (.A(net1379),
    .X(net1358));
 sky130_fd_sc_hd__buf_2 hold774 (.A(net3901),
    .X(net2055));
 sky130_fd_sc_hd__buf_2 hold78 (.A(net1351),
    .X(net1359));
 sky130_fd_sc_hd__buf_2 hold782 (.A(net3888),
    .X(net2063));
 sky130_fd_sc_hd__buf_2 hold786 (.A(net3125),
    .X(net2067));
 sky130_fd_sc_hd__buf_2 hold787 (.A(net3129),
    .X(net2068));
 sky130_fd_sc_hd__buf_2 hold79 (.A(net1339),
    .X(net1360));
 sky130_fd_sc_hd__buf_2 hold793 (.A(net3768),
    .X(net2074));
 sky130_fd_sc_hd__buf_2 hold799 (.A(net3781),
    .X(net2080));
 sky130_fd_sc_hd__buf_2 hold8 (.A(net2826),
    .X(net1289));
 sky130_fd_sc_hd__buf_2 hold80 (.A(net1352),
    .X(net1361));
 sky130_fd_sc_hd__buf_2 hold803 (.A(net3230),
    .X(net2084));
 sky130_fd_sc_hd__buf_2 hold804 (.A(net3234),
    .X(net2085));
 sky130_fd_sc_hd__buf_2 hold81 (.A(_1010_),
    .X(net1362));
 sky130_fd_sc_hd__buf_2 hold810 (.A(net3755),
    .X(net2091));
 sky130_fd_sc_hd__buf_2 hold816 (.A(net3794),
    .X(net2097));
 sky130_fd_sc_hd__buf_2 hold82 (.A(wbs_sel_i[0]),
    .X(net1363));
 sky130_fd_sc_hd__buf_2 hold821 (.A(net485),
    .X(net2102));
 sky130_fd_sc_hd__buf_2 hold822 (.A(net1968),
    .X(net2103));
 sky130_fd_sc_hd__buf_2 hold823 (.A(net1851),
    .X(net2104));
 sky130_fd_sc_hd__buf_2 hold824 (.A(net1969),
    .X(net2105));
 sky130_fd_sc_hd__buf_2 hold825 (.A(net1749),
    .X(net2106));
 sky130_fd_sc_hd__buf_2 hold826 (.A(net1970),
    .X(net2107));
 sky130_fd_sc_hd__buf_2 hold827 (.A(_0944_),
    .X(net2108));
 sky130_fd_sc_hd__buf_2 hold83 (.A(net1343),
    .X(net1364));
 sky130_fd_sc_hd__buf_2 hold833 (.A(net3807),
    .X(net2114));
 sky130_fd_sc_hd__buf_2 hold84 (.A(net1335),
    .X(net1365));
 sky130_fd_sc_hd__buf_2 hold841 (.A(net3175),
    .X(net2122));
 sky130_fd_sc_hd__buf_2 hold842 (.A(net3179),
    .X(net2123));
 sky130_fd_sc_hd__buf_2 hold848 (.A(net3820),
    .X(net2129));
 sky130_fd_sc_hd__buf_2 hold85 (.A(net1344),
    .X(net1366));
 sky130_fd_sc_hd__buf_2 hold852 (.A(net3197),
    .X(net2133));
 sky130_fd_sc_hd__buf_2 hold853 (.A(net3201),
    .X(net2134));
 sky130_fd_sc_hd__buf_2 hold857 (.A(net3186),
    .X(net2138));
 sky130_fd_sc_hd__buf_2 hold858 (.A(net3190),
    .X(net2139));
 sky130_fd_sc_hd__buf_2 hold86 (.A(net1290),
    .X(net1367));
 sky130_fd_sc_hd__buf_2 hold862 (.A(net3219),
    .X(net2143));
 sky130_fd_sc_hd__buf_2 hold863 (.A(net3223),
    .X(net2144));
 sky130_fd_sc_hd__buf_2 hold867 (.A(net3164),
    .X(net2148));
 sky130_fd_sc_hd__buf_2 hold868 (.A(net3168),
    .X(net2149));
 sky130_fd_sc_hd__buf_2 hold87 (.A(net1345),
    .X(net1368));
 sky130_fd_sc_hd__buf_2 hold872 (.A(net2160),
    .X(net2153));
 sky130_fd_sc_hd__buf_2 hold873 (.A(net1989),
    .X(net2154));
 sky130_fd_sc_hd__buf_2 hold874 (.A(net1953),
    .X(net2155));
 sky130_fd_sc_hd__buf_2 hold875 (.A(net1990),
    .X(net2156));
 sky130_fd_sc_hd__buf_2 hold879 (.A(_1374_),
    .X(net2160));
 sky130_fd_sc_hd__buf_2 hold88 (.A(net1336),
    .X(net1369));
 sky130_fd_sc_hd__buf_2 hold89 (.A(net1346),
    .X(net1370));
 sky130_fd_sc_hd__buf_2 hold9 (.A(net1366),
    .X(net1290));
 sky130_fd_sc_hd__buf_2 hold90 (.A(net200),
    .X(net1371));
 sky130_fd_sc_hd__buf_2 hold903 (.A(net3685),
    .X(net2184));
 sky130_fd_sc_hd__buf_2 hold909 (.A(net3662),
    .X(net2190));
 sky130_fd_sc_hd__buf_2 hold91 (.A(net1347),
    .X(net1372));
 sky130_fd_sc_hd__buf_2 hold92 (.A(net1337),
    .X(net1373));
 sky130_fd_sc_hd__buf_2 hold929 (.A(net3990),
    .X(net2210));
 sky130_fd_sc_hd__buf_2 hold93 (.A(net1348),
    .X(net1374));
 sky130_fd_sc_hd__buf_2 hold94 (.A(net1291),
    .X(net1375));
 sky130_fd_sc_hd__buf_2 hold95 (.A(net1349),
    .X(net1376));
 sky130_fd_sc_hd__buf_2 hold953 (.A(net3445),
    .X(net2234));
 sky130_fd_sc_hd__buf_2 hold954 (.A(net3449),
    .X(net2235));
 sky130_fd_sc_hd__buf_2 hold955 (.A(net3516),
    .X(net2236));
 sky130_fd_sc_hd__buf_2 hold956 (.A(net3520),
    .X(net2237));
 sky130_fd_sc_hd__buf_2 hold957 (.A(net3524),
    .X(net2238));
 sky130_fd_sc_hd__buf_2 hold958 (.A(net2751),
    .X(net2239));
 sky130_fd_sc_hd__buf_2 hold959 (.A(net2753),
    .X(net2240));
 sky130_fd_sc_hd__buf_2 hold96 (.A(net1338),
    .X(net1377));
 sky130_fd_sc_hd__buf_2 hold960 (.A(net2755),
    .X(net2241));
 sky130_fd_sc_hd__buf_2 hold961 (.A(net3527),
    .X(net2242));
 sky130_fd_sc_hd__buf_2 hold962 (.A(net3531),
    .X(net2243));
 sky130_fd_sc_hd__buf_2 hold963 (.A(net3535),
    .X(net2244));
 sky130_fd_sc_hd__buf_2 hold964 (.A(net2763),
    .X(net2245));
 sky130_fd_sc_hd__buf_2 hold965 (.A(net2765),
    .X(net2246));
 sky130_fd_sc_hd__buf_2 hold966 (.A(net2767),
    .X(net2247));
 sky130_fd_sc_hd__buf_2 hold967 (.A(net3538),
    .X(net2248));
 sky130_fd_sc_hd__buf_2 hold968 (.A(net3542),
    .X(net2249));
 sky130_fd_sc_hd__buf_2 hold969 (.A(net3546),
    .X(net2250));
 sky130_fd_sc_hd__buf_2 hold97 (.A(net1350),
    .X(net1378));
 sky130_fd_sc_hd__buf_2 hold970 (.A(net2775),
    .X(net2251));
 sky130_fd_sc_hd__buf_2 hold971 (.A(net2777),
    .X(net2252));
 sky130_fd_sc_hd__buf_2 hold972 (.A(net2779),
    .X(net2253));
 sky130_fd_sc_hd__buf_2 hold973 (.A(net3548),
    .X(net2254));
 sky130_fd_sc_hd__buf_2 hold974 (.A(net3552),
    .X(net2255));
 sky130_fd_sc_hd__buf_2 hold975 (.A(net3556),
    .X(net2256));
 sky130_fd_sc_hd__buf_2 hold976 (.A(net2787),
    .X(net2257));
 sky130_fd_sc_hd__buf_2 hold977 (.A(net2789),
    .X(net2258));
 sky130_fd_sc_hd__buf_2 hold978 (.A(net2791),
    .X(net2259));
 sky130_fd_sc_hd__buf_2 hold979 (.A(net3570),
    .X(net2260));
 sky130_fd_sc_hd__buf_2 hold98 (.A(_2038_),
    .X(net1379));
 sky130_fd_sc_hd__buf_2 hold980 (.A(net3574),
    .X(net2261));
 sky130_fd_sc_hd__buf_2 hold981 (.A(net3578),
    .X(net2262));
 sky130_fd_sc_hd__buf_2 hold982 (.A(net2799),
    .X(net2263));
 sky130_fd_sc_hd__buf_2 hold983 (.A(net2801),
    .X(net2264));
 sky130_fd_sc_hd__buf_2 hold984 (.A(net2803),
    .X(net2265));
 sky130_fd_sc_hd__buf_2 hold985 (.A(net3668),
    .X(net2266));
 sky130_fd_sc_hd__buf_2 hold986 (.A(net3672),
    .X(net2267));
 sky130_fd_sc_hd__buf_2 hold987 (.A(net3676),
    .X(net2268));
 sky130_fd_sc_hd__buf_2 hold988 (.A(net2823),
    .X(net2269));
 sky130_fd_sc_hd__buf_2 hold989 (.A(net2825),
    .X(net2270));
 sky130_fd_sc_hd__buf_2 hold99 (.A(net1358),
    .X(net1380));
 sky130_fd_sc_hd__buf_2 hold990 (.A(net2827),
    .X(net2271));
 sky130_fd_sc_hd__buf_2 hold991 (.A(net3606),
    .X(net2272));
 sky130_fd_sc_hd__buf_2 hold992 (.A(net3610),
    .X(net2273));
 sky130_fd_sc_hd__buf_2 hold993 (.A(net3614),
    .X(net2274));
 sky130_fd_sc_hd__buf_2 hold994 (.A(net2811),
    .X(net2275));
 sky130_fd_sc_hd__buf_2 hold995 (.A(net2813),
    .X(net2276));
 sky130_fd_sc_hd__buf_2 hold996 (.A(net2815),
    .X(net2277));
 sky130_fd_sc_hd__buf_2 hold997 (.A(net3701),
    .X(net2278));
 sky130_fd_sc_hd__buf_2 hold998 (.A(net3705),
    .X(net2279));
 sky130_fd_sc_hd__buf_2 hold999 (.A(net3709),
    .X(net2280));
 sky130_fd_sc_hd__buf_4 input1 (.A(caravel_uart_rx),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(caravel_wb_data_i[16]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(probe_out[68]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(probe_out[69]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(probe_out[6]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(probe_out[70]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(probe_out[71]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(probe_out[72]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(probe_out[73]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(probe_out[74]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(probe_out[75]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(probe_out[76]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(caravel_wb_data_i[17]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(probe_out[77]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(probe_out[78]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 input112 (.A(probe_out[79]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 input113 (.A(probe_out[7]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(probe_out[80]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(probe_out[81]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(probe_out[82]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(probe_out[83]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(probe_out[84]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(probe_out[85]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(caravel_wb_data_i[18]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(probe_out[86]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(probe_out[87]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(probe_out[88]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(probe_out[89]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(probe_out[8]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(probe_out[90]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(probe_out[91]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(probe_out[92]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(probe_out[93]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(probe_out[94]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(caravel_wb_data_i[19]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(probe_out[95]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(probe_out[96]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(probe_out[97]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(probe_out[9]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input134 (.A(wb_rst_i),
    .X(net134));
 sky130_fd_sc_hd__buf_4 input135 (.A(wbs_adr_i[0]),
    .X(net135));
 sky130_fd_sc_hd__buf_6 input136 (.A(net3674),
    .X(net136));
 sky130_fd_sc_hd__buf_6 input137 (.A(net3707),
    .X(net137));
 sky130_fd_sc_hd__buf_4 input138 (.A(net3727),
    .X(net138));
 sky130_fd_sc_hd__buf_4 input139 (.A(net3736),
    .X(net139));
 sky130_fd_sc_hd__buf_2 input14 (.A(caravel_wb_data_i[1]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input140 (.A(net3745),
    .X(net140));
 sky130_fd_sc_hd__buf_6 input141 (.A(wbs_adr_i[15]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(wbs_adr_i[16]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(wbs_adr_i[17]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 input144 (.A(wbs_adr_i[18]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(wbs_adr_i[19]),
    .X(net145));
 sky130_fd_sc_hd__buf_4 input146 (.A(wbs_adr_i[1]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(wbs_adr_i[20]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 input148 (.A(wbs_adr_i[21]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 input149 (.A(wbs_adr_i[22]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(caravel_wb_data_i[20]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input150 (.A(wbs_adr_i[23]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 input151 (.A(wbs_adr_i[24]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 input152 (.A(wbs_adr_i[25]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 input153 (.A(wbs_adr_i[26]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 input154 (.A(wbs_adr_i[27]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 input155 (.A(wbs_adr_i[28]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 input156 (.A(wbs_adr_i[29]),
    .X(net156));
 sky130_fd_sc_hd__buf_4 input157 (.A(net3697),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 input158 (.A(wbs_adr_i[30]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 input159 (.A(wbs_adr_i[31]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(caravel_wb_data_i[21]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input160 (.A(net3717),
    .X(net160));
 sky130_fd_sc_hd__buf_4 input161 (.A(net3522),
    .X(net161));
 sky130_fd_sc_hd__buf_4 input162 (.A(net3533),
    .X(net162));
 sky130_fd_sc_hd__buf_4 input163 (.A(net3544),
    .X(net163));
 sky130_fd_sc_hd__buf_4 input164 (.A(net3554),
    .X(net164));
 sky130_fd_sc_hd__buf_4 input165 (.A(net3576),
    .X(net165));
 sky130_fd_sc_hd__buf_4 input166 (.A(net3612),
    .X(net166));
 sky130_fd_sc_hd__buf_6 input167 (.A(wbs_cyc_i),
    .X(net167));
 sky130_fd_sc_hd__buf_8 input168 (.A(wbs_data_i[0]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 input169 (.A(wbs_data_i[10]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(caravel_wb_data_i[22]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_8 input170 (.A(wbs_data_i[11]),
    .X(net170));
 sky130_fd_sc_hd__buf_4 input171 (.A(wbs_data_i[12]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_8 input172 (.A(wbs_data_i[13]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_8 input173 (.A(wbs_data_i[14]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_8 input174 (.A(wbs_data_i[15]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_8 input175 (.A(wbs_data_i[16]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_8 input176 (.A(wbs_data_i[17]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_8 input177 (.A(wbs_data_i[18]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_8 input178 (.A(wbs_data_i[19]),
    .X(net178));
 sky130_fd_sc_hd__buf_8 input179 (.A(wbs_data_i[1]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(caravel_wb_data_i[23]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_8 input180 (.A(wbs_data_i[20]),
    .X(net180));
 sky130_fd_sc_hd__buf_4 input181 (.A(wbs_data_i[21]),
    .X(net181));
 sky130_fd_sc_hd__buf_4 input182 (.A(wbs_data_i[22]),
    .X(net182));
 sky130_fd_sc_hd__buf_4 input183 (.A(wbs_data_i[23]),
    .X(net183));
 sky130_fd_sc_hd__buf_4 input184 (.A(wbs_data_i[24]),
    .X(net184));
 sky130_fd_sc_hd__buf_4 input185 (.A(wbs_data_i[25]),
    .X(net185));
 sky130_fd_sc_hd__buf_4 input186 (.A(wbs_data_i[26]),
    .X(net186));
 sky130_fd_sc_hd__buf_4 input187 (.A(wbs_data_i[27]),
    .X(net187));
 sky130_fd_sc_hd__buf_4 input188 (.A(wbs_data_i[28]),
    .X(net188));
 sky130_fd_sc_hd__buf_4 input189 (.A(wbs_data_i[29]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(caravel_wb_data_i[24]),
    .X(net19));
 sky130_fd_sc_hd__buf_6 input190 (.A(wbs_data_i[2]),
    .X(net190));
 sky130_fd_sc_hd__buf_4 input191 (.A(wbs_data_i[30]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_8 input192 (.A(wbs_data_i[31]),
    .X(net192));
 sky130_fd_sc_hd__buf_6 input193 (.A(wbs_data_i[3]),
    .X(net193));
 sky130_fd_sc_hd__buf_6 input194 (.A(wbs_data_i[4]),
    .X(net194));
 sky130_fd_sc_hd__buf_6 input195 (.A(wbs_data_i[5]),
    .X(net195));
 sky130_fd_sc_hd__buf_6 input196 (.A(wbs_data_i[6]),
    .X(net196));
 sky130_fd_sc_hd__buf_6 input197 (.A(wbs_data_i[7]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 input198 (.A(wbs_data_i[8]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_8 input199 (.A(wbs_data_i[9]),
    .X(net199));
 sky130_fd_sc_hd__buf_2 input2 (.A(caravel_wb_ack_i),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(caravel_wb_data_i[25]),
    .X(net20));
 sky130_fd_sc_hd__buf_8 input200 (.A(net1370),
    .X(net200));
 sky130_fd_sc_hd__buf_8 input201 (.A(net1451),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_16 input202 (.A(net1410),
    .X(net202));
 sky130_fd_sc_hd__buf_4 input203 (.A(net1505),
    .X(net203));
 sky130_fd_sc_hd__buf_6 input204 (.A(net1576),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_8 input205 (.A(net2325),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(caravel_wb_data_i[26]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(caravel_wb_data_i[27]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(caravel_wb_data_i[28]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(caravel_wb_data_i[29]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(caravel_wb_data_i[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(caravel_wb_data_i[30]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(caravel_wb_data_i[31]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(caravel_wb_data_i[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(caravel_wb_data_i[4]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input3 (.A(caravel_wb_data_i[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(caravel_wb_data_i[5]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(caravel_wb_data_i[6]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(caravel_wb_data_i[7]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(caravel_wb_data_i[8]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(caravel_wb_data_i[9]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(caravel_wb_error_i),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(probe_out[0]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(probe_out[10]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(probe_out[11]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(probe_out[12]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(caravel_wb_data_i[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(probe_out[13]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(probe_out[14]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(probe_out[15]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(probe_out[16]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(probe_out[17]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(probe_out[18]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(probe_out[19]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(probe_out[1]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(probe_out[20]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(probe_out[21]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(caravel_wb_data_i[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(probe_out[22]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(probe_out[23]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(probe_out[24]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(probe_out[25]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(probe_out[26]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(probe_out[27]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(probe_out[28]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(probe_out[29]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(probe_out[2]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(probe_out[30]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(caravel_wb_data_i[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(probe_out[31]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(probe_out[32]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(probe_out[33]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(probe_out[34]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(probe_out[35]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(probe_out[36]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(probe_out[37]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(probe_out[38]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(probe_out[39]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(probe_out[3]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input7 (.A(caravel_wb_data_i[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(probe_out[40]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(probe_out[41]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(probe_out[42]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(probe_out[43]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(probe_out[44]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(probe_out[45]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input76 (.A(probe_out[46]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(probe_out[47]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(probe_out[48]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(probe_out[49]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input8 (.A(caravel_wb_data_i[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(probe_out[4]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(probe_out[50]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(probe_out[51]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(probe_out[52]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(probe_out[53]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(probe_out[54]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(probe_out[55]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(probe_out[56]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(probe_out[57]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(probe_out[58]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(caravel_wb_data_i[15]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(probe_out[59]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 input91 (.A(probe_out[5]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(probe_out[60]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(probe_out[61]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(probe_out[62]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(probe_out[63]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(probe_out[64]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(probe_out[65]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(probe_out[66]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(probe_out[67]),
    .X(net99));
 sky130_fd_sc_hd__buf_12 max_cap405 (.A(_1461_),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_2 max_cap458 (.A(_1441_),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_2 max_cap459 (.A(_1441_),
    .X(net459));
 sky130_fd_sc_hd__buf_2 max_cap460 (.A(_2406_),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_2 output206 (.A(net206),
    .X(caravel_uart_tx));
 sky130_fd_sc_hd__clkbuf_2 output207 (.A(net207),
    .X(caravel_wb_adr_o[0]));
 sky130_fd_sc_hd__clkbuf_2 output208 (.A(net208),
    .X(caravel_wb_adr_o[10]));
 sky130_fd_sc_hd__clkbuf_2 output209 (.A(net209),
    .X(caravel_wb_adr_o[11]));
 sky130_fd_sc_hd__clkbuf_2 output210 (.A(net210),
    .X(caravel_wb_adr_o[12]));
 sky130_fd_sc_hd__clkbuf_2 output211 (.A(net211),
    .X(caravel_wb_adr_o[13]));
 sky130_fd_sc_hd__clkbuf_2 output212 (.A(net212),
    .X(caravel_wb_adr_o[14]));
 sky130_fd_sc_hd__clkbuf_2 output213 (.A(net213),
    .X(caravel_wb_adr_o[15]));
 sky130_fd_sc_hd__clkbuf_2 output214 (.A(net214),
    .X(caravel_wb_adr_o[16]));
 sky130_fd_sc_hd__clkbuf_2 output215 (.A(net215),
    .X(caravel_wb_adr_o[17]));
 sky130_fd_sc_hd__clkbuf_2 output216 (.A(net216),
    .X(caravel_wb_adr_o[18]));
 sky130_fd_sc_hd__clkbuf_2 output217 (.A(net217),
    .X(caravel_wb_adr_o[19]));
 sky130_fd_sc_hd__clkbuf_2 output218 (.A(net218),
    .X(caravel_wb_adr_o[1]));
 sky130_fd_sc_hd__clkbuf_2 output219 (.A(net219),
    .X(caravel_wb_adr_o[20]));
 sky130_fd_sc_hd__clkbuf_2 output220 (.A(net220),
    .X(caravel_wb_adr_o[21]));
 sky130_fd_sc_hd__clkbuf_2 output221 (.A(net221),
    .X(caravel_wb_adr_o[22]));
 sky130_fd_sc_hd__clkbuf_2 output222 (.A(net222),
    .X(caravel_wb_adr_o[23]));
 sky130_fd_sc_hd__clkbuf_2 output223 (.A(net223),
    .X(caravel_wb_adr_o[24]));
 sky130_fd_sc_hd__clkbuf_2 output224 (.A(net224),
    .X(caravel_wb_adr_o[25]));
 sky130_fd_sc_hd__clkbuf_2 output225 (.A(net225),
    .X(caravel_wb_adr_o[26]));
 sky130_fd_sc_hd__clkbuf_2 output226 (.A(net226),
    .X(caravel_wb_adr_o[27]));
 sky130_fd_sc_hd__clkbuf_2 output227 (.A(net227),
    .X(caravel_wb_adr_o[2]));
 sky130_fd_sc_hd__clkbuf_2 output228 (.A(net228),
    .X(caravel_wb_adr_o[3]));
 sky130_fd_sc_hd__clkbuf_2 output229 (.A(net229),
    .X(caravel_wb_adr_o[4]));
 sky130_fd_sc_hd__clkbuf_2 output230 (.A(net230),
    .X(caravel_wb_adr_o[5]));
 sky130_fd_sc_hd__clkbuf_2 output231 (.A(net231),
    .X(caravel_wb_adr_o[6]));
 sky130_fd_sc_hd__clkbuf_2 output232 (.A(net232),
    .X(caravel_wb_adr_o[7]));
 sky130_fd_sc_hd__clkbuf_2 output233 (.A(net233),
    .X(caravel_wb_adr_o[8]));
 sky130_fd_sc_hd__clkbuf_2 output234 (.A(net234),
    .X(caravel_wb_adr_o[9]));
 sky130_fd_sc_hd__clkbuf_2 output235 (.A(net414),
    .X(caravel_wb_cyc_o));
 sky130_fd_sc_hd__clkbuf_2 output236 (.A(net236),
    .X(caravel_wb_data_o[0]));
 sky130_fd_sc_hd__clkbuf_2 output237 (.A(net237),
    .X(caravel_wb_data_o[10]));
 sky130_fd_sc_hd__clkbuf_2 output238 (.A(net238),
    .X(caravel_wb_data_o[11]));
 sky130_fd_sc_hd__clkbuf_2 output239 (.A(net239),
    .X(caravel_wb_data_o[12]));
 sky130_fd_sc_hd__clkbuf_2 output240 (.A(net240),
    .X(caravel_wb_data_o[13]));
 sky130_fd_sc_hd__clkbuf_2 output241 (.A(net241),
    .X(caravel_wb_data_o[14]));
 sky130_fd_sc_hd__clkbuf_2 output242 (.A(net242),
    .X(caravel_wb_data_o[15]));
 sky130_fd_sc_hd__clkbuf_2 output243 (.A(net243),
    .X(caravel_wb_data_o[16]));
 sky130_fd_sc_hd__clkbuf_2 output244 (.A(net244),
    .X(caravel_wb_data_o[17]));
 sky130_fd_sc_hd__clkbuf_2 output245 (.A(net245),
    .X(caravel_wb_data_o[18]));
 sky130_fd_sc_hd__clkbuf_2 output246 (.A(net246),
    .X(caravel_wb_data_o[19]));
 sky130_fd_sc_hd__clkbuf_2 output247 (.A(net247),
    .X(caravel_wb_data_o[1]));
 sky130_fd_sc_hd__clkbuf_2 output248 (.A(net248),
    .X(caravel_wb_data_o[20]));
 sky130_fd_sc_hd__clkbuf_2 output249 (.A(net249),
    .X(caravel_wb_data_o[21]));
 sky130_fd_sc_hd__clkbuf_2 output250 (.A(net250),
    .X(caravel_wb_data_o[22]));
 sky130_fd_sc_hd__clkbuf_2 output251 (.A(net251),
    .X(caravel_wb_data_o[23]));
 sky130_fd_sc_hd__clkbuf_2 output252 (.A(net252),
    .X(caravel_wb_data_o[24]));
 sky130_fd_sc_hd__clkbuf_2 output253 (.A(net253),
    .X(caravel_wb_data_o[25]));
 sky130_fd_sc_hd__clkbuf_2 output254 (.A(net254),
    .X(caravel_wb_data_o[26]));
 sky130_fd_sc_hd__clkbuf_2 output255 (.A(net255),
    .X(caravel_wb_data_o[27]));
 sky130_fd_sc_hd__clkbuf_2 output256 (.A(net256),
    .X(caravel_wb_data_o[28]));
 sky130_fd_sc_hd__clkbuf_2 output257 (.A(net257),
    .X(caravel_wb_data_o[29]));
 sky130_fd_sc_hd__clkbuf_2 output258 (.A(net258),
    .X(caravel_wb_data_o[2]));
 sky130_fd_sc_hd__clkbuf_2 output259 (.A(net259),
    .X(caravel_wb_data_o[30]));
 sky130_fd_sc_hd__clkbuf_2 output260 (.A(net260),
    .X(caravel_wb_data_o[31]));
 sky130_fd_sc_hd__clkbuf_2 output261 (.A(net261),
    .X(caravel_wb_data_o[3]));
 sky130_fd_sc_hd__clkbuf_2 output262 (.A(net262),
    .X(caravel_wb_data_o[4]));
 sky130_fd_sc_hd__clkbuf_2 output263 (.A(net263),
    .X(caravel_wb_data_o[5]));
 sky130_fd_sc_hd__clkbuf_2 output264 (.A(net264),
    .X(caravel_wb_data_o[6]));
 sky130_fd_sc_hd__clkbuf_2 output265 (.A(net265),
    .X(caravel_wb_data_o[7]));
 sky130_fd_sc_hd__clkbuf_2 output266 (.A(net266),
    .X(caravel_wb_data_o[8]));
 sky130_fd_sc_hd__clkbuf_2 output267 (.A(net267),
    .X(caravel_wb_data_o[9]));
 sky130_fd_sc_hd__clkbuf_2 output268 (.A(net268),
    .X(caravel_wb_sel_o[0]));
 sky130_fd_sc_hd__clkbuf_2 output269 (.A(net269),
    .X(caravel_wb_sel_o[1]));
 sky130_fd_sc_hd__clkbuf_2 output270 (.A(net270),
    .X(caravel_wb_sel_o[2]));
 sky130_fd_sc_hd__clkbuf_2 output271 (.A(net271),
    .X(caravel_wb_sel_o[3]));
 sky130_fd_sc_hd__clkbuf_2 output272 (.A(net272),
    .X(caravel_wb_stb_o));
 sky130_fd_sc_hd__clkbuf_2 output273 (.A(net273),
    .X(caravel_wb_we_o));
 sky130_fd_sc_hd__buf_12 output274 (.A(net274),
    .X(la_data_out[0]));
 sky130_fd_sc_hd__buf_12 output275 (.A(net275),
    .X(la_data_out[10]));
 sky130_fd_sc_hd__buf_12 output276 (.A(net276),
    .X(la_data_out[11]));
 sky130_fd_sc_hd__buf_12 output277 (.A(net277),
    .X(la_data_out[12]));
 sky130_fd_sc_hd__buf_12 output278 (.A(net278),
    .X(la_data_out[13]));
 sky130_fd_sc_hd__buf_12 output279 (.A(net279),
    .X(la_data_out[14]));
 sky130_fd_sc_hd__buf_12 output280 (.A(net280),
    .X(la_data_out[15]));
 sky130_fd_sc_hd__buf_12 output281 (.A(net281),
    .X(la_data_out[16]));
 sky130_fd_sc_hd__buf_12 output282 (.A(net282),
    .X(la_data_out[17]));
 sky130_fd_sc_hd__buf_12 output283 (.A(net283),
    .X(la_data_out[18]));
 sky130_fd_sc_hd__buf_12 output284 (.A(net284),
    .X(la_data_out[19]));
 sky130_fd_sc_hd__buf_12 output285 (.A(net285),
    .X(la_data_out[1]));
 sky130_fd_sc_hd__buf_12 output286 (.A(net286),
    .X(la_data_out[20]));
 sky130_fd_sc_hd__buf_12 output287 (.A(net287),
    .X(la_data_out[21]));
 sky130_fd_sc_hd__buf_12 output288 (.A(net288),
    .X(la_data_out[22]));
 sky130_fd_sc_hd__buf_12 output289 (.A(net289),
    .X(la_data_out[23]));
 sky130_fd_sc_hd__buf_12 output290 (.A(net290),
    .X(la_data_out[24]));
 sky130_fd_sc_hd__buf_12 output291 (.A(net291),
    .X(la_data_out[25]));
 sky130_fd_sc_hd__buf_12 output292 (.A(net292),
    .X(la_data_out[26]));
 sky130_fd_sc_hd__buf_12 output293 (.A(net293),
    .X(la_data_out[27]));
 sky130_fd_sc_hd__buf_12 output294 (.A(net294),
    .X(la_data_out[28]));
 sky130_fd_sc_hd__buf_12 output295 (.A(net295),
    .X(la_data_out[29]));
 sky130_fd_sc_hd__buf_12 output296 (.A(net296),
    .X(la_data_out[2]));
 sky130_fd_sc_hd__buf_12 output297 (.A(net297),
    .X(la_data_out[30]));
 sky130_fd_sc_hd__buf_12 output298 (.A(net298),
    .X(la_data_out[31]));
 sky130_fd_sc_hd__buf_12 output299 (.A(net299),
    .X(la_data_out[32]));
 sky130_fd_sc_hd__buf_12 output300 (.A(net300),
    .X(la_data_out[33]));
 sky130_fd_sc_hd__buf_12 output301 (.A(net301),
    .X(la_data_out[34]));
 sky130_fd_sc_hd__buf_12 output302 (.A(net302),
    .X(la_data_out[35]));
 sky130_fd_sc_hd__buf_12 output303 (.A(net303),
    .X(la_data_out[36]));
 sky130_fd_sc_hd__buf_12 output304 (.A(net304),
    .X(la_data_out[37]));
 sky130_fd_sc_hd__buf_12 output305 (.A(net305),
    .X(la_data_out[38]));
 sky130_fd_sc_hd__buf_12 output306 (.A(net306),
    .X(la_data_out[39]));
 sky130_fd_sc_hd__buf_12 output307 (.A(net307),
    .X(la_data_out[3]));
 sky130_fd_sc_hd__buf_12 output308 (.A(net308),
    .X(la_data_out[40]));
 sky130_fd_sc_hd__buf_12 output309 (.A(net309),
    .X(la_data_out[41]));
 sky130_fd_sc_hd__buf_12 output310 (.A(net310),
    .X(la_data_out[42]));
 sky130_fd_sc_hd__buf_12 output311 (.A(net311),
    .X(la_data_out[43]));
 sky130_fd_sc_hd__buf_12 output312 (.A(net312),
    .X(la_data_out[44]));
 sky130_fd_sc_hd__buf_12 output313 (.A(net313),
    .X(la_data_out[45]));
 sky130_fd_sc_hd__buf_12 output314 (.A(net314),
    .X(la_data_out[46]));
 sky130_fd_sc_hd__buf_12 output315 (.A(net315),
    .X(la_data_out[47]));
 sky130_fd_sc_hd__buf_12 output316 (.A(net316),
    .X(la_data_out[48]));
 sky130_fd_sc_hd__buf_12 output317 (.A(net317),
    .X(la_data_out[49]));
 sky130_fd_sc_hd__buf_12 output318 (.A(net318),
    .X(la_data_out[4]));
 sky130_fd_sc_hd__buf_12 output319 (.A(net319),
    .X(la_data_out[50]));
 sky130_fd_sc_hd__buf_12 output320 (.A(net320),
    .X(la_data_out[51]));
 sky130_fd_sc_hd__buf_12 output321 (.A(net321),
    .X(la_data_out[52]));
 sky130_fd_sc_hd__buf_12 output322 (.A(net322),
    .X(la_data_out[53]));
 sky130_fd_sc_hd__buf_12 output323 (.A(net323),
    .X(la_data_out[54]));
 sky130_fd_sc_hd__buf_12 output324 (.A(net324),
    .X(la_data_out[55]));
 sky130_fd_sc_hd__buf_12 output325 (.A(net325),
    .X(la_data_out[56]));
 sky130_fd_sc_hd__buf_12 output326 (.A(net326),
    .X(la_data_out[57]));
 sky130_fd_sc_hd__buf_12 output327 (.A(net327),
    .X(la_data_out[58]));
 sky130_fd_sc_hd__buf_12 output328 (.A(net328),
    .X(la_data_out[59]));
 sky130_fd_sc_hd__buf_12 output329 (.A(net329),
    .X(la_data_out[5]));
 sky130_fd_sc_hd__buf_12 output330 (.A(net330),
    .X(la_data_out[60]));
 sky130_fd_sc_hd__buf_12 output331 (.A(net331),
    .X(la_data_out[61]));
 sky130_fd_sc_hd__buf_12 output332 (.A(net332),
    .X(la_data_out[62]));
 sky130_fd_sc_hd__buf_12 output333 (.A(net333),
    .X(la_data_out[63]));
 sky130_fd_sc_hd__buf_12 output334 (.A(net334),
    .X(la_data_out[64]));
 sky130_fd_sc_hd__buf_12 output335 (.A(net335),
    .X(la_data_out[65]));
 sky130_fd_sc_hd__buf_12 output336 (.A(net336),
    .X(la_data_out[66]));
 sky130_fd_sc_hd__buf_12 output337 (.A(net337),
    .X(la_data_out[67]));
 sky130_fd_sc_hd__buf_12 output338 (.A(net338),
    .X(la_data_out[68]));
 sky130_fd_sc_hd__buf_12 output339 (.A(net339),
    .X(la_data_out[69]));
 sky130_fd_sc_hd__buf_12 output340 (.A(net340),
    .X(la_data_out[6]));
 sky130_fd_sc_hd__buf_12 output341 (.A(net341),
    .X(la_data_out[70]));
 sky130_fd_sc_hd__buf_12 output342 (.A(net342),
    .X(la_data_out[71]));
 sky130_fd_sc_hd__buf_12 output343 (.A(net343),
    .X(la_data_out[72]));
 sky130_fd_sc_hd__buf_12 output344 (.A(net344),
    .X(la_data_out[73]));
 sky130_fd_sc_hd__buf_12 output345 (.A(net345),
    .X(la_data_out[74]));
 sky130_fd_sc_hd__buf_12 output346 (.A(net346),
    .X(la_data_out[75]));
 sky130_fd_sc_hd__buf_12 output347 (.A(net347),
    .X(la_data_out[76]));
 sky130_fd_sc_hd__buf_12 output348 (.A(net348),
    .X(la_data_out[77]));
 sky130_fd_sc_hd__buf_12 output349 (.A(net349),
    .X(la_data_out[78]));
 sky130_fd_sc_hd__buf_12 output350 (.A(net350),
    .X(la_data_out[79]));
 sky130_fd_sc_hd__buf_12 output351 (.A(net351),
    .X(la_data_out[7]));
 sky130_fd_sc_hd__buf_12 output352 (.A(net352),
    .X(la_data_out[80]));
 sky130_fd_sc_hd__buf_12 output353 (.A(net353),
    .X(la_data_out[81]));
 sky130_fd_sc_hd__buf_12 output354 (.A(net354),
    .X(la_data_out[82]));
 sky130_fd_sc_hd__buf_12 output355 (.A(net355),
    .X(la_data_out[83]));
 sky130_fd_sc_hd__buf_12 output356 (.A(net356),
    .X(la_data_out[84]));
 sky130_fd_sc_hd__buf_12 output357 (.A(net357),
    .X(la_data_out[85]));
 sky130_fd_sc_hd__buf_12 output358 (.A(net358),
    .X(la_data_out[86]));
 sky130_fd_sc_hd__buf_12 output359 (.A(net359),
    .X(la_data_out[87]));
 sky130_fd_sc_hd__buf_12 output360 (.A(net360),
    .X(la_data_out[88]));
 sky130_fd_sc_hd__buf_12 output361 (.A(net361),
    .X(la_data_out[89]));
 sky130_fd_sc_hd__buf_12 output362 (.A(net362),
    .X(la_data_out[8]));
 sky130_fd_sc_hd__buf_12 output363 (.A(net363),
    .X(la_data_out[90]));
 sky130_fd_sc_hd__buf_12 output364 (.A(net364),
    .X(la_data_out[91]));
 sky130_fd_sc_hd__buf_12 output365 (.A(net365),
    .X(la_data_out[92]));
 sky130_fd_sc_hd__buf_12 output366 (.A(net366),
    .X(la_data_out[93]));
 sky130_fd_sc_hd__buf_12 output367 (.A(net367),
    .X(la_data_out[94]));
 sky130_fd_sc_hd__buf_12 output368 (.A(net368),
    .X(la_data_out[95]));
 sky130_fd_sc_hd__buf_12 output369 (.A(net369),
    .X(la_data_out[96]));
 sky130_fd_sc_hd__buf_12 output370 (.A(net370),
    .X(la_data_out[97]));
 sky130_fd_sc_hd__buf_12 output371 (.A(net371),
    .X(la_data_out[9]));
 sky130_fd_sc_hd__buf_12 output372 (.A(net372),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__clkbuf_2 output373 (.A(net373),
    .X(wbs_data_o[0]));
 sky130_fd_sc_hd__clkbuf_2 output374 (.A(net374),
    .X(wbs_data_o[10]));
 sky130_fd_sc_hd__clkbuf_2 output375 (.A(net375),
    .X(wbs_data_o[11]));
 sky130_fd_sc_hd__clkbuf_2 output376 (.A(net376),
    .X(wbs_data_o[12]));
 sky130_fd_sc_hd__clkbuf_2 output377 (.A(net377),
    .X(wbs_data_o[13]));
 sky130_fd_sc_hd__clkbuf_2 output378 (.A(net378),
    .X(wbs_data_o[14]));
 sky130_fd_sc_hd__clkbuf_2 output379 (.A(net379),
    .X(wbs_data_o[15]));
 sky130_fd_sc_hd__clkbuf_2 output380 (.A(net380),
    .X(wbs_data_o[16]));
 sky130_fd_sc_hd__clkbuf_2 output381 (.A(net381),
    .X(wbs_data_o[17]));
 sky130_fd_sc_hd__clkbuf_2 output382 (.A(net382),
    .X(wbs_data_o[18]));
 sky130_fd_sc_hd__clkbuf_2 output383 (.A(net383),
    .X(wbs_data_o[19]));
 sky130_fd_sc_hd__clkbuf_2 output384 (.A(net384),
    .X(wbs_data_o[1]));
 sky130_fd_sc_hd__clkbuf_2 output385 (.A(net385),
    .X(wbs_data_o[20]));
 sky130_fd_sc_hd__clkbuf_2 output386 (.A(net386),
    .X(wbs_data_o[21]));
 sky130_fd_sc_hd__clkbuf_2 output387 (.A(net387),
    .X(wbs_data_o[22]));
 sky130_fd_sc_hd__clkbuf_2 output388 (.A(net388),
    .X(wbs_data_o[23]));
 sky130_fd_sc_hd__clkbuf_2 output389 (.A(net389),
    .X(wbs_data_o[24]));
 sky130_fd_sc_hd__clkbuf_2 output390 (.A(net390),
    .X(wbs_data_o[25]));
 sky130_fd_sc_hd__clkbuf_2 output391 (.A(net391),
    .X(wbs_data_o[26]));
 sky130_fd_sc_hd__clkbuf_2 output392 (.A(net392),
    .X(wbs_data_o[27]));
 sky130_fd_sc_hd__clkbuf_2 output393 (.A(net393),
    .X(wbs_data_o[28]));
 sky130_fd_sc_hd__clkbuf_2 output394 (.A(net394),
    .X(wbs_data_o[29]));
 sky130_fd_sc_hd__clkbuf_2 output395 (.A(net395),
    .X(wbs_data_o[2]));
 sky130_fd_sc_hd__clkbuf_2 output396 (.A(net396),
    .X(wbs_data_o[30]));
 sky130_fd_sc_hd__clkbuf_2 output397 (.A(net397),
    .X(wbs_data_o[31]));
 sky130_fd_sc_hd__clkbuf_2 output398 (.A(net398),
    .X(wbs_data_o[3]));
 sky130_fd_sc_hd__clkbuf_2 output399 (.A(net399),
    .X(wbs_data_o[4]));
 sky130_fd_sc_hd__clkbuf_2 output400 (.A(net400),
    .X(wbs_data_o[5]));
 sky130_fd_sc_hd__clkbuf_2 output401 (.A(net401),
    .X(wbs_data_o[6]));
 sky130_fd_sc_hd__clkbuf_2 output402 (.A(net402),
    .X(wbs_data_o[7]));
 sky130_fd_sc_hd__clkbuf_2 output403 (.A(net403),
    .X(wbs_data_o[8]));
 sky130_fd_sc_hd__clkbuf_2 output404 (.A(net404),
    .X(wbs_data_o[9]));
 sky130_fd_sc_hd__buf_4 split1 (.A(net486),
    .X(net1282));
 sky130_fd_sc_hd__buf_4 split2 (.A(net503),
    .X(net1283));
 sky130_fd_sc_hd__buf_2 split3 (.A(net442),
    .X(net1284));
 sky130_fd_sc_hd__buf_2 split4 (.A(net502),
    .X(net1285));
 sky130_fd_sc_hd__clkbuf_2 split5 (.A(net484),
    .X(net1286));
 assign caravel_irq[0] = net651;
 assign caravel_irq[1] = net652;
 assign caravel_irq[2] = net653;
 assign caravel_irq[3] = net654;
 assign core0Index[0] = net655;
 assign core0Index[1] = net656;
 assign core0Index[2] = net657;
 assign core0Index[3] = net658;
 assign core0Index[4] = net659;
 assign core0Index[5] = net660;
 assign core0Index[6] = net661;
 assign core0Index[7] = net662;
 assign core1Index[0] = net722;
 assign core1Index[1] = net663;
 assign core1Index[2] = net664;
 assign core1Index[3] = net665;
 assign core1Index[4] = net666;
 assign core1Index[5] = net667;
 assign core1Index[6] = net668;
 assign core1Index[7] = net669;
 assign la_data_out[100] = net672;
 assign la_data_out[101] = net673;
 assign la_data_out[102] = net674;
 assign la_data_out[103] = net675;
 assign la_data_out[104] = net676;
 assign la_data_out[105] = net677;
 assign la_data_out[106] = net678;
 assign la_data_out[107] = net679;
 assign la_data_out[108] = net680;
 assign la_data_out[109] = net681;
 assign la_data_out[110] = net682;
 assign la_data_out[111] = net683;
 assign la_data_out[112] = net684;
 assign la_data_out[113] = net685;
 assign la_data_out[114] = net686;
 assign la_data_out[115] = net687;
 assign la_data_out[116] = net688;
 assign la_data_out[117] = net689;
 assign la_data_out[118] = net690;
 assign la_data_out[119] = net691;
 assign la_data_out[120] = net692;
 assign la_data_out[121] = net693;
 assign la_data_out[122] = net694;
 assign la_data_out[123] = net695;
 assign la_data_out[124] = net696;
 assign la_data_out[125] = net697;
 assign la_data_out[126] = net698;
 assign la_data_out[127] = net699;
 assign la_data_out[98] = net670;
 assign la_data_out[99] = net671;
 assign manufacturerID[0] = net700;
 assign manufacturerID[10] = net710;
 assign manufacturerID[1] = net701;
 assign manufacturerID[2] = net702;
 assign manufacturerID[3] = net703;
 assign manufacturerID[4] = net704;
 assign manufacturerID[5] = net705;
 assign manufacturerID[6] = net706;
 assign manufacturerID[7] = net707;
 assign manufacturerID[8] = net708;
 assign manufacturerID[9] = net709;
 assign partID[0] = net723;
 assign partID[10] = net728;
 assign partID[11] = net729;
 assign partID[12] = net716;
 assign partID[13] = net717;
 assign partID[14] = net730;
 assign partID[15] = net731;
 assign partID[1] = net711;
 assign partID[2] = net724;
 assign partID[3] = net712;
 assign partID[4] = net725;
 assign partID[5] = net713;
 assign partID[6] = net726;
 assign partID[7] = net714;
 assign partID[8] = net727;
 assign partID[9] = net715;
 assign versionID[0] = net718;
 assign versionID[1] = net719;
 assign versionID[2] = net720;
 assign versionID[3] = net721;
endmodule

