* NGSPICE file created from CaravelHost.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

.subckt CaravelHost caravel_irq[0] caravel_irq[1] caravel_irq[2] caravel_irq[3] caravel_uart_rx
+ caravel_uart_tx caravel_wb_ack_i caravel_wb_adr_o[0] caravel_wb_adr_o[10] caravel_wb_adr_o[11]
+ caravel_wb_adr_o[12] caravel_wb_adr_o[13] caravel_wb_adr_o[14] caravel_wb_adr_o[15]
+ caravel_wb_adr_o[16] caravel_wb_adr_o[17] caravel_wb_adr_o[18] caravel_wb_adr_o[19]
+ caravel_wb_adr_o[1] caravel_wb_adr_o[20] caravel_wb_adr_o[21] caravel_wb_adr_o[22]
+ caravel_wb_adr_o[23] caravel_wb_adr_o[24] caravel_wb_adr_o[25] caravel_wb_adr_o[26]
+ caravel_wb_adr_o[27] caravel_wb_adr_o[2] caravel_wb_adr_o[3] caravel_wb_adr_o[4]
+ caravel_wb_adr_o[5] caravel_wb_adr_o[6] caravel_wb_adr_o[7] caravel_wb_adr_o[8]
+ caravel_wb_adr_o[9] caravel_wb_cyc_o caravel_wb_data_i[0] caravel_wb_data_i[10]
+ caravel_wb_data_i[11] caravel_wb_data_i[12] caravel_wb_data_i[13] caravel_wb_data_i[14]
+ caravel_wb_data_i[15] caravel_wb_data_i[16] caravel_wb_data_i[17] caravel_wb_data_i[18]
+ caravel_wb_data_i[19] caravel_wb_data_i[1] caravel_wb_data_i[20] caravel_wb_data_i[21]
+ caravel_wb_data_i[22] caravel_wb_data_i[23] caravel_wb_data_i[24] caravel_wb_data_i[25]
+ caravel_wb_data_i[26] caravel_wb_data_i[27] caravel_wb_data_i[28] caravel_wb_data_i[29]
+ caravel_wb_data_i[2] caravel_wb_data_i[30] caravel_wb_data_i[31] caravel_wb_data_i[3]
+ caravel_wb_data_i[4] caravel_wb_data_i[5] caravel_wb_data_i[6] caravel_wb_data_i[7]
+ caravel_wb_data_i[8] caravel_wb_data_i[9] caravel_wb_data_o[0] caravel_wb_data_o[10]
+ caravel_wb_data_o[11] caravel_wb_data_o[12] caravel_wb_data_o[13] caravel_wb_data_o[14]
+ caravel_wb_data_o[15] caravel_wb_data_o[16] caravel_wb_data_o[17] caravel_wb_data_o[18]
+ caravel_wb_data_o[19] caravel_wb_data_o[1] caravel_wb_data_o[20] caravel_wb_data_o[21]
+ caravel_wb_data_o[22] caravel_wb_data_o[23] caravel_wb_data_o[24] caravel_wb_data_o[25]
+ caravel_wb_data_o[26] caravel_wb_data_o[27] caravel_wb_data_o[28] caravel_wb_data_o[29]
+ caravel_wb_data_o[2] caravel_wb_data_o[30] caravel_wb_data_o[31] caravel_wb_data_o[3]
+ caravel_wb_data_o[4] caravel_wb_data_o[5] caravel_wb_data_o[6] caravel_wb_data_o[7]
+ caravel_wb_data_o[8] caravel_wb_data_o[9] caravel_wb_error_i caravel_wb_sel_o[0]
+ caravel_wb_sel_o[1] caravel_wb_sel_o[2] caravel_wb_sel_o[3] caravel_wb_stall_i caravel_wb_stb_o
+ caravel_wb_we_o core0Index[0] core0Index[1] core0Index[2] core0Index[3] core0Index[4]
+ core0Index[5] core0Index[6] core0Index[7] core1Index[0] core1Index[1] core1Index[2]
+ core1Index[3] core1Index[4] core1Index[5] core1Index[6] core1Index[7] manufacturerID[0]
+ manufacturerID[10] manufacturerID[1] manufacturerID[2] manufacturerID[3] manufacturerID[4]
+ manufacturerID[5] manufacturerID[6] manufacturerID[7] manufacturerID[8] manufacturerID[9]
+ partID[0] partID[10] partID[11] partID[12] partID[13] partID[14] partID[15] partID[1]
+ partID[2] partID[3] partID[4] partID[5] partID[6] partID[7] partID[8] partID[9]
+ vccd1 versionID[0] versionID[1] versionID[2] versionID[3] vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_data_i[0] wbs_data_i[10] wbs_data_i[11] wbs_data_i[12]
+ wbs_data_i[13] wbs_data_i[14] wbs_data_i[15] wbs_data_i[16] wbs_data_i[17] wbs_data_i[18]
+ wbs_data_i[19] wbs_data_i[1] wbs_data_i[20] wbs_data_i[21] wbs_data_i[22] wbs_data_i[23]
+ wbs_data_i[24] wbs_data_i[25] wbs_data_i[26] wbs_data_i[27] wbs_data_i[28] wbs_data_i[29]
+ wbs_data_i[2] wbs_data_i[30] wbs_data_i[31] wbs_data_i[3] wbs_data_i[4] wbs_data_i[5]
+ wbs_data_i[6] wbs_data_i[7] wbs_data_i[8] wbs_data_i[9] wbs_data_o[0] wbs_data_o[10]
+ wbs_data_o[11] wbs_data_o[12] wbs_data_o[13] wbs_data_o[14] wbs_data_o[15] wbs_data_o[16]
+ wbs_data_o[17] wbs_data_o[18] wbs_data_o[19] wbs_data_o[1] wbs_data_o[20] wbs_data_o[21]
+ wbs_data_o[22] wbs_data_o[23] wbs_data_o[24] wbs_data_o[25] wbs_data_o[26] wbs_data_o[27]
+ wbs_data_o[28] wbs_data_o[29] wbs_data_o[2] wbs_data_o[30] wbs_data_o[31] wbs_data_o[3]
+ wbs_data_o[4] wbs_data_o[5] wbs_data_o[6] wbs_data_o[7] wbs_data_o[8] wbs_data_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7963_ _7963_/CLK _7963_/D vssd1 vssd1 vccd1 vccd1 _7963_/Q sky130_fd_sc_hd__dfxtp_1
X_6914_ _6914_/A vssd1 vssd1 vccd1 vccd1 _8113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7894_ _8520_/CLK _7894_/D vssd1 vssd1 vccd1 vccd1 _7894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8570__217 vssd1 vssd1 vccd1 vccd1 _8570__217/HI core0Index[4] sky130_fd_sc_hd__conb_1
X_6845_ _6838_/X _6839_/Y _6842_/Y _6843_/Y _6844_/X vssd1 vssd1 vccd1 vccd1 _6845_/X
+ sky130_fd_sc_hd__o2111a_1
X_3988_ _3831_/X _8450_/Q _3996_/S vssd1 vssd1 vccd1 vccd1 _3989_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8515_ _8515_/CLK _8515_/D vssd1 vssd1 vccd1 vccd1 _8515_/Q sky130_fd_sc_hd__dfxtp_1
X_5727_ _7920_/Q _5593_/X _5731_/S vssd1 vssd1 vccd1 vccd1 _5728_/A sky130_fd_sc_hd__mux2_1
X_8446_ _8446_/CLK _8446_/D vssd1 vssd1 vccd1 vccd1 _8446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5658_ _5658_/A vssd1 vssd1 vccd1 vccd1 _7951_/D sky130_fd_sc_hd__clkbuf_1
X_8377_ _8377_/CLK _8377_/D vssd1 vssd1 vccd1 vccd1 _8377_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3456_ _7083_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3456_/X sky130_fd_sc_hd__clkbuf_16
X_5589_ _5589_/A vssd1 vssd1 vccd1 vccd1 _7986_/D sky130_fd_sc_hd__clkbuf_1
X_4609_ _4609_/A vssd1 vssd1 vccd1 vccd1 _8195_/D sky130_fd_sc_hd__clkbuf_1
X_6947__414 _6948__415/A vssd1 vssd1 vccd1 vccd1 _8138_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3773_ clkbuf_0__3773_/X vssd1 vssd1 vccd1 vccd1 _7657__35/A sky130_fd_sc_hd__clkbuf_4
X_7328_ _7336_/A _7328_/B vssd1 vssd1 vccd1 vccd1 _8350_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7259_ _8352_/Q vssd1 vssd1 vccd1 vccd1 _7259_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6887__383 _6887__383/A vssd1 vssd1 vccd1 vccd1 _8097_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _4975_/S vssd1 vssd1 vccd1 vccd1 _4969_/S sky130_fd_sc_hd__buf_2
XFILLER_51_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4891_ _4901_/S vssd1 vssd1 vccd1 vccd1 _4909_/S sky130_fd_sc_hd__clkbuf_4
X_3911_ _8488_/Q vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__buf_4
XFILLER_20_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3842_ _5345_/A _8114_/Q vssd1 vssd1 vccd1 vccd1 _5034_/D sky130_fd_sc_hd__nand2_1
X_5512_ _8040_/Q _4292_/A _5516_/S vssd1 vssd1 vccd1 vccd1 _5513_/A sky130_fd_sc_hd__mux2_1
X_8300_ _8300_/CLK _8300_/D vssd1 vssd1 vccd1 vccd1 _8300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3273_ clkbuf_0__3273_/X vssd1 vssd1 vccd1 vccd1 _6643__303/A sky130_fd_sc_hd__clkbuf_4
X_6751__347 _6754__350/A vssd1 vssd1 vccd1 vccd1 _8057_/CLK sky130_fd_sc_hd__inv_2
X_6492_ _6000_/A _7888_/Q _6498_/S vssd1 vssd1 vccd1 vccd1 _6493_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3310_ _6731_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3310_/X sky130_fd_sc_hd__clkbuf_16
X_5443_ _5443_/A vssd1 vssd1 vccd1 vccd1 _8074_/D sky130_fd_sc_hd__clkbuf_1
X_8231_ _8231_/CLK _8231_/D vssd1 vssd1 vccd1 vccd1 _8231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7487__20 _7487__20/A vssd1 vssd1 vccd1 vccd1 _8452_/CLK sky130_fd_sc_hd__inv_2
X_5374_ _8109_/Q vssd1 vssd1 vccd1 vccd1 _5566_/A sky130_fd_sc_hd__buf_2
X_8162_ _8162_/CLK _8162_/D vssd1 vssd1 vccd1 vccd1 _8162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4325_ _4325_/A vssd1 vssd1 vccd1 vccd1 _8307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8093_ _8093_/CLK _8093_/D vssd1 vssd1 vccd1 vccd1 _8093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4256_ _4256_/A _4301_/B _4256_/C vssd1 vssd1 vccd1 vccd1 _5787_/B sky130_fd_sc_hd__nand3_4
X_4187_ _8491_/Q vssd1 vssd1 vccd1 vccd1 _4187_/X sky130_fd_sc_hd__buf_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7946_ _7946_/CLK _7946_/D vssd1 vssd1 vccd1 vccd1 _7946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7877_ _8345_/CLK _7877_/D vssd1 vssd1 vccd1 vccd1 _7877_/Q sky130_fd_sc_hd__dfxtp_1
X_6828_ _7576_/A _7576_/B _8544_/Q vssd1 vssd1 vccd1 vccd1 _6828_/X sky130_fd_sc_hd__a21bo_1
XFILLER_11_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6759_ _6759_/A vssd1 vssd1 vccd1 vccd1 _8062_/D sky130_fd_sc_hd__clkbuf_1
X_8429_ _8429_/CLK _8429_/D vssd1 vssd1 vccd1 vccd1 _8429_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3439_ _6994_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3439_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_78_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7181__99 _7181__99/A vssd1 vssd1 vccd1 vccd1 _8326_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4031_/X _8404_/Q _4112_/S vssd1 vssd1 vccd1 vccd1 _4111_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _5169_/A _5090_/B vssd1 vssd1 vccd1 vccd1 _5090_/X sky130_fd_sc_hd__and2_1
XFILLER_69_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4041_ _4005_/X _8434_/Q _4049_/S vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5992_ _5992_/A vssd1 vssd1 vccd1 vccd1 _5992_/X sky130_fd_sc_hd__clkbuf_1
X_7800_ _8531_/CLK _7800_/D vssd1 vssd1 vccd1 vccd1 _7800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7731_ _7731_/A vssd1 vssd1 vccd1 vccd1 _7731_/X sky130_fd_sc_hd__clkbuf_2
X_4943_ _4943_/A _4943_/B vssd1 vssd1 vccd1 vccd1 _8174_/D sky130_fd_sc_hd__nor2_1
X_4874_ _8230_/Q _4775_/X _4777_/X _8214_/Q _4654_/A vssd1 vssd1 vccd1 vccd1 _4874_/X
+ sky130_fd_sc_hd__o221a_1
X_6613_ _8182_/Q _8167_/D vssd1 vssd1 vccd1 vccd1 _6614_/A sky130_fd_sc_hd__and2_1
X_7593_ _6812_/B _7588_/X _7547_/X _6793_/B vssd1 vssd1 vccd1 vccd1 _7594_/B sky130_fd_sc_hd__o22a_1
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3256_ clkbuf_0__3256_/X vssd1 vssd1 vccd1 vccd1 _6632_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6475_ _6475_/A vssd1 vssd1 vccd1 vccd1 _7880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8214_ _8214_/CLK _8214_/D vssd1 vssd1 vccd1 vccd1 _8214_/Q sky130_fd_sc_hd__dfxtp_1
X_5426_ _5387_/X _8082_/Q _5426_/S vssd1 vssd1 vccd1 vccd1 _5427_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8145_ _8145_/CLK _8145_/D vssd1 vssd1 vccd1 vccd1 _8145_/Q sky130_fd_sc_hd__dfxtp_1
X_5357_ _5061_/X _5348_/X _5356_/Y _5339_/X vssd1 vssd1 vccd1 vccd1 _8115_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8076_ _8076_/CLK _8076_/D vssd1 vssd1 vccd1 vccd1 _8076_/Q sky130_fd_sc_hd__dfxtp_1
X_5288_ _8497_/Q _5232_/A _5214_/X _8513_/Q _5100_/A vssd1 vssd1 vccd1 vccd1 _5288_/X
+ sky130_fd_sc_hd__o221a_1
X_7044__489 _7045__490/A vssd1 vssd1 vccd1 vccd1 _8216_/CLK sky130_fd_sc_hd__inv_2
X_4308_ _4283_/X _8314_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4309_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_4 _7821_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4239_ _4254_/S vssd1 vssd1 vccd1 vccd1 _4248_/S sky130_fd_sc_hd__buf_2
X_7027_ _7058_/A vssd1 vssd1 vccd1 vccd1 _7027_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3086_ _6291_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3086_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3472_ clkbuf_0__3472_/X vssd1 vssd1 vccd1 vccd1 _7164__85/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8576__223 vssd1 vssd1 vccd1 vccd1 _8576__223/HI core1Index[3] sky130_fd_sc_hd__conb_1
X_7929_ _7929_/CLK _7929_/D vssd1 vssd1 vccd1 vccd1 _7929_/Q sky130_fd_sc_hd__dfxtp_1
X_6990__448 _6992__450/A vssd1 vssd1 vccd1 vccd1 _8173_/CLK sky130_fd_sc_hd__inv_2
X_7448__163 _7450__165/A vssd1 vssd1 vccd1 vccd1 _8420_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7481__15 _7481__15/A vssd1 vssd1 vccd1 vccd1 _8447_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6301__203 _6303__205/A vssd1 vssd1 vccd1 vccd1 _7833_/CLK sky130_fd_sc_hd__inv_2
X_4590_ _4424_/X _8203_/Q _4596_/S vssd1 vssd1 vccd1 vccd1 _4591_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6260_ _7642_/A _7816_/Q _6264_/S vssd1 vssd1 vccd1 vccd1 _6261_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5211_ _8382_/Q _8390_/Q _5315_/S vssd1 vssd1 vccd1 vccd1 _5211_/X sky130_fd_sc_hd__mux2_2
X_6191_ _6202_/A vssd1 vssd1 vccd1 vccd1 _6191_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5142_ _8517_/Q _8070_/Q _8043_/Q _8501_/Q _5290_/S _5129_/X vssd1 vssd1 vccd1 vccd1
+ _5142_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5073_ _5354_/B _5069_/X _5235_/A vssd1 vssd1 vccd1 vccd1 _5073_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4024_ _4023_/X _8438_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4025_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5975_ _5975_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__and2_1
XFILLER_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3773_ _7652_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3773_/X sky130_fd_sc_hd__clkbuf_16
X_7714_ _8535_/Q _7701_/X _7713_/X _7704_/X vssd1 vssd1 vccd1 vccd1 _8535_/D sky130_fd_sc_hd__o211a_1
X_4926_ _8178_/Q _8187_/Q _4924_/X _4925_/Y vssd1 vssd1 vccd1 vccd1 _8178_/D sky130_fd_sc_hd__o211a_1
X_4857_ _6900_/B vssd1 vssd1 vccd1 vccd1 _4857_/X sky130_fd_sc_hd__clkbuf_2
X_7645_ _7645_/A vssd1 vssd1 vccd1 vccd1 _8494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7576_ _7576_/A _7576_/B vssd1 vssd1 vccd1 vccd1 _7576_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3308_ clkbuf_0__3308_/X vssd1 vssd1 vccd1 vccd1 _6737_/A sky130_fd_sc_hd__clkbuf_4
X_4788_ _7937_/Q _4784_/X _4785_/X _4787_/X vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__o22a_1
X_6527_ _6589_/A vssd1 vssd1 vccd1 vccd1 _6527_/X sky130_fd_sc_hd__buf_1
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6458_ _7875_/Q _6388_/X _6422_/X vssd1 vssd1 vccd1 vccd1 _7875_/D sky130_fd_sc_hd__a21o_1
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5409_ _5409_/A vssd1 vssd1 vccd1 vccd1 _8090_/D sky130_fd_sc_hd__clkbuf_1
X_6389_ _8546_/Q vssd1 vssd1 vccd1 vccd1 _7522_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8128_ _8128_/CLK _8128_/D vssd1 vssd1 vccd1 vccd1 _8128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8059_ _8059_/CLK _8059_/D vssd1 vssd1 vccd1 vccd1 _8059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3455_ clkbuf_0__3455_/X vssd1 vssd1 vccd1 vccd1 _7079__517/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7092__527 _7093__528/A vssd1 vssd1 vccd1 vccd1 _8254_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6927__401 _6930__404/A vssd1 vssd1 vccd1 vccd1 _8123_/CLK sky130_fd_sc_hd__inv_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5760_ _5760_/A vssd1 vssd1 vccd1 vccd1 _7906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _7936_/Q _5593_/X _5695_/S vssd1 vssd1 vccd1 vccd1 _5692_/A sky130_fd_sc_hd__mux2_1
X_4711_ _4424_/X _4629_/X _4710_/X _4690_/X vssd1 vssd1 vccd1 vccd1 _8185_/D sky130_fd_sc_hd__o211a_1
X_4642_ _4726_/A vssd1 vssd1 vccd1 vccd1 _4677_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ _3966_/X _8210_/Q _4577_/S vssd1 vssd1 vccd1 vccd1 _4574_/A sky130_fd_sc_hd__mux2_1
X_7127__55 _7127__55/A vssd1 vssd1 vccd1 vccd1 _8282_/CLK sky130_fd_sc_hd__inv_2
X_7361_ _7361_/A _7361_/B vssd1 vssd1 vccd1 vccd1 _7361_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3024_ clkbuf_0__3024_/X vssd1 vssd1 vccd1 vccd1 _6171__180/A sky130_fd_sc_hd__clkbuf_4
X_6243_ _8018_/Q _6238_/X _6236_/X _6239_/X _7807_/Q vssd1 vssd1 vccd1 vccd1 _7807_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_103_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5125_ _5125_/A vssd1 vssd1 vccd1 vccd1 _5205_/S sky130_fd_sc_hd__buf_2
X_5056_ _5182_/B vssd1 vssd1 vccd1 vccd1 _5252_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4007_ _4036_/S vssd1 vssd1 vccd1 vccd1 _4024_/S sky130_fd_sc_hd__buf_2
X_6308__209 _6309__210/A vssd1 vssd1 vccd1 vccd1 _7839_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5958_ _5958_/A vssd1 vssd1 vccd1 vccd1 _5958_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _7958_/Q _7942_/Q _4909_/S vssd1 vssd1 vccd1 vccd1 _4909_/X sky130_fd_sc_hd__mux2_1
X_5889_ _5889_/A vssd1 vssd1 vccd1 vccd1 _5889_/X sky130_fd_sc_hd__clkbuf_1
X_7628_ _8487_/Q _7613_/A _7627_/X _7543_/X vssd1 vssd1 vccd1 vccd1 _8486_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7559_ _6847_/A _7542_/X _7555_/X _7521_/B vssd1 vssd1 vccd1 vccd1 _7560_/B sky130_fd_sc_hd__o22a_1
X_7669__45 _7669__45/A vssd1 vssd1 vccd1 vccd1 _8514_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6881__378 _6881__378/A vssd1 vssd1 vccd1 vccd1 _8092_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7100__534 _7101__535/A vssd1 vssd1 vccd1 vccd1 _8261_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3438_ clkbuf_0__3438_/X vssd1 vssd1 vccd1 vccd1 _7006_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_wb_clk_i clkbuf_opt_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8479_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6294__198 _6294__198/A vssd1 vssd1 vccd1 vccd1 _7828_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3642_ clkbuf_0__3642_/X vssd1 vssd1 vccd1 vccd1 _7416__137/A sky130_fd_sc_hd__clkbuf_4
X_6861_ _7505_/A _8459_/Q _6860_/X vssd1 vssd1 vccd1 vccd1 _7614_/A sky130_fd_sc_hd__or3b_2
X_5812_ _5812_/A vssd1 vssd1 vccd1 vccd1 _7835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6792_ _8474_/Q _6857_/D vssd1 vssd1 vccd1 vccd1 _6793_/B sky130_fd_sc_hd__xnor2_4
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5743_ _7913_/Q _5566_/A _5743_/S vssd1 vssd1 vccd1 vccd1 _5744_/A sky130_fd_sc_hd__mux2_1
X_8531_ _8531_/CLK _8531_/D vssd1 vssd1 vccd1 vccd1 _8531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5674_ _5674_/A vssd1 vssd1 vccd1 vccd1 _7944_/D sky130_fd_sc_hd__clkbuf_1
X_8462_ _8487_/CLK _8462_/D vssd1 vssd1 vccd1 vccd1 _8462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6715__318 _6716__319/A vssd1 vssd1 vccd1 vccd1 _8028_/CLK sky130_fd_sc_hd__inv_2
X_8393_ _8393_/CLK _8393_/D vssd1 vssd1 vccd1 vccd1 _8393_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3472_ _7159_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3472_/X sky130_fd_sc_hd__clkbuf_16
X_4625_ _4876_/A vssd1 vssd1 vccd1 vccd1 _4810_/S sky130_fd_sc_hd__buf_4
X_4556_ _4556_/A vssd1 vssd1 vccd1 vccd1 _8218_/D sky130_fd_sc_hd__clkbuf_1
X_7344_ _7344_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _7344_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4487_ _8106_/Q vssd1 vssd1 vccd1 vccd1 _4487_/X sky130_fd_sc_hd__clkbuf_2
X_7275_ _7727_/B _7258_/B _7272_/X _7273_/Y _7274_/Y vssd1 vssd1 vccd1 vccd1 _7275_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6226_ _6225_/X _8008_/Q _6219_/X _6221_/X _7797_/Q vssd1 vssd1 vccd1 vccd1 _7797_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_58_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6034_/X _7901_/Q _6063_/A _6156_/X vssd1 vssd1 vccd1 vccd1 _6157_/X sky130_fd_sc_hd__a31o_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _8132_/Q _5040_/X _5348_/A _5105_/X _5107_/X vssd1 vssd1 vccd1 vccd1 _5108_/X
+ sky130_fd_sc_hd__a221o_1
X_6088_ _7866_/Q input6/X _6092_/S vssd1 vssd1 vccd1 vccd1 _6088_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5039_ _8134_/Q vssd1 vssd1 vccd1 vccd1 _5041_/A sky130_fd_sc_hd__inv_2
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6167__176 _6170__179/A vssd1 vssd1 vccd1 vccd1 _7763_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8556__254 vssd1 vssd1 vccd1 vccd1 partID[6] _8556__254/LO sky130_fd_sc_hd__conb_1
XFILLER_44_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4410_ _4388_/X _8272_/Q _4410_/S vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5390_ _5859_/A _5733_/B vssd1 vssd1 vccd1 vccd1 _5408_/S sky130_fd_sc_hd__or2_2
X_4341_ _4341_/A vssd1 vssd1 vccd1 vccd1 _8300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4272_ _4272_/A vssd1 vssd1 vccd1 vccd1 _8326_/D sky130_fd_sc_hd__clkbuf_1
X_6011_ _8008_/Q _6019_/B vssd1 vssd1 vccd1 vccd1 _6012_/A sky130_fd_sc_hd__and2_1
XFILLER_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7962_ _7962_/CLK _7962_/D vssd1 vssd1 vccd1 vccd1 _7962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6913_ _8487_/Q _7008_/C vssd1 vssd1 vccd1 vccd1 _6914_/A sky130_fd_sc_hd__and2_1
X_7893_ _8520_/CLK _7893_/D vssd1 vssd1 vccd1 vccd1 _7893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6844_ _7247_/A _7548_/S vssd1 vssd1 vccd1 vccd1 _6844_/X sky130_fd_sc_hd__or2_1
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3987_ _4002_/S vssd1 vssd1 vccd1 vccd1 _3996_/S sky130_fd_sc_hd__buf_2
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8514_ _8514_/CLK _8514_/D vssd1 vssd1 vccd1 vccd1 _8514_/Q sky130_fd_sc_hd__dfxtp_1
X_5726_ _5726_/A vssd1 vssd1 vccd1 vccd1 _7921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6574__263 _6574__263/A vssd1 vssd1 vccd1 vccd1 _7941_/CLK sky130_fd_sc_hd__inv_2
X_8445_ _8445_/CLK _8445_/D vssd1 vssd1 vccd1 vccd1 _8445_/Q sky130_fd_sc_hd__dfxtp_1
X_5657_ _7951_/Q _5596_/X _5659_/S vssd1 vssd1 vccd1 vccd1 _5658_/A sky130_fd_sc_hd__mux2_1
X_8376_ _8376_/CLK _8376_/D vssd1 vssd1 vccd1 vccd1 _8376_/Q sky130_fd_sc_hd__dfxtp_1
X_7442__158 _7444__160/A vssd1 vssd1 vccd1 vccd1 _8415_/CLK sky130_fd_sc_hd__inv_2
X_5588_ _7986_/Q _4520_/X _5591_/S vssd1 vssd1 vccd1 vccd1 _5589_/A sky130_fd_sc_hd__mux2_1
X_4608_ _8195_/Q _4178_/X _4614_/S vssd1 vssd1 vccd1 vccd1 _4609_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3455_ _7077_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3455_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4539_ _4385_/X _8225_/Q _4541_/S vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7327_ _8350_/Q _7318_/X _7326_/X _7216_/B vssd1 vssd1 vccd1 vccd1 _7328_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7258_ _8539_/Q _7258_/B vssd1 vssd1 vccd1 vccd1 _7262_/C sky130_fd_sc_hd__nand2_1
XFILLER_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6209_ _6208_/X _7998_/Q _6202_/X _6204_/X _7787_/Q vssd1 vssd1 vccd1 vccd1 _7787_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_100_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3410_ clkbuf_0__3410_/X vssd1 vssd1 vccd1 vccd1 _6895__390/A sky130_fd_sc_hd__clkbuf_4
X_3910_ _3910_/A vssd1 vssd1 vccd1 vccd1 _8513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4890_ _4441_/X _4629_/X _4889_/X _4857_/X vssd1 vssd1 vccd1 vccd1 _8180_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3841_ _5345_/A _8114_/Q vssd1 vssd1 vccd1 vccd1 _5034_/C sky130_fd_sc_hd__or2_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5511_ _5511_/A vssd1 vssd1 vccd1 vccd1 _8041_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3272_ clkbuf_0__3272_/X vssd1 vssd1 vccd1 vccd1 _6718_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6491_ _6491_/A vssd1 vssd1 vccd1 vccd1 _7887_/D sky130_fd_sc_hd__clkbuf_1
X_5442_ _3978_/X _8074_/Q _5444_/S vssd1 vssd1 vccd1 vccd1 _5443_/A sky130_fd_sc_hd__mux2_1
X_8230_ _8230_/CLK _8230_/D vssd1 vssd1 vccd1 vccd1 _8230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5373_ _5373_/A vssd1 vssd1 vccd1 vccd1 _8102_/D sky130_fd_sc_hd__clkbuf_1
X_8161_ _8161_/CLK _8161_/D vssd1 vssd1 vccd1 vccd1 _8161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8092_ _8092_/CLK _8092_/D vssd1 vssd1 vccd1 vccd1 _8092_/Q sky130_fd_sc_hd__dfxtp_1
X_4324_ _4280_/X _8307_/Q _4330_/S vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4255_ _4255_/A vssd1 vssd1 vccd1 vccd1 _8335_/D sky130_fd_sc_hd__clkbuf_1
X_4186_ _4186_/A vssd1 vssd1 vccd1 vccd1 _8391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7945_ _7945_/CLK _7945_/D vssd1 vssd1 vccd1 vccd1 _7945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7876_ _8551_/CLK _7876_/D vssd1 vssd1 vccd1 vccd1 _7876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6827_ _8544_/Q _7576_/A _7576_/B vssd1 vssd1 vccd1 vccd1 _6827_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6758_ _6248_/A _7747_/A _6762_/S vssd1 vssd1 vccd1 vccd1 _6759_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5709_ _7928_/Q _5593_/X _5713_/S vssd1 vssd1 vccd1 vccd1 _5710_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6689_ _6689_/A vssd1 vssd1 vccd1 vccd1 _8013_/D sky130_fd_sc_hd__clkbuf_1
X_8428_ _8428_/CLK _8428_/D vssd1 vssd1 vccd1 vccd1 _8428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3438_ _6993_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3438_/X sky130_fd_sc_hd__clkbuf_16
X_8359_ _8368_/CLK _8359_/D vssd1 vssd1 vccd1 vccd1 _8359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6767__355 _6767__355/A vssd1 vssd1 vccd1 vccd1 _8068_/CLK sky130_fd_sc_hd__inv_2
X_6728__328 _6730__330/A vssd1 vssd1 vccd1 vccd1 _8038_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7166__86 _7170__90/A vssd1 vssd1 vccd1 vccd1 _8313_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4040_ _4055_/S vssd1 vssd1 vccd1 vccd1 _4049_/S sky130_fd_sc_hd__buf_2
XFILLER_84_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6525__224 _6526__225/A vssd1 vssd1 vccd1 vccd1 _7902_/CLK sky130_fd_sc_hd__inv_2
X_5991_ _5991_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5992_/A sky130_fd_sc_hd__and2_1
XFILLER_91_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7730_ _7730_/A vssd1 vssd1 vccd1 vccd1 _8539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4942_ _4929_/A _4945_/B _7010_/A vssd1 vssd1 vccd1 vccd1 _4943_/B sky130_fd_sc_hd__a21o_1
X_4873_ _8160_/Q _8198_/Q _4873_/S vssd1 vssd1 vccd1 vccd1 _4873_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6612_ _6612_/A vssd1 vssd1 vccd1 vccd1 _7968_/D sky130_fd_sc_hd__clkbuf_1
X_7592_ _7600_/A _7592_/B vssd1 vssd1 vccd1 vccd1 _8473_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1_0__3255_ clkbuf_0__3255_/X vssd1 vssd1 vccd1 vccd1 _6584__271/A sky130_fd_sc_hd__clkbuf_4
X_6474_ _5982_/A _7880_/Q _6476_/S vssd1 vssd1 vccd1 vccd1 _6475_/A sky130_fd_sc_hd__mux2_1
X_8213_ _8213_/CLK _8213_/D vssd1 vssd1 vccd1 vccd1 _8213_/Q sky130_fd_sc_hd__dfxtp_1
X_5425_ _5425_/A vssd1 vssd1 vccd1 vccd1 _8083_/D sky130_fd_sc_hd__clkbuf_1
X_8144_ _8144_/CLK _8144_/D vssd1 vssd1 vccd1 vccd1 _8144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5356_ _5356_/A _5356_/B vssd1 vssd1 vccd1 vccd1 _5356_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8075_ _8075_/CLK _8075_/D vssd1 vssd1 vccd1 vccd1 _8075_/Q sky130_fd_sc_hd__dfxtp_1
X_5287_ _8039_/Q _8066_/Q _5290_/S vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4307_ _4307_/A vssd1 vssd1 vccd1 vccd1 _8315_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_5 _7821_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4238_ _5641_/A _5555_/A vssd1 vssd1 vccd1 vccd1 _4254_/S sky130_fd_sc_hd__nor2_2
Xclkbuf_1_0_0__3471_ clkbuf_0__3471_/X vssd1 vssd1 vccd1 vccd1 _7158__80/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4169_ _8106_/Q vssd1 vssd1 vccd1 vccd1 _4169_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7928_ _7928_/CLK _7928_/D vssd1 vssd1 vccd1 vccd1 _7928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7859_ _8551_/CLK _7859_/D vssd1 vssd1 vccd1 vccd1 _7859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6628__292 _6628__292/A vssd1 vssd1 vccd1 vccd1 _7978_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967__429 _6968__430/A vssd1 vssd1 vccd1 vccd1 _8153_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5210_ _8438_/Q _5207_/X _5101_/S _5209_/X vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__o211a_1
XFILLER_6_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6190_ _6210_/A vssd1 vssd1 vccd1 vccd1 _6202_/A sky130_fd_sc_hd__buf_4
X_5141_ _7843_/Q _8051_/Q _8330_/Q _8078_/Q _5273_/S _5068_/X vssd1 vssd1 vccd1 vccd1
+ _5141_/X sky130_fd_sc_hd__mux4_2
X_5072_ _5221_/A vssd1 vssd1 vccd1 vccd1 _5235_/A sky130_fd_sc_hd__buf_2
X_8599__246 vssd1 vssd1 vccd1 vccd1 _8599__246/HI versionID[0] sky130_fd_sc_hd__conb_1
X_4023_ _4289_/A vssd1 vssd1 vccd1 vccd1 _4023_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7119__550 _7119__550/A vssd1 vssd1 vccd1 vccd1 _8277_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5974_ _5974_/A vssd1 vssd1 vccd1 vccd1 _5974_/X sky130_fd_sc_hd__clkbuf_1
X_7713_ _5937_/A _7710_/X _7700_/A vssd1 vssd1 vccd1 vccd1 _7713_/X sky130_fd_sc_hd__a21bo_1
X_4925_ _4944_/B vssd1 vssd1 vccd1 vccd1 _4925_/Y sky130_fd_sc_hd__inv_2
X_4856_ _4713_/X _8181_/Q _4712_/X _4855_/X vssd1 vssd1 vccd1 vccd1 _4856_/X sky130_fd_sc_hd__a211o_1
X_7644_ _7644_/A _7646_/B _7646_/C vssd1 vssd1 vccd1 vccd1 _7645_/A sky130_fd_sc_hd__and3_1
X_7575_ _7575_/A vssd1 vssd1 vccd1 vccd1 _7575_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3307_ clkbuf_0__3307_/X vssd1 vssd1 vccd1 vccd1 _6723__325/A sky130_fd_sc_hd__clkbuf_4
X_4787_ _4803_/A vssd1 vssd1 vccd1 vccd1 _4787_/X sky130_fd_sc_hd__clkbuf_2
X_7050__494 _7051__495/A vssd1 vssd1 vccd1 vccd1 _8221_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6457_ _7874_/Q _6328_/A _6437_/A _6456_/X _6435_/A vssd1 vssd1 vccd1 vccd1 _7874_/D
+ sky130_fd_sc_hd__a221o_1
X_5408_ _5387_/X _8090_/Q _5408_/S vssd1 vssd1 vccd1 vccd1 _5409_/A sky130_fd_sc_hd__mux2_1
X_6388_ _6521_/A vssd1 vssd1 vccd1 vccd1 _6388_/X sky130_fd_sc_hd__buf_2
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8127_ _8127_/CLK _8127_/D vssd1 vssd1 vccd1 vccd1 _8127_/Q sky130_fd_sc_hd__dfxtp_1
X_5339_ _6941_/B vssd1 vssd1 vccd1 vccd1 _5339_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8058_ _8058_/CLK _8058_/D vssd1 vssd1 vccd1 vccd1 _8058_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3454_ clkbuf_0__3454_/X vssd1 vssd1 vccd1 vccd1 _7076__515/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7009_ _7009_/A vssd1 vssd1 vccd1 vccd1 _8187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5690_ _5690_/A vssd1 vssd1 vccd1 vccd1 _7937_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4710_ _4713_/A _8185_/Q _4947_/A _4709_/X _4712_/A vssd1 vssd1 vccd1 vccd1 _4710_/X
+ sky130_fd_sc_hd__a221o_1
X_4641_ _4658_/B _4783_/A vssd1 vssd1 vccd1 vccd1 _4726_/A sky130_fd_sc_hd__or2_1
XFILLER_116_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4572_ _4572_/A vssd1 vssd1 vccd1 vccd1 _8211_/D sky130_fd_sc_hd__clkbuf_1
X_7360_ _8361_/Q _7360_/B _7360_/C _7360_/D vssd1 vssd1 vccd1 vccd1 _7361_/B sky130_fd_sc_hd__or4_1
Xclkbuf_1_1_0__3023_ clkbuf_0__3023_/X vssd1 vssd1 vccd1 vccd1 _6184_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6242_ _8017_/Q _6238_/X _6236_/X _6239_/X _7806_/Q vssd1 vssd1 vccd1 vccd1 _7806_/D
+ sky130_fd_sc_hd__o32a_1
X_7397__122 _7400__125/A vssd1 vssd1 vccd1 vccd1 _8379_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5124_ _8307_/Q _8299_/Q _8291_/Q _8315_/Q _5095_/X _5088_/X vssd1 vssd1 vccd1 vccd1
+ _5124_/X sky130_fd_sc_hd__mux4_1
X_5055_ _5055_/A vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4006_ _5787_/A _5805_/B vssd1 vssd1 vccd1 vccd1 _4036_/S sky130_fd_sc_hd__or2_2
XFILLER_84_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5957_ _5957_/A _5965_/B vssd1 vssd1 vccd1 vccd1 _5958_/A sky130_fd_sc_hd__or2_1
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4908_ _4955_/B _4906_/X _4907_/X vssd1 vssd1 vccd1 vccd1 _4908_/Y sky130_fd_sc_hd__o21ai_1
X_5888_ _6248_/A _5890_/B vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__and2_1
XFILLER_21_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7627_ _8486_/Q _7601_/X vssd1 vssd1 vccd1 vccd1 _7627_/X sky130_fd_sc_hd__or2b_1
X_4839_ _4833_/X _4835_/X _4694_/X _4838_/X vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__a211o_1
X_6538__234 _6538__234/A vssd1 vssd1 vccd1 vccd1 _7912_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7406__129 _7407__130/A vssd1 vssd1 vccd1 vccd1 _8386_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7558_ _7567_/A _7558_/B vssd1 vssd1 vccd1 vccd1 _8463_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6509_ _8011_/Q _7896_/Q _6509_/S vssd1 vssd1 vccd1 vccd1 _6510_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3437_ clkbuf_0__3437_/X vssd1 vssd1 vccd1 vccd1 _6992__450/A sky130_fd_sc_hd__clkbuf_4
X_6922__398 _6924__400/A vssd1 vssd1 vccd1 vccd1 _8120_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3641_ clkbuf_0__3641_/X vssd1 vssd1 vccd1 vccd1 _7413__135/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6860_ _6860_/A _6860_/B _6860_/C _6860_/D vssd1 vssd1 vccd1 vccd1 _6860_/X sky130_fd_sc_hd__and4_1
XFILLER_35_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5811_ _3966_/X _7835_/Q _5815_/S vssd1 vssd1 vccd1 vccd1 _5812_/A sky130_fd_sc_hd__mux2_1
X_6791_ _8473_/Q _6796_/A _6818_/A _6795_/A vssd1 vssd1 vccd1 vccd1 _6857_/D sky130_fd_sc_hd__and4_2
XFILLER_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8530_ _8530_/CLK _8530_/D vssd1 vssd1 vccd1 vccd1 _8530_/Q sky130_fd_sc_hd__dfxtp_1
X_5742_ _5742_/A vssd1 vssd1 vccd1 vccd1 _7914_/D sky130_fd_sc_hd__clkbuf_1
X_5673_ _5569_/X _7944_/Q _5677_/S vssd1 vssd1 vccd1 vccd1 _5674_/A sky130_fd_sc_hd__mux2_1
X_8461_ _8487_/CLK _8461_/D vssd1 vssd1 vccd1 vccd1 _8461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8392_ _8392_/CLK _8392_/D vssd1 vssd1 vccd1 vccd1 _8392_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3471_ _7153_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3471_/X sky130_fd_sc_hd__clkbuf_16
X_4624_ _4766_/B vssd1 vssd1 vccd1 vccd1 _4876_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4555_ _4428_/X _8218_/Q _4559_/S vssd1 vssd1 vccd1 vccd1 _4556_/A sky130_fd_sc_hd__mux2_1
X_7343_ _7348_/A _7343_/B vssd1 vssd1 vccd1 vccd1 _8356_/D sky130_fd_sc_hd__nor2_1
X_6314__214 _6315__215/A vssd1 vssd1 vccd1 vccd1 _7844_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4486_ _4486_/A vssd1 vssd1 vccd1 vccd1 _8246_/D sky130_fd_sc_hd__clkbuf_1
X_7274_ _7220_/A _7220_/B _8541_/Q vssd1 vssd1 vccd1 vccd1 _7274_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6225_ _6235_/A vssd1 vssd1 vccd1 vccd1 _6225_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ input35/X input2/X _5969_/B _6153_/X _7637_/B vssd1 vssd1 vccd1 vccd1 _6156_/X
+ sky130_fd_sc_hd__o311a_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5107_/A vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6087_ _6075_/X _6085_/X _6086_/X _6083_/X vssd1 vssd1 vccd1 vccd1 _6087_/X sky130_fd_sc_hd__o211a_1
XFILLER_85_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5038_ _5038_/A vssd1 vssd1 vccd1 vccd1 _5038_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7648__27 _7651__30/A vssd1 vssd1 vccd1 vccd1 _8496_/CLK sky130_fd_sc_hd__inv_2
X_4340_ _4275_/X _8300_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4341_/A sky130_fd_sc_hd__mux2_1
X_4271_ _8326_/Q _4193_/X _4273_/S vssd1 vssd1 vccd1 vccd1 _4272_/A sky130_fd_sc_hd__mux2_1
X_6010_ _6010_/A vssd1 vssd1 vccd1 vccd1 _6019_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7961_ _7961_/CLK _7961_/D vssd1 vssd1 vccd1 vccd1 _7961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6721__323 _6723__325/A vssd1 vssd1 vccd1 vccd1 _8033_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6912_ _6912_/A vssd1 vssd1 vccd1 vccd1 _8112_/D sky130_fd_sc_hd__clkbuf_1
X_7892_ _8520_/CLK _7892_/D vssd1 vssd1 vccd1 vccd1 _7892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6843_ _7247_/A _7548_/S vssd1 vssd1 vccd1 vccd1 _6843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6774_ _6780_/A vssd1 vssd1 vccd1 vccd1 _6774_/X sky130_fd_sc_hd__buf_1
X_3986_ _4531_/A _5805_/B vssd1 vssd1 vccd1 vccd1 _4002_/S sky130_fd_sc_hd__or2_2
X_8513_ _8513_/CLK _8513_/D vssd1 vssd1 vccd1 vccd1 _8513_/Q sky130_fd_sc_hd__dfxtp_1
X_5725_ _7921_/Q _5590_/X _5725_/S vssd1 vssd1 vccd1 vccd1 _5726_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8444_ _8444_/CLK _8444_/D vssd1 vssd1 vccd1 vccd1 _8444_/Q sky130_fd_sc_hd__dfxtp_1
X_5656_ _5656_/A vssd1 vssd1 vccd1 vccd1 _7952_/D sky130_fd_sc_hd__clkbuf_1
X_4607_ _4607_/A vssd1 vssd1 vccd1 vccd1 _8196_/D sky130_fd_sc_hd__clkbuf_1
X_8375_ _8375_/CLK _8375_/D vssd1 vssd1 vccd1 vccd1 _8375_/Q sky130_fd_sc_hd__dfxtp_1
X_5587_ _5587_/A vssd1 vssd1 vccd1 vccd1 _7987_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3454_ _7071_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3454_/X sky130_fd_sc_hd__clkbuf_16
X_4538_ _4538_/A vssd1 vssd1 vccd1 vccd1 _8226_/D sky130_fd_sc_hd__clkbuf_1
X_7326_ _7326_/A vssd1 vssd1 vccd1 vccd1 _7326_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4469_ _8252_/Q _4465_/X _4479_/S vssd1 vssd1 vccd1 vccd1 _4470_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7257_ _7257_/A _7255_/X vssd1 vssd1 vccd1 vccd1 _7258_/B sky130_fd_sc_hd__or2b_1
X_6173__181 _6175__183/A vssd1 vssd1 vccd1 vccd1 _7768_/CLK sky130_fd_sc_hd__inv_2
X_6208_ _6235_/A vssd1 vssd1 vccd1 vccd1 _6208_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6139_ _6139_/A vssd1 vssd1 vccd1 vccd1 _6139_/X sky130_fd_sc_hd__clkbuf_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6894__389 _6895__390/A vssd1 vssd1 vccd1 vccd1 _8103_/CLK sky130_fd_sc_hd__inv_2
X_3840_ _8119_/Q vssd1 vssd1 vccd1 vccd1 _5345_/A sky130_fd_sc_hd__inv_2
X_7113__545 _7113__545/A vssd1 vssd1 vccd1 vccd1 _8272_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5510_ _8041_/Q _4289_/A _5510_/S vssd1 vssd1 vccd1 vccd1 _5511_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3271_ clkbuf_0__3271_/X vssd1 vssd1 vccd1 vccd1 _6755_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6490_ _5997_/A _7887_/Q _6498_/S vssd1 vssd1 vccd1 vccd1 _6491_/A sky130_fd_sc_hd__mux2_1
X_5441_ _5441_/A vssd1 vssd1 vccd1 vccd1 _8075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5372_ _4432_/X _8102_/Q _5376_/S vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__mux2_1
X_8160_ _8160_/CLK _8160_/D vssd1 vssd1 vccd1 vccd1 _8160_/Q sky130_fd_sc_hd__dfxtp_1
X_8091_ _8091_/CLK _8091_/D vssd1 vssd1 vccd1 vccd1 _8091_/Q sky130_fd_sc_hd__dfxtp_1
X_4323_ _4323_/A vssd1 vssd1 vccd1 vccd1 _8308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4254_ _8335_/Q _4169_/X _4254_/S vssd1 vssd1 vccd1 vccd1 _4255_/A sky130_fd_sc_hd__mux2_1
X_7007__461 _7011__462/A vssd1 vssd1 vccd1 vccd1 _8186_/CLK sky130_fd_sc_hd__inv_2
X_4185_ _8391_/Q _4184_/X _4188_/S vssd1 vssd1 vccd1 vccd1 _4186_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7944_ _7944_/CLK _7944_/D vssd1 vssd1 vccd1 vccd1 _7944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7875_ _8063_/CLK _7875_/D vssd1 vssd1 vccd1 vccd1 _7875_/Q sky130_fd_sc_hd__dfxtp_1
X_6826_ _8467_/Q _6849_/B _6830_/B _8468_/Q vssd1 vssd1 vccd1 vccd1 _7576_/B sky130_fd_sc_hd__a31o_1
XFILLER_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5708_ _5708_/A vssd1 vssd1 vccd1 vccd1 _7929_/D sky130_fd_sc_hd__clkbuf_1
X_7014__465 _7014__465/A vssd1 vssd1 vccd1 vccd1 _8192_/CLK sky130_fd_sc_hd__inv_2
X_3969_ _8492_/Q vssd1 vssd1 vccd1 vccd1 _3969_/X sky130_fd_sc_hd__buf_4
Xclkbuf_1_1_0__3469_ clkbuf_0__3469_/X vssd1 vssd1 vccd1 vccd1 _7151__75/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6688_ _5952_/A _8013_/Q _6688_/S vssd1 vssd1 vccd1 vccd1 _6689_/A sky130_fd_sc_hd__mux2_1
X_5639_ _5575_/X _7958_/Q _5639_/S vssd1 vssd1 vccd1 vccd1 _5640_/A sky130_fd_sc_hd__mux2_1
X_8427_ _8427_/CLK _8427_/D vssd1 vssd1 vccd1 vccd1 _8427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8358_ _8358_/CLK _8358_/D vssd1 vssd1 vccd1 vccd1 _8358_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3437_ _6987_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3437_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_5_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7309_ _7326_/A vssd1 vssd1 vccd1 vccd1 _7310_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7493__25 _7493__25/A vssd1 vssd1 vccd1 vccd1 _8457_/CLK sky130_fd_sc_hd__inv_2
X_8289_ _8289_/CLK _8289_/D vssd1 vssd1 vccd1 vccd1 _8289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7391__117 _7392__118/A vssd1 vssd1 vccd1 vccd1 _8374_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8601__248 vssd1 vssd1 vccd1 vccd1 _8601__248/HI versionID[2] sky130_fd_sc_hd__conb_1
XFILLER_49_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5990_ _5990_/A vssd1 vssd1 vccd1 vccd1 _5990_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ _6902_/A vssd1 vssd1 vccd1 vccd1 _7010_/A sky130_fd_sc_hd__inv_2
X_4872_ _4673_/X _4861_/X _4864_/X _4871_/X _4684_/X vssd1 vssd1 vccd1 vccd1 _4872_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_60_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6611_ _8181_/Q _8167_/D vssd1 vssd1 vccd1 vccd1 _6612_/A sky130_fd_sc_hd__and2_1
X_7591_ _6802_/A _7588_/X _7547_/X _7528_/B vssd1 vssd1 vccd1 vccd1 _7592_/B sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_9_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8480_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3254_ clkbuf_0__3254_/X vssd1 vssd1 vccd1 vccd1 _6582__270/A sky130_fd_sc_hd__clkbuf_4
X_6473_ _6473_/A vssd1 vssd1 vccd1 vccd1 _7879_/D sky130_fd_sc_hd__clkbuf_1
X_8212_ _8212_/CLK _8212_/D vssd1 vssd1 vccd1 vccd1 _8212_/Q sky130_fd_sc_hd__dfxtp_1
X_5424_ _5383_/X _8083_/Q _5426_/S vssd1 vssd1 vccd1 vccd1 _5425_/A sky130_fd_sc_hd__mux2_1
Xoutput200 _6150_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[30] sky130_fd_sc_hd__buf_2
X_6532__229 _6533__230/A vssd1 vssd1 vccd1 vccd1 _7907_/CLK sky130_fd_sc_hd__inv_2
X_8143_ _8143_/CLK _8143_/D vssd1 vssd1 vccd1 vccd1 _8143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5355_ _5270_/X _5348_/X _5354_/Y _5339_/X vssd1 vssd1 vccd1 vccd1 _8116_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8074_ _8074_/CLK _8074_/D vssd1 vssd1 vccd1 vccd1 _8074_/Q sky130_fd_sc_hd__dfxtp_1
X_5286_ _5356_/B _5284_/X _5285_/X vssd1 vssd1 vccd1 vccd1 _5286_/Y sky130_fd_sc_hd__o21ai_1
X_4306_ _4280_/X _8315_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4307_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_6 _4379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_0__3470_ clkbuf_0__3470_/X vssd1 vssd1 vccd1 vccd1 _7165_/A sky130_fd_sc_hd__clkbuf_4
X_4237_ _5622_/A _4466_/B _4933_/C vssd1 vssd1 vccd1 vccd1 _5555_/A sky130_fd_sc_hd__or3b_4
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4168_ _4168_/A vssd1 vssd1 vccd1 vccd1 _8396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4099_ _4099_/A vssd1 vssd1 vccd1 vccd1 _8410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7927_ _7927_/CLK _7927_/D vssd1 vssd1 vccd1 vccd1 _7927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7858_ _8345_/CLK _7858_/D vssd1 vssd1 vccd1 vccd1 _7858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6809_ _8474_/Q _6857_/D _8475_/Q vssd1 vssd1 vccd1 vccd1 _7532_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6773__360 _6773__360/A vssd1 vssd1 vccd1 vccd1 _8073_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7789_ _8540_/CLK _7789_/D vssd1 vssd1 vccd1 vccd1 _7789_/Q sky130_fd_sc_hd__dfxtp_1
X_6734__333 _6736__335/A vssd1 vssd1 vccd1 vccd1 _8043_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7062__503 _7063__504/A vssd1 vssd1 vccd1 vccd1 _8230_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6587__274 _6588__275/A vssd1 vssd1 vccd1 vccd1 _7952_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7455__169 _7456__170/A vssd1 vssd1 vccd1 vccd1 _8426_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7139__65 _7139__65/A vssd1 vssd1 vccd1 vccd1 _8292_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5140_ _5055_/X _5137_/X _5139_/X vssd1 vssd1 vccd1 vccd1 _5140_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5071_ _5103_/B _5082_/B vssd1 vssd1 vccd1 vccd1 _5221_/A sky130_fd_sc_hd__or2_2
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4022_ _8491_/Q vssd1 vssd1 vccd1 vccd1 _4289_/A sky130_fd_sc_hd__buf_4
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5973_ _5973_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5974_/A sky130_fd_sc_hd__and2_1
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7712_ _7008_/A _7701_/X _7711_/X _7704_/X vssd1 vssd1 vccd1 vccd1 _8534_/D sky130_fd_sc_hd__o211a_1
X_4924_ _7008_/C vssd1 vssd1 vccd1 vccd1 _4924_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4855_ _4840_/X _4854_/X _4948_/A vssd1 vssd1 vccd1 vccd1 _4855_/X sky130_fd_sc_hd__o21a_1
X_7643_ _7643_/A vssd1 vssd1 vccd1 vccd1 _8493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4786_ _4786_/A vssd1 vssd1 vccd1 vccd1 _4803_/A sky130_fd_sc_hd__clkbuf_2
X_7574_ _8468_/Q vssd1 vssd1 vccd1 vccd1 _7574_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3306_ clkbuf_0__3306_/X vssd1 vssd1 vccd1 vccd1 _6717__320/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6456_ _8531_/Q _6456_/B _8064_/Q vssd1 vssd1 vccd1 vccd1 _6456_/X sky130_fd_sc_hd__and3_1
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5407_ _5407_/A vssd1 vssd1 vccd1 vccd1 _8091_/D sky130_fd_sc_hd__clkbuf_1
X_6387_ _7858_/Q _6328_/X _6386_/X vssd1 vssd1 vccd1 vccd1 _7858_/D sky130_fd_sc_hd__a21o_1
X_8126_ _8126_/CLK _8126_/D vssd1 vssd1 vccd1 vccd1 _8126_/Q sky130_fd_sc_hd__dfxtp_1
X_5338_ _5338_/A vssd1 vssd1 vccd1 vccd1 _8122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8057_ _8057_/CLK _8057_/D vssd1 vssd1 vccd1 vccd1 _8057_/Q sky130_fd_sc_hd__dfxtp_1
X_5269_ _8452_/Q _8190_/Q _5281_/S vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__mux2_1
X_7008_ _7008_/A _8081_/Q _7008_/C vssd1 vssd1 vccd1 vccd1 _7009_/A sky130_fd_sc_hd__and3_1
Xclkbuf_1_0_0__3453_ clkbuf_0__3453_/X vssd1 vssd1 vccd1 vccd1 _7070__510/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6973__434 _6973__434/A vssd1 vssd1 vccd1 vccd1 _8158_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6934__407 _6937__410/A vssd1 vssd1 vccd1 vccd1 _8129_/CLK sky130_fd_sc_hd__inv_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _4767_/A _4766_/B _8170_/Q vssd1 vssd1 vccd1 vccd1 _4783_/A sky130_fd_sc_hd__a21oi_2
X_7069__509 _7069__509/A vssd1 vssd1 vccd1 vccd1 _8236_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3314_ clkbuf_0__3314_/X vssd1 vssd1 vccd1 vccd1 _6780_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6310_ _6310_/A vssd1 vssd1 vccd1 vccd1 _6310_/X sky130_fd_sc_hd__buf_1
X_4571_ _3963_/X _8211_/Q _4577_/S vssd1 vssd1 vccd1 vccd1 _4572_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8566__213 vssd1 vssd1 vccd1 vccd1 _8566__213/HI core0Index[0] sky130_fd_sc_hd__conb_1
XFILLER_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6241_ _8016_/Q _6238_/X _6236_/X _6239_/X _7805_/Q vssd1 vssd1 vccd1 vccd1 _7805_/D
+ sky130_fd_sc_hd__o32a_1
X_6172_ _6184_/A vssd1 vssd1 vccd1 vccd1 _6172_/X sky130_fd_sc_hd__buf_1
XFILLER_111_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5123_ _8425_/Q _8323_/Q _8060_/Q _8275_/Q _5129_/A _5305_/S vssd1 vssd1 vccd1 vccd1
+ _5123_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7293__110 _7293__110/A vssd1 vssd1 vccd1 vccd1 _8339_/CLK sky130_fd_sc_hd__inv_2
X_5054_ _5167_/S vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__clkbuf_2
X_4005_ _4275_/A vssd1 vssd1 vccd1 vccd1 _4005_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _5956_/A vssd1 vssd1 vccd1 vccd1 _5965_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5887_ _5887_/A vssd1 vssd1 vccd1 vccd1 _5887_/X sky130_fd_sc_hd__clkbuf_1
X_4907_ _4811_/X _7950_/Q _7763_/Q _4791_/X _4739_/S vssd1 vssd1 vccd1 vccd1 _4907_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4838_ _4794_/X _4836_/X _4837_/X vssd1 vssd1 vccd1 vccd1 _4838_/X sky130_fd_sc_hd__o21a_1
X_7626_ _8486_/Q _7613_/A _7625_/X _7543_/X vssd1 vssd1 vccd1 vccd1 _8485_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4769_ _4786_/A vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__clkbuf_2
X_7557_ _7554_/Y _7542_/X _7555_/X _7556_/Y vssd1 vssd1 vccd1 vccd1 _7558_/B sky130_fd_sc_hd__o22a_1
XFILLER_107_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7488_ _7488_/A vssd1 vssd1 vccd1 vccd1 _7488_/X sky130_fd_sc_hd__buf_1
XFILLER_20_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6508_ _6508_/A vssd1 vssd1 vccd1 vccd1 _7895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6439_ _6456_/B vssd1 vssd1 vccd1 vccd1 _6452_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_96_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8109_ _8480_/CLK _8109_/D vssd1 vssd1 vccd1 vccd1 _8109_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_88_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3436_ clkbuf_0__3436_/X vssd1 vssd1 vccd1 vccd1 _6983__442/A sky130_fd_sc_hd__clkbuf_4
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _8358_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3640_ clkbuf_0__3640_/X vssd1 vssd1 vccd1 vccd1 _7405__128/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7001__456 _7002__457/A vssd1 vssd1 vccd1 vccd1 _8181_/CLK sky130_fd_sc_hd__inv_2
X_5810_ _5810_/A vssd1 vssd1 vccd1 vccd1 _7836_/D sky130_fd_sc_hd__clkbuf_1
X_6790_ _8468_/Q _8467_/Q _8466_/Q _8465_/Q vssd1 vssd1 vccd1 vccd1 _6795_/A sky130_fd_sc_hd__and4_1
XFILLER_35_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5741_ _7914_/Q _5650_/X _5743_/S vssd1 vssd1 vccd1 vccd1 _5742_/A sky130_fd_sc_hd__mux2_1
X_8460_ _8479_/CLK _8460_/D vssd1 vssd1 vccd1 vccd1 _8460_/Q sky130_fd_sc_hd__dfxtp_1
X_5672_ _5672_/A vssd1 vssd1 vccd1 vccd1 _7945_/D sky130_fd_sc_hd__clkbuf_1
X_8391_ _8391_/CLK _8391_/D vssd1 vssd1 vccd1 vccd1 _8391_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3470_ _7152_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3470_/X sky130_fd_sc_hd__clkbuf_16
X_4623_ _8168_/Q vssd1 vssd1 vccd1 vccd1 _4766_/B sky130_fd_sc_hd__clkbuf_2
X_4554_ _4554_/A vssd1 vssd1 vccd1 vccd1 _8219_/D sky130_fd_sc_hd__clkbuf_1
X_7342_ _8356_/Q _7334_/X _7310_/A _7205_/B vssd1 vssd1 vccd1 vccd1 _7343_/B sky130_fd_sc_hd__o2bb2a_1
X_7273_ _7272_/B _7272_/C _7216_/A vssd1 vssd1 vccd1 vccd1 _7273_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4485_ _8246_/Q _4484_/X _4488_/S vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__mux2_1
X_6224_ _6217_/X _8007_/Q _6219_/X _6221_/X _7796_/Q vssd1 vssd1 vccd1 vccd1 _7796_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_112_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _7702_/A vssd1 vssd1 vccd1 vccd1 _7637_/B sky130_fd_sc_hd__buf_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _7790_/Q _6086_/B vssd1 vssd1 vccd1 vccd1 _6086_/X sky130_fd_sc_hd__or2_1
X_5106_ _5106_/A _7363_/A vssd1 vssd1 vccd1 vccd1 _5107_/A sky130_fd_sc_hd__and2_1
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5037_ _5106_/A _7363_/A vssd1 vssd1 vccd1 vccd1 _5038_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7412__134 _7413__135/A vssd1 vssd1 vccd1 vccd1 _8391_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5939_ _5939_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5940_/A sky130_fd_sc_hd__or2_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7609_ _7609_/A _7609_/B vssd1 vssd1 vccd1 vccd1 _7609_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput100 wbs_data_i[8] vssd1 vssd1 vccd1 vccd1 _5919_/A sky130_fd_sc_hd__buf_4
XFILLER_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4270_ _4270_/A vssd1 vssd1 vccd1 vccd1 _8327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7960_ _7960_/CLK _7960_/D vssd1 vssd1 vccd1 vccd1 _7960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6911_ _8486_/Q _6911_/B vssd1 vssd1 vccd1 vccd1 _6912_/A sky130_fd_sc_hd__and2_1
X_7891_ _8520_/CLK _7891_/D vssd1 vssd1 vccd1 vccd1 _7891_/Q sky130_fd_sc_hd__dfxtp_1
X_6842_ _7550_/A _6842_/B vssd1 vssd1 vccd1 vccd1 _6842_/Y sky130_fd_sc_hd__xnor2_1
X_3985_ _4301_/B _4076_/A _4301_/A vssd1 vssd1 vccd1 vccd1 _5805_/B sky130_fd_sc_hd__or3b_4
X_8512_ _8512_/CLK _8512_/D vssd1 vssd1 vccd1 vccd1 _8512_/Q sky130_fd_sc_hd__dfxtp_1
X_5724_ _5724_/A vssd1 vssd1 vccd1 vccd1 _7922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8443_ _8443_/CLK _8443_/D vssd1 vssd1 vccd1 vccd1 _8443_/Q sky130_fd_sc_hd__dfxtp_1
X_5655_ _7952_/Q _5593_/X _5659_/S vssd1 vssd1 vccd1 vccd1 _5656_/A sky130_fd_sc_hd__mux2_1
X_8374_ _8374_/CLK _8374_/D vssd1 vssd1 vccd1 vccd1 _8374_/Q sky130_fd_sc_hd__dfxtp_1
X_4606_ _8196_/Q _4172_/X _4614_/S vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3453_ _7065_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3453_/X sky130_fd_sc_hd__clkbuf_16
X_5586_ _7987_/Q _4517_/X _5591_/S vssd1 vssd1 vccd1 vccd1 _5587_/A sky130_fd_sc_hd__mux2_1
X_7325_ _7336_/A _7325_/B vssd1 vssd1 vccd1 vccd1 _8349_/D sky130_fd_sc_hd__nor2_1
X_4537_ _4382_/X _8226_/Q _4541_/S vssd1 vssd1 vccd1 vccd1 _4538_/A sky130_fd_sc_hd__mux2_1
X_4468_ _4488_/S vssd1 vssd1 vccd1 vccd1 _4479_/S sky130_fd_sc_hd__buf_2
X_7256_ _8539_/Q _7257_/A _7255_/X vssd1 vssd1 vccd1 vccd1 _7262_/B sky130_fd_sc_hd__or3b_1
XFILLER_89_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6207_ _6200_/X _7818_/Q _6202_/X _6204_/X _7786_/Q vssd1 vssd1 vccd1 vccd1 _7786_/D
+ sky130_fd_sc_hd__o32a_1
X_4399_ _4399_/A vssd1 vssd1 vccd1 vccd1 _8277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6138_ _6138_/A vssd1 vssd1 vccd1 vccd1 _6138_/X sky130_fd_sc_hd__clkbuf_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6069_ _6138_/A vssd1 vssd1 vccd1 vccd1 _6086_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6581__269 _6582__270/A vssd1 vssd1 vccd1 vccd1 _7947_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7178__96 _7179__97/A vssd1 vssd1 vccd1 vccd1 _8323_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7653__31 _7657__35/A vssd1 vssd1 vccd1 vccd1 _8500_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3270_ clkbuf_0__3270_/X vssd1 vssd1 vccd1 vccd1 _6637__300/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5440_ _3975_/X _8075_/Q _5444_/S vssd1 vssd1 vccd1 vccd1 _5441_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5371_ _5371_/A vssd1 vssd1 vccd1 vccd1 _8103_/D sky130_fd_sc_hd__clkbuf_1
X_8090_ _8090_/CLK _8090_/D vssd1 vssd1 vccd1 vccd1 _8090_/Q sky130_fd_sc_hd__dfxtp_1
X_4322_ _4275_/X _8308_/Q _4330_/S vssd1 vssd1 vccd1 vccd1 _4323_/A sky130_fd_sc_hd__mux2_1
X_4253_ _4253_/A vssd1 vssd1 vccd1 vccd1 _8336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4184_ _8492_/Q vssd1 vssd1 vccd1 vccd1 _4184_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7943_ _7943_/CLK _7943_/D vssd1 vssd1 vccd1 vccd1 _7943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7874_ _8548_/CLK _7874_/D vssd1 vssd1 vccd1 vccd1 _7874_/Q sky130_fd_sc_hd__dfxtp_1
X_6825_ _6853_/B vssd1 vssd1 vccd1 vccd1 _7576_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6756_ _6780_/A vssd1 vssd1 vccd1 vccd1 _6756_/X sky130_fd_sc_hd__buf_1
X_3968_ _3968_/A vssd1 vssd1 vccd1 vccd1 _8456_/D sky130_fd_sc_hd__clkbuf_1
X_7186__102 _7186__102/A vssd1 vssd1 vccd1 vccd1 _8329_/CLK sky130_fd_sc_hd__inv_2
X_5707_ _7929_/Q _5590_/X _5707_/S vssd1 vssd1 vccd1 vccd1 _5708_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3468_ clkbuf_0__3468_/X vssd1 vssd1 vccd1 vccd1 _7142__67/A sky130_fd_sc_hd__clkbuf_4
X_6687_ _6687_/A vssd1 vssd1 vccd1 vccd1 _8012_/D sky130_fd_sc_hd__clkbuf_1
X_3899_ _8492_/Q vssd1 vssd1 vccd1 vccd1 _3899_/X sky130_fd_sc_hd__buf_4
X_5638_ _5638_/A vssd1 vssd1 vccd1 vccd1 _7959_/D sky130_fd_sc_hd__clkbuf_1
X_8426_ _8426_/CLK _8426_/D vssd1 vssd1 vccd1 vccd1 _8426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7478__12 _7479__13/A vssd1 vssd1 vccd1 vccd1 _8444_/CLK sky130_fd_sc_hd__inv_2
X_5569_ _5569_/A vssd1 vssd1 vccd1 vccd1 _5569_/X sky130_fd_sc_hd__clkbuf_4
X_8357_ _8358_/CLK _8357_/D vssd1 vssd1 vccd1 vccd1 _8357_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3436_ _6981_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3436_/X sky130_fd_sc_hd__clkbuf_16
X_7308_ _7308_/A _7308_/B vssd1 vssd1 vccd1 vccd1 _7326_/A sky130_fd_sc_hd__or2_1
X_8288_ _8288_/CLK _8288_/D vssd1 vssd1 vccd1 vccd1 _8288_/Q sky130_fd_sc_hd__dfxtp_1
X_6960__425 _6960__425/A vssd1 vssd1 vccd1 vccd1 _8149_/CLK sky130_fd_sc_hd__inv_2
X_7239_ _8346_/Q _7311_/A vssd1 vssd1 vccd1 vccd1 _7240_/B sky130_fd_sc_hd__xor2_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4940_ _4141_/A _4925_/Y _4939_/X _4857_/X vssd1 vssd1 vccd1 vccd1 _8175_/D sky130_fd_sc_hd__o211a_1
X_4871_ _4865_/X _4867_/X _4694_/X _4870_/X vssd1 vssd1 vccd1 vccd1 _4871_/X sky130_fd_sc_hd__a211o_1
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7590_ _7600_/A _7590_/B vssd1 vssd1 vccd1 vccd1 _8472_/D sky130_fd_sc_hd__nor2_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6610_ _6610_/A vssd1 vssd1 vccd1 vccd1 _7967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3253_ clkbuf_0__3253_/X vssd1 vssd1 vccd1 vccd1 _6574__263/A sky130_fd_sc_hd__clkbuf_4
X_6472_ _5980_/A _7879_/Q _6476_/S vssd1 vssd1 vccd1 vccd1 _6473_/A sky130_fd_sc_hd__mux2_1
X_8211_ _8211_/CLK _8211_/D vssd1 vssd1 vccd1 vccd1 _8211_/Q sky130_fd_sc_hd__dfxtp_1
X_5423_ _5423_/A vssd1 vssd1 vccd1 vccd1 _8084_/D sky130_fd_sc_hd__clkbuf_1
Xoutput201 _6152_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[31] sky130_fd_sc_hd__buf_2
X_5354_ _5356_/A _5354_/B vssd1 vssd1 vccd1 vccd1 _5354_/Y sky130_fd_sc_hd__nand2_1
X_8142_ _8142_/CLK _8142_/D vssd1 vssd1 vccd1 vccd1 _8142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4305_ _4305_/A vssd1 vssd1 vccd1 vccd1 _8316_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_7 _5969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8073_ _8073_/CLK _8073_/D vssd1 vssd1 vccd1 vccd1 _8073_/Q sky130_fd_sc_hd__dfxtp_1
X_6647__306 _6649__308/A vssd1 vssd1 vccd1 vccd1 _7992_/CLK sky130_fd_sc_hd__inv_2
X_5285_ _8444_/Q _5180_/X _5239_/X _8436_/Q _5101_/S vssd1 vssd1 vccd1 vccd1 _5285_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4236_ _4236_/A vssd1 vssd1 vccd1 vccd1 _8371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4167_ _8396_/Q _4166_/X _4170_/S vssd1 vssd1 vccd1 vccd1 _4168_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4098_ _4005_/X _8410_/Q _4106_/S vssd1 vssd1 vccd1 vccd1 _4099_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7020__470 _7020__470/A vssd1 vssd1 vccd1 vccd1 _8197_/CLK sky130_fd_sc_hd__inv_2
X_7926_ _7926_/CLK _7926_/D vssd1 vssd1 vccd1 vccd1 _7926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7857_ _8345_/CLK _7857_/D vssd1 vssd1 vccd1 vccd1 _7857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6808_ _6808_/A _6808_/B _6808_/C _6808_/D vssd1 vssd1 vccd1 vccd1 _6860_/A sky130_fd_sc_hd__and4_1
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7788_ _8540_/CLK _7788_/D vssd1 vssd1 vccd1 vccd1 _7788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8409_ _8409_/CLK _8409_/D vssd1 vssd1 vccd1 vccd1 _8409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6594__279 _6594__279/A vssd1 vssd1 vccd1 vccd1 _7957_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6635__298 _6635__298/A vssd1 vssd1 vccd1 vccd1 _7984_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5070_ _5070_/A _5070_/B vssd1 vssd1 vccd1 vccd1 _5082_/B sky130_fd_sc_hd__nor2_1
X_4021_ _4021_/A vssd1 vssd1 vccd1 vccd1 _8439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5972_ _5972_/A vssd1 vssd1 vccd1 vccd1 _5972_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7711_ _5939_/A _7710_/X _7701_/A vssd1 vssd1 vccd1 vccd1 _7711_/X sky130_fd_sc_hd__a21bo_1
X_4923_ _6902_/A vssd1 vssd1 vccd1 vccd1 _7008_/C sky130_fd_sc_hd__clkbuf_2
X_4854_ _4740_/X _4843_/X _4846_/X _4853_/X _4638_/A vssd1 vssd1 vccd1 vccd1 _4854_/X
+ sky130_fd_sc_hd__o311a_1
X_7642_ _7642_/A _7646_/B _7646_/C vssd1 vssd1 vccd1 vccd1 _7643_/A sky130_fd_sc_hd__and3_1
X_4785_ _7985_/Q _8033_/Q _4866_/S vssd1 vssd1 vccd1 vccd1 _4785_/X sky130_fd_sc_hd__mux2_1
X_7573_ _7585_/A _7573_/B vssd1 vssd1 vccd1 vccd1 _8467_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6524_ _6191_/X _6272_/B _7680_/A vssd1 vssd1 vccd1 vccd1 _7901_/D sky130_fd_sc_hd__a21oi_1
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6455_ _7873_/Q _6442_/X _6437_/A _6454_/X _6435_/A vssd1 vssd1 vccd1 vccd1 _7873_/D
+ sky130_fd_sc_hd__a221o_1
X_5406_ _5383_/X _8091_/Q _5408_/S vssd1 vssd1 vccd1 vccd1 _5407_/A sky130_fd_sc_hd__mux2_1
X_6386_ _6331_/A _6383_/X _6385_/X _6367_/X vssd1 vssd1 vccd1 vccd1 _6386_/X sky130_fd_sc_hd__a31o_1
X_8125_ _8125_/CLK _8125_/D vssd1 vssd1 vccd1 vccd1 _8125_/Q sky130_fd_sc_hd__dfxtp_1
X_5337_ _5343_/A _5337_/B _5337_/C vssd1 vssd1 vccd1 vccd1 _5338_/A sky130_fd_sc_hd__and3_1
X_8056_ _8056_/CLK _8056_/D vssd1 vssd1 vccd1 vccd1 _8056_/Q sky130_fd_sc_hd__dfxtp_1
X_5268_ _5356_/B _5266_/X _5267_/X vssd1 vssd1 vccd1 vccd1 _5268_/Y sky130_fd_sc_hd__o21ai_1
X_4219_ _5602_/A _5823_/A vssd1 vssd1 vccd1 vccd1 _4235_/S sky130_fd_sc_hd__nor2_2
X_5199_ _8224_/Q _5196_/X _5198_/X _8208_/Q _5167_/S vssd1 vssd1 vccd1 vccd1 _5199_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3452_ clkbuf_0__3452_/X vssd1 vssd1 vccd1 vccd1 _7064__505/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7909_ _7909_/CLK _7909_/D vssd1 vssd1 vccd1 vccd1 _7909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7461__174 _7462__175/A vssd1 vssd1 vccd1 vccd1 _8431_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4570_ _4570_/A vssd1 vssd1 vccd1 vccd1 _8212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3021_ clkbuf_0__3021_/X vssd1 vssd1 vccd1 vccd1 _6961_/A sky130_fd_sc_hd__clkbuf_4
X_6240_ _8015_/Q _6238_/X _6236_/X _6239_/X _7804_/Q vssd1 vssd1 vccd1 vccd1 _7804_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5122_ _5318_/S vssd1 vssd1 vccd1 vccd1 _5305_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_69_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5053_ _5125_/A vssd1 vssd1 vccd1 vccd1 _5167_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_38_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4004_ _8495_/Q vssd1 vssd1 vccd1 vccd1 _4275_/A sky130_fd_sc_hd__buf_4
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5955_ _5955_/A vssd1 vssd1 vccd1 vccd1 _5955_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5886_ _6269_/C _5890_/B vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__and2_1
X_4906_ _7846_/Q _7771_/Q _4909_/S vssd1 vssd1 vccd1 vccd1 _4906_/X sky130_fd_sc_hd__mux2_1
X_4837_ _4811_/A _7952_/Q _7765_/Q _4797_/X _4733_/A vssd1 vssd1 vccd1 vccd1 _4837_/X
+ sky130_fd_sc_hd__o221a_1
X_7625_ _8485_/Q _7601_/X vssd1 vssd1 vccd1 vccd1 _7625_/X sky130_fd_sc_hd__or2b_1
XFILLER_119_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4768_ _4768_/A _4797_/A vssd1 vssd1 vccd1 vccd1 _4786_/A sky130_fd_sc_hd__nand2_2
X_7556_ _7556_/A _7556_/B vssd1 vssd1 vccd1 vccd1 _7556_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4699_ _4714_/A _4698_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _4699_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6507_ _8010_/Q _7895_/Q _6509_/S vssd1 vssd1 vccd1 vccd1 _6508_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6438_ _8537_/Q vssd1 vssd1 vccd1 vccd1 _6440_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6369_ _7855_/Q _6328_/X _6368_/X vssd1 vssd1 vccd1 vccd1 _7855_/D sky130_fd_sc_hd__a21o_1
X_8108_ _8480_/CLK _8108_/D vssd1 vssd1 vccd1 vccd1 _8108_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8039_ _8039_/CLK _8039_/D vssd1 vssd1 vccd1 vccd1 _8039_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3435_ clkbuf_0__3435_/X vssd1 vssd1 vccd1 vccd1 _6980__440/A sky130_fd_sc_hd__clkbuf_4
XFILLER_45_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7033__480 _7033__480/A vssd1 vssd1 vccd1 vccd1 _8207_/CLK sky130_fd_sc_hd__inv_2
X_8589__236 vssd1 vssd1 vccd1 vccd1 _8589__236/HI manufacturerID[8] sky130_fd_sc_hd__conb_1
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6747__344 _6748__345/A vssd1 vssd1 vccd1 vccd1 _8054_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7075__514 _7076__515/A vssd1 vssd1 vccd1 vccd1 _8241_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5740_ _5740_/A vssd1 vssd1 vccd1 vccd1 _7915_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5566_/X _7945_/Q _5671_/S vssd1 vssd1 vccd1 vccd1 _5672_/A sky130_fd_sc_hd__mux2_1
X_8390_ _8390_/CLK _8390_/D vssd1 vssd1 vccd1 vccd1 _8390_/Q sky130_fd_sc_hd__dfxtp_1
X_4622_ _4622_/A _4622_/B _4622_/C vssd1 vssd1 vccd1 vccd1 _4622_/X sky130_fd_sc_hd__or3_1
X_4553_ _4424_/X _8219_/Q _4559_/S vssd1 vssd1 vccd1 vccd1 _4554_/A sky130_fd_sc_hd__mux2_1
X_7341_ _7348_/A _7341_/B vssd1 vssd1 vccd1 vccd1 _8355_/D sky130_fd_sc_hd__nor2_1
X_4484_ _8107_/Q vssd1 vssd1 vccd1 vccd1 _4484_/X sky130_fd_sc_hd__clkbuf_2
X_7272_ _7216_/A _7272_/B _7272_/C vssd1 vssd1 vccd1 vccd1 _7272_/X sky130_fd_sc_hd__and3b_1
X_6223_ _6217_/X _8006_/Q _6219_/X _6221_/X _7795_/Q vssd1 vssd1 vccd1 vccd1 _7795_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _7731_/A vssd1 vssd1 vccd1 vccd1 _7702_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5105_ _5047_/X _5074_/X _5085_/X _5104_/X vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__a31o_2
XFILLER_85_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _7865_/Q input5/X _6092_/S vssd1 vssd1 vccd1 vccd1 _6085_/X sky130_fd_sc_hd__mux2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _6941_/C vssd1 vssd1 vccd1 vccd1 _7363_/A sky130_fd_sc_hd__inv_2
XFILLER_72_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6987_ _6987_/A vssd1 vssd1 vccd1 vccd1 _6987_/X sky130_fd_sc_hd__buf_1
X_5938_ _5938_/A vssd1 vssd1 vccd1 vccd1 _5938_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5869_ _4160_/X _7766_/Q _5869_/S vssd1 vssd1 vccd1 vccd1 _5870_/A sky130_fd_sc_hd__mux2_1
X_7608_ _6865_/A _7602_/Y _7607_/X _7568_/A vssd1 vssd1 vccd1 vccd1 _8478_/D sky130_fd_sc_hd__a211oi_1
XFILLER_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7539_ _7552_/A _7539_/B _7539_/C vssd1 vssd1 vccd1 vccd1 _7540_/A sky130_fd_sc_hd__and3_1
XFILLER_107_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput101 wbs_data_i[9] vssd1 vssd1 vccd1 vccd1 _5921_/A sky130_fd_sc_hd__buf_4
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7890_ _8063_/CLK _7890_/D vssd1 vssd1 vccd1 vccd1 _7890_/Q sky130_fd_sc_hd__dfxtp_1
X_6910_ _6910_/A vssd1 vssd1 vccd1 vccd1 _8111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6841_ _8550_/Q _7548_/S vssd1 vssd1 vccd1 vccd1 _6842_/B sky130_fd_sc_hd__xor2_1
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3984_ _5428_/A vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__buf_2
X_8511_ _8511_/CLK _8511_/D vssd1 vssd1 vccd1 vccd1 _8511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5723_ _7922_/Q _5650_/X _5725_/S vssd1 vssd1 vccd1 vccd1 _5724_/A sky130_fd_sc_hd__mux2_1
X_8442_ _8442_/CLK _8442_/D vssd1 vssd1 vccd1 vccd1 _8442_/Q sky130_fd_sc_hd__dfxtp_1
X_5654_ _5654_/A vssd1 vssd1 vccd1 vccd1 _7953_/D sky130_fd_sc_hd__clkbuf_1
X_8373_ _8373_/CLK _8373_/D vssd1 vssd1 vccd1 vccd1 _8373_/Q sky130_fd_sc_hd__dfxtp_1
X_4605_ _4620_/S vssd1 vssd1 vccd1 vccd1 _4614_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3452_ _7059_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3452_/X sky130_fd_sc_hd__clkbuf_16
X_5585_ _5585_/A vssd1 vssd1 vccd1 vccd1 _7988_/D sky130_fd_sc_hd__clkbuf_1
X_7324_ _8349_/Q _7318_/X _7310_/X _7323_/Y vssd1 vssd1 vccd1 vccd1 _7325_/B sky130_fd_sc_hd__o2bb2a_1
X_6986__445 _6986__445/A vssd1 vssd1 vccd1 vccd1 _8170_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4536_ _4536_/A vssd1 vssd1 vccd1 vccd1 _8227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4467_ _5823_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _4488_/S sky130_fd_sc_hd__nor2_2
X_7255_ _7210_/A _7210_/B _7197_/D _8355_/Q vssd1 vssd1 vccd1 vccd1 _7255_/X sky130_fd_sc_hd__a31o_1
XFILLER_104_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4398_ _4397_/X _8277_/Q _4398_/S vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__mux2_1
X_6206_ _6200_/X _7817_/Q _6202_/X _6204_/X _7785_/Q vssd1 vssd1 vccd1 vccd1 _7785_/D
+ sky130_fd_sc_hd__o32a_1
X_6137_ _7804_/Q _6122_/X _6126_/X _6135_/X _6136_/X vssd1 vssd1 vccd1 vccd1 _6137_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6068_ _7861_/Q input32/X _6072_/S vssd1 vssd1 vccd1 vccd1 _6068_/X sky130_fd_sc_hd__mux2_1
X_5019_ _4424_/X _8141_/Q _5025_/S vssd1 vssd1 vccd1 vccd1 _5020_/A sky130_fd_sc_hd__mux2_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6180__187 _6180__187/A vssd1 vssd1 vccd1 vccd1 _7774_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5370_ _4428_/X _8103_/Q _5376_/S vssd1 vssd1 vccd1 vccd1 _5371_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4321_ _4336_/S vssd1 vssd1 vccd1 vccd1 _4330_/S sky130_fd_sc_hd__buf_2
XFILLER_113_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4252_ _8336_/Q _4166_/X _4254_/S vssd1 vssd1 vccd1 vccd1 _4253_/A sky130_fd_sc_hd__mux2_1
X_7040_ _7040_/A vssd1 vssd1 vccd1 vccd1 _7040_/X sky130_fd_sc_hd__buf_1
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ _4183_/A vssd1 vssd1 vccd1 vccd1 _8392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7942_ _7942_/CLK _7942_/D vssd1 vssd1 vccd1 vccd1 _7942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7873_ _8548_/CLK _7873_/D vssd1 vssd1 vccd1 vccd1 _7873_/Q sky130_fd_sc_hd__dfxtp_1
X_6824_ _6849_/B _6824_/B vssd1 vssd1 vccd1 vccd1 _6853_/B sky130_fd_sc_hd__nand2_1
X_6755_ _6755_/A vssd1 vssd1 vccd1 vccd1 _6755_/X sky130_fd_sc_hd__buf_1
X_3967_ _8456_/Q _3966_/X _3973_/S vssd1 vssd1 vccd1 vccd1 _3968_/A sky130_fd_sc_hd__mux2_1
X_5706_ _5706_/A vssd1 vssd1 vccd1 vccd1 _7930_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3467_ clkbuf_0__3467_/X vssd1 vssd1 vccd1 vccd1 _7136__62/A sky130_fd_sc_hd__clkbuf_4
X_3898_ _3898_/A vssd1 vssd1 vccd1 vccd1 _8517_/D sky130_fd_sc_hd__clkbuf_1
X_8425_ _8425_/CLK _8425_/D vssd1 vssd1 vccd1 vccd1 _8425_/Q sky130_fd_sc_hd__dfxtp_1
X_6686_ _5950_/A _8012_/Q _6688_/S vssd1 vssd1 vccd1 vccd1 _6687_/A sky130_fd_sc_hd__mux2_1
X_5637_ _5572_/X _7959_/Q _5639_/S vssd1 vssd1 vccd1 vccd1 _5638_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5568_ _5568_/A vssd1 vssd1 vccd1 vccd1 _7993_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3435_ _6975_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3435_/X sky130_fd_sc_hd__clkbuf_16
X_8356_ _8543_/CLK _8356_/D vssd1 vssd1 vccd1 vccd1 _8356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8287_ _8287_/CLK _8287_/D vssd1 vssd1 vccd1 vccd1 _8287_/Q sky130_fd_sc_hd__dfxtp_1
X_4519_ _4519_/A vssd1 vssd1 vccd1 vccd1 _8234_/D sky130_fd_sc_hd__clkbuf_1
X_7307_ _7321_/A _7307_/B vssd1 vssd1 vccd1 vccd1 _8344_/D sky130_fd_sc_hd__nor2_1
X_5499_ _5499_/A vssd1 vssd1 vccd1 vccd1 _8046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7238_ _8345_/Q _8344_/Q _8343_/Q vssd1 vssd1 vccd1 vccd1 _7311_/A sky130_fd_sc_hd__nand3_2
XFILLER_86_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6557__250 _6557__250/A vssd1 vssd1 vccd1 vccd1 _7928_/CLK sky130_fd_sc_hd__inv_2
X_7425__145 _7425__145/A vssd1 vssd1 vccd1 vccd1 _8402_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4870_ _4787_/X _4868_/X _4869_/X vssd1 vssd1 vccd1 vccd1 _4870_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6540_ _6540_/A vssd1 vssd1 vccd1 vccd1 _6540_/X sky130_fd_sc_hd__buf_1
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3252_ clkbuf_0__3252_/X vssd1 vssd1 vccd1 vccd1 _6570__260/A sky130_fd_sc_hd__clkbuf_4
X_6471_ _6471_/A vssd1 vssd1 vccd1 vccd1 _7878_/D sky130_fd_sc_hd__clkbuf_1
X_8210_ _8210_/CLK _8210_/D vssd1 vssd1 vccd1 vccd1 _8210_/Q sky130_fd_sc_hd__dfxtp_1
X_5422_ _5379_/X _8084_/Q _5426_/S vssd1 vssd1 vccd1 vccd1 _5423_/A sky130_fd_sc_hd__mux2_1
X_8141_ _8141_/CLK _8141_/D vssd1 vssd1 vccd1 vccd1 _8141_/Q sky130_fd_sc_hd__dfxtp_1
X_5353_ _5070_/A _5348_/X _5352_/Y _5339_/X vssd1 vssd1 vccd1 vccd1 _8117_/D sky130_fd_sc_hd__o211a_1
Xoutput202 _6055_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[3] sky130_fd_sc_hd__buf_2
X_4304_ _4275_/X _8316_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__mux2_1
X_8072_ _8072_/CLK _8072_/D vssd1 vssd1 vccd1 vccd1 _8072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5284_ _7831_/Q _8428_/Q _5284_/S vssd1 vssd1 vccd1 vccd1 _5284_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_8 _5969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4235_ _8371_/Q _4169_/X _4235_/S vssd1 vssd1 vccd1 vccd1 _4236_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4166_ _8107_/Q vssd1 vssd1 vccd1 vccd1 _4166_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4097_ _4112_/S vssd1 vssd1 vccd1 vccd1 _4106_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7925_ _7925_/CLK _7925_/D vssd1 vssd1 vccd1 vccd1 _7925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7856_ _8345_/CLK _7856_/D vssd1 vssd1 vccd1 vccd1 _7856_/Q sky130_fd_sc_hd__dfxtp_1
X_6807_ _8542_/Q _7529_/B vssd1 vssd1 vccd1 vccd1 _6808_/D sky130_fd_sc_hd__xor2_1
X_4999_ _4999_/A vssd1 vssd1 vccd1 vccd1 _8150_/D sky130_fd_sc_hd__clkbuf_1
X_7787_ _8540_/CLK _7787_/D vssd1 vssd1 vccd1 vccd1 _7787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6669_ _6669_/A vssd1 vssd1 vccd1 vccd1 _8004_/D sky130_fd_sc_hd__clkbuf_1
X_8408_ _8408_/CLK _8408_/D vssd1 vssd1 vccd1 vccd1 _8408_/Q sky130_fd_sc_hd__dfxtp_1
X_8339_ _8339_/CLK _8339_/D vssd1 vssd1 vccd1 vccd1 _8339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6741__339 _6742__340/A vssd1 vssd1 vccd1 vccd1 _8049_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6999__455 _6999__455/A vssd1 vssd1 vccd1 vccd1 _8180_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8548_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4020_ _4019_/X _8439_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4021_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5971_ _5971_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5972_/A sky130_fd_sc_hd__and2_1
XFILLER_52_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7710_ _7731_/A vssd1 vssd1 vccd1 vccd1 _7710_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4922_ _4444_/X _4764_/B _4921_/X _4857_/X vssd1 vssd1 vccd1 vccd1 _8179_/D sky130_fd_sc_hd__o211a_1
X_7641_ _7641_/A vssd1 vssd1 vccd1 vccd1 _8492_/D sky130_fd_sc_hd__clkbuf_1
X_4853_ _4886_/A _4853_/B _4853_/C vssd1 vssd1 vccd1 vccd1 _4853_/X sky130_fd_sc_hd__or3_1
X_4784_ _4784_/A vssd1 vssd1 vccd1 vccd1 _4784_/X sky130_fd_sc_hd__clkbuf_2
X_7572_ _7569_/Y _7570_/X _7555_/X _7571_/Y vssd1 vssd1 vccd1 vccd1 _7573_/B sky130_fd_sc_hd__o22a_1
XFILLER_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6653__311 _6653__311/A vssd1 vssd1 vccd1 vccd1 _7997_/CLK sky130_fd_sc_hd__inv_2
X_6523_ _6523_/A vssd1 vssd1 vccd1 vccd1 _7900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6454_ _8532_/Q _6456_/B _6454_/C vssd1 vssd1 vccd1 vccd1 _6454_/X sky130_fd_sc_hd__and3_1
XFILLER_106_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5405_ _5405_/A vssd1 vssd1 vccd1 vccd1 _8092_/D sky130_fd_sc_hd__clkbuf_1
X_6385_ _8529_/Q _6356_/X _6384_/X _6350_/X _6358_/X vssd1 vssd1 vccd1 vccd1 _6385_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8124_ _8124_/CLK _8124_/D vssd1 vssd1 vccd1 vccd1 _8124_/Q sky130_fd_sc_hd__dfxtp_1
X_5336_ _5106_/A _3849_/B _7680_/B _5334_/A vssd1 vssd1 vccd1 vccd1 _5337_/C sky130_fd_sc_hd__a31o_1
XFILLER_87_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8055_ _8055_/CLK _8055_/D vssd1 vssd1 vccd1 vccd1 _8055_/Q sky130_fd_sc_hd__dfxtp_1
X_5267_ _8278_/Q _5180_/X _5207_/X _8505_/Q _5250_/X vssd1 vssd1 vccd1 vccd1 _5267_/X
+ sky130_fd_sc_hd__o221a_1
X_4218_ _5859_/A vssd1 vssd1 vccd1 vccd1 _5823_/A sky130_fd_sc_hd__buf_4
XFILLER_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3451_ clkbuf_0__3451_/X vssd1 vssd1 vccd1 vccd1 _7077_/A sky130_fd_sc_hd__clkbuf_4
X_7006_ _7006_/A vssd1 vssd1 vccd1 vccd1 _7006_/X sky130_fd_sc_hd__buf_1
X_5198_ _5319_/B vssd1 vssd1 vccd1 vccd1 _5198_/X sky130_fd_sc_hd__buf_2
X_4149_ _8402_/Q _4114_/X _4161_/S vssd1 vssd1 vccd1 vccd1 _4150_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7908_ _7908_/CLK _7908_/D vssd1 vssd1 vccd1 vccd1 _7908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7839_ _7839_/CLK _7839_/D vssd1 vssd1 vccd1 vccd1 _7839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3649_ clkbuf_0__3649_/X vssd1 vssd1 vccd1 vccd1 _7453__167/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5121_ _5055_/A _5117_/X _5120_/X vssd1 vssd1 vccd1 vccd1 _5121_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7438__155 _7438__155/A vssd1 vssd1 vccd1 vccd1 _8412_/CLK sky130_fd_sc_hd__inv_2
X_5052_ _5091_/A vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4003_ _4003_/A vssd1 vssd1 vccd1 vccd1 _8443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5954_ _5954_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__or2_4
X_5885_ _5885_/A vssd1 vssd1 vccd1 vccd1 _5885_/X sky130_fd_sc_hd__clkbuf_1
X_4905_ _4949_/B _4894_/Y _4897_/Y _4904_/X vssd1 vssd1 vccd1 vccd1 _4920_/A sky130_fd_sc_hd__a31o_1
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4836_ _7848_/Q _7773_/Q _4868_/S vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__mux2_1
X_7624_ _8485_/Q _7613_/X _7623_/X _7543_/X vssd1 vssd1 vccd1 vccd1 _8484_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7555_ _7575_/A vssd1 vssd1 vccd1 vccd1 _7555_/X sky130_fd_sc_hd__clkbuf_2
X_4767_ _4767_/A _8168_/Q vssd1 vssd1 vccd1 vccd1 _4797_/A sky130_fd_sc_hd__or2_2
X_6506_ _6506_/A vssd1 vssd1 vccd1 vccd1 _7894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4698_ _8377_/Q _8267_/Q _7980_/Q _8401_/Q _4666_/X _4667_/X vssd1 vssd1 vccd1 vccd1
+ _4698_/X sky130_fd_sc_hd__mux4_2
XFILLER_105_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6437_ _6437_/A vssd1 vssd1 vccd1 vccd1 _6437_/X sky130_fd_sc_hd__clkbuf_2
X_6368_ _6331_/X _6363_/X _6366_/X _6367_/X vssd1 vssd1 vccd1 vccd1 _6368_/X sky130_fd_sc_hd__a31o_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5319_ _8435_/Q _5319_/B vssd1 vssd1 vccd1 vccd1 _5319_/X sky130_fd_sc_hd__or2_1
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8107_ _8480_/CLK _8107_/D vssd1 vssd1 vccd1 vccd1 _8107_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8038_ _8038_/CLK _8038_/D vssd1 vssd1 vccd1 vccd1 _8038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3434_ clkbuf_0__3434_/X vssd1 vssd1 vccd1 vccd1 _6973__434/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7109__541 _7109__541/A vssd1 vssd1 vccd1 vccd1 _8268_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5670_ _5670_/A vssd1 vssd1 vccd1 vccd1 _7946_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4621_ _4621_/A vssd1 vssd1 vccd1 vccd1 _8189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4552_ _4552_/A vssd1 vssd1 vccd1 vccd1 _8220_/D sky130_fd_sc_hd__clkbuf_1
X_7340_ _8355_/Q _7334_/X _7310_/A _7258_/B vssd1 vssd1 vccd1 vccd1 _7341_/B sky130_fd_sc_hd__o2bb2a_1
X_4483_ _4483_/A vssd1 vssd1 vccd1 vccd1 _8247_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7271_ _7298_/A vssd1 vssd1 vccd1 vccd1 _7271_/Y sky130_fd_sc_hd__inv_2
X_6222_ _6217_/X _8005_/Q _6219_/X _6221_/X _7794_/Q vssd1 vssd1 vccd1 vccd1 _7794_/D
+ sky130_fd_sc_hd__o32a_1
X_7123__51 _7124__52/A vssd1 vssd1 vccd1 vccd1 _8278_/CLK sky130_fd_sc_hd__inv_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _7876_/Q _6153_/B vssd1 vssd1 vccd1 vccd1 _6153_/X sky130_fd_sc_hd__or2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5104_ _5090_/X _5094_/X _5101_/X _5206_/A _5177_/A vssd1 vssd1 vccd1 vccd1 _5104_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6075_/X _6080_/X _6081_/X _6083_/X vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__o211a_1
XFILLER_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5035_/A _5035_/B _5034_/X vssd1 vssd1 vccd1 vccd1 _6941_/C sky130_fd_sc_hd__or3b_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5937_ _5937_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5938_/A sky130_fd_sc_hd__or2_1
X_7467__3 _7469__5/A vssd1 vssd1 vccd1 vccd1 _8435_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5868_ _5868_/A vssd1 vssd1 vccd1 vccd1 _7767_/D sky130_fd_sc_hd__clkbuf_1
X_7607_ _7601_/X _6867_/C _7597_/X _7606_/X vssd1 vssd1 vccd1 vccd1 _7607_/X sky130_fd_sc_hd__o211a_1
X_5799_ _7840_/Q _4292_/A _5803_/S vssd1 vssd1 vccd1 vccd1 _5800_/A sky130_fd_sc_hd__mux2_1
X_4819_ _8154_/Q _4784_/A _4818_/X _4786_/A vssd1 vssd1 vccd1 vccd1 _4819_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7538_ _8460_/Q _7535_/X _7504_/X _7550_/C vssd1 vssd1 vccd1 vccd1 _7539_/C sky130_fd_sc_hd__o211ai_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6551__245 _6551__245/A vssd1 vssd1 vccd1 vccd1 _7923_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7665__41 _7666__42/A vssd1 vssd1 vccd1 vccd1 _8510_/CLK sky130_fd_sc_hd__inv_2
Xinput102 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _6248_/A sky130_fd_sc_hd__buf_6
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6840_ _8461_/Q vssd1 vssd1 vccd1 vccd1 _7548_/S sky130_fd_sc_hd__buf_2
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3983_ _3983_/A vssd1 vssd1 vccd1 vccd1 _8451_/D sky130_fd_sc_hd__clkbuf_1
X_8510_ _8510_/CLK _8510_/D vssd1 vssd1 vccd1 vccd1 _8510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5722_ _5722_/A vssd1 vssd1 vccd1 vccd1 _7923_/D sky130_fd_sc_hd__clkbuf_1
X_8441_ _8441_/CLK _8441_/D vssd1 vssd1 vccd1 vccd1 _8441_/Q sky130_fd_sc_hd__dfxtp_1
X_5653_ _7953_/Q _5590_/X _5653_/S vssd1 vssd1 vccd1 vccd1 _5654_/A sky130_fd_sc_hd__mux2_1
X_8372_ _8372_/CLK _8372_/D vssd1 vssd1 vccd1 vccd1 _8372_/Q sky130_fd_sc_hd__dfxtp_1
X_5584_ _7988_/Q _5583_/X _5591_/S vssd1 vssd1 vccd1 vccd1 _5585_/A sky130_fd_sc_hd__mux2_1
X_4604_ _4604_/A _5482_/A vssd1 vssd1 vccd1 vccd1 _4620_/S sky130_fd_sc_hd__nor2_2
Xclkbuf_0__3451_ _7058_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3451_/X sky130_fd_sc_hd__clkbuf_16
X_4535_ _4379_/X _8227_/Q _4541_/S vssd1 vssd1 vccd1 vccd1 _4536_/A sky130_fd_sc_hd__mux2_1
X_7323_ _7323_/A _7323_/B vssd1 vssd1 vccd1 vccd1 _7323_/Y sky130_fd_sc_hd__nand2_1
X_4466_ _5622_/A _4466_/B _4933_/C vssd1 vssd1 vccd1 vccd1 _5679_/B sky130_fd_sc_hd__or3_4
X_7254_ _8540_/Q _7254_/B vssd1 vssd1 vccd1 vccd1 _7277_/B sky130_fd_sc_hd__xor2_1
XFILLER_89_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4397_ _8488_/Q vssd1 vssd1 vccd1 vccd1 _4397_/X sky130_fd_sc_hd__clkbuf_2
X_6205_ _6200_/X _7816_/Q _6202_/X _6204_/X _7784_/Q vssd1 vssd1 vccd1 vccd1 _7784_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_98_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6136_ _7633_/C vssd1 vssd1 vccd1 vccd1 _6136_/X sky130_fd_sc_hd__clkbuf_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6067_ _6056_/X _6065_/X _6066_/X _6063_/X vssd1 vssd1 vccd1 vccd1 _6067_/X sky130_fd_sc_hd__o211a_1
X_5018_ _5018_/A vssd1 vssd1 vccd1 vccd1 _8142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6969_ _6987_/A vssd1 vssd1 vccd1 vccd1 _6969_/X sky130_fd_sc_hd__buf_1
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3649_ _7451_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3649_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6870__370 _6870__370/A vssd1 vssd1 vccd1 vccd1 _8084_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4320_ _4567_/A _4356_/B vssd1 vssd1 vccd1 vccd1 _4336_/S sky130_fd_sc_hd__or2_2
X_4251_ _4251_/A vssd1 vssd1 vccd1 vccd1 _8337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4182_ _8392_/Q _4181_/X _4188_/S vssd1 vssd1 vccd1 vccd1 _4183_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7941_ _7941_/CLK _7941_/D vssd1 vssd1 vccd1 vccd1 _7941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7872_ _8548_/CLK _7872_/D vssd1 vssd1 vccd1 vccd1 _7872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6823_ _8545_/Q _7571_/A _7571_/B vssd1 vssd1 vccd1 vccd1 _6823_/X sky130_fd_sc_hd__and3_1
X_6992__450 _6992__450/A vssd1 vssd1 vccd1 vccd1 _8175_/CLK sky130_fd_sc_hd__inv_2
X_3966_ _8493_/Q vssd1 vssd1 vccd1 vccd1 _3966_/X sky130_fd_sc_hd__buf_4
X_5705_ _7930_/Q _5650_/X _5707_/S vssd1 vssd1 vccd1 vccd1 _5706_/A sky130_fd_sc_hd__mux2_1
X_7088__525 _7088__525/A vssd1 vssd1 vccd1 vccd1 _8252_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3466_ clkbuf_0__3466_/X vssd1 vssd1 vccd1 vccd1 _7130__57/A sky130_fd_sc_hd__clkbuf_4
X_6685_ _6685_/A vssd1 vssd1 vccd1 vccd1 _8011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5636_ _5636_/A vssd1 vssd1 vccd1 vccd1 _7960_/D sky130_fd_sc_hd__clkbuf_1
X_3897_ _3896_/X _8517_/Q _3903_/S vssd1 vssd1 vccd1 vccd1 _3898_/A sky130_fd_sc_hd__mux2_1
X_8424_ _8424_/CLK _8424_/D vssd1 vssd1 vccd1 vccd1 _8424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5567_ _5566_/X _7993_/Q _5567_/S vssd1 vssd1 vccd1 vccd1 _5568_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3434_ _6969_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3434_/X sky130_fd_sc_hd__clkbuf_16
X_8355_ _8355_/CLK _8355_/D vssd1 vssd1 vccd1 vccd1 _8355_/Q sky130_fd_sc_hd__dfxtp_1
X_5498_ _8046_/Q _4298_/A _5498_/S vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__mux2_1
X_8286_ _8286_/CLK _8286_/D vssd1 vssd1 vccd1 vccd1 _8286_/Q sky130_fd_sc_hd__dfxtp_1
X_4518_ _8234_/Q _4517_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4519_/A sky130_fd_sc_hd__mux2_1
X_7306_ _7299_/B _7246_/B _7303_/Y _7301_/X _8344_/Q vssd1 vssd1 vccd1 vccd1 _7307_/B
+ sky130_fd_sc_hd__a32oi_1
XFILLER_78_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4449_ _4374_/X _8260_/Q _4457_/S vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__mux2_1
X_7237_ _8547_/Q _7237_/B vssd1 vssd1 vccd1 vccd1 _7281_/C sky130_fd_sc_hd__xor2_1
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _7799_/Q _6122_/A vssd1 vssd1 vccd1 vccd1 _6119_/X sky130_fd_sc_hd__or2_1
XFILLER_39_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7484__17 _7485__18/A vssd1 vssd1 vccd1 vccd1 _8449_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6564__255 _6564__255/A vssd1 vssd1 vccd1 vccd1 _7933_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3320_ clkbuf_0__3320_/X vssd1 vssd1 vccd1 vccd1 _6779__365/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3251_ clkbuf_0__3251_/X vssd1 vssd1 vccd1 vccd1 _6563__254/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7157__79 _7158__80/A vssd1 vssd1 vccd1 vccd1 _8306_/CLK sky130_fd_sc_hd__inv_2
X_6470_ _5978_/A _7878_/Q _6476_/S vssd1 vssd1 vccd1 vccd1 _6471_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5421_ _5421_/A vssd1 vssd1 vccd1 vccd1 _8085_/D sky130_fd_sc_hd__clkbuf_1
X_5352_ _5356_/A _5352_/B vssd1 vssd1 vccd1 vccd1 _5352_/Y sky130_fd_sc_hd__nand2_1
X_8140_ _8140_/CLK _8140_/D vssd1 vssd1 vccd1 vccd1 _8140_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput203 _6060_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_114_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8071_ _8071_/CLK _8071_/D vssd1 vssd1 vccd1 vccd1 _8071_/Q sky130_fd_sc_hd__dfxtp_1
X_4303_ _4318_/S vssd1 vssd1 vccd1 vccd1 _4312_/S sky130_fd_sc_hd__buf_2
X_5283_ _5356_/B _5281_/X _5282_/X vssd1 vssd1 vccd1 vccd1 _5283_/Y sky130_fd_sc_hd__o21ai_1
XINSDIODE2_9 _5947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4234_ _4234_/A vssd1 vssd1 vccd1 vccd1 _8372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4165_ _4165_/A vssd1 vssd1 vccd1 vccd1 _8397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4096_ _5787_/A _4199_/B vssd1 vssd1 vccd1 vccd1 _4112_/S sky130_fd_sc_hd__or2_2
XFILLER_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7924_ _7924_/CLK _7924_/D vssd1 vssd1 vccd1 vccd1 _7924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7855_ _8370_/CLK _7855_/D vssd1 vssd1 vccd1 vccd1 _7855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6806_ _6816_/B _6806_/B vssd1 vssd1 vccd1 vccd1 _7529_/B sky130_fd_sc_hd__nand2_2
X_4998_ _8150_/Q _4465_/X _5006_/S vssd1 vssd1 vccd1 vccd1 _4999_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6918__395 _6918__395/A vssd1 vssd1 vccd1 vccd1 _8117_/CLK sky130_fd_sc_hd__inv_2
X_7786_ _8543_/CLK _7786_/D vssd1 vssd1 vccd1 vccd1 _7786_/Q sky130_fd_sc_hd__dfxtp_1
X_8552__250 vssd1 vssd1 vccd1 vccd1 core1Index[0] _8552__250/LO sky130_fd_sc_hd__conb_1
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6737_ _6737_/A vssd1 vssd1 vccd1 vccd1 _6737_/X sky130_fd_sc_hd__buf_1
X_3949_ _3949_/A vssd1 vssd1 vccd1 vccd1 _8498_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3449_ clkbuf_0__3449_/X vssd1 vssd1 vccd1 vccd1 _7049__493/A sky130_fd_sc_hd__clkbuf_4
X_6668_ _5932_/A _8004_/Q _6670_/S vssd1 vssd1 vccd1 vccd1 _6669_/A sky130_fd_sc_hd__mux2_1
X_8407_ _8407_/CLK _8407_/D vssd1 vssd1 vccd1 vccd1 _8407_/Q sky130_fd_sc_hd__dfxtp_1
X_5619_ _5619_/A vssd1 vssd1 vccd1 vccd1 _7975_/D sky130_fd_sc_hd__clkbuf_1
X_8338_ _8338_/CLK _8338_/D vssd1 vssd1 vccd1 vccd1 _8338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8269_ _8269_/CLK _8269_/D vssd1 vssd1 vccd1 vccd1 _8269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7103__536 _7107__540/A vssd1 vssd1 vccd1 vccd1 _8263_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7431__150 _7431__150/A vssd1 vssd1 vccd1 vccd1 _8407_/CLK sky130_fd_sc_hd__inv_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5970_ _5970_/A vssd1 vssd1 vccd1 vccd1 _5970_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4921_ _4713_/A _8179_/Q _4948_/A _4920_/Y _4712_/A vssd1 vssd1 vccd1 vccd1 _4921_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4852_ _8092_/Q _4781_/A _4782_/A _4851_/X vssd1 vssd1 vccd1 vccd1 _4853_/C sky130_fd_sc_hd__o211a_1
XFILLER_21_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7640_ _7640_/A _7646_/B _7640_/C vssd1 vssd1 vccd1 vccd1 _7641_/A sky130_fd_sc_hd__and3_1
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4783_ _4783_/A vssd1 vssd1 vccd1 vccd1 _4784_/A sky130_fd_sc_hd__clkbuf_2
X_7571_ _7571_/A _7571_/B vssd1 vssd1 vccd1 vccd1 _7571_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6522_ _6522_/A _6522_/B _6522_/C vssd1 vssd1 vccd1 vccd1 _6523_/A sky130_fd_sc_hd__and3_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6453_ _7872_/Q _6442_/X _6437_/X _6452_/X _6435_/A vssd1 vssd1 vccd1 vccd1 _7872_/D
+ sky130_fd_sc_hd__a221o_1
X_5404_ _5379_/X _8092_/Q _5408_/S vssd1 vssd1 vccd1 vccd1 _5405_/A sky130_fd_sc_hd__mux2_1
X_8123_ _8123_/CLK _8123_/D vssd1 vssd1 vccd1 vccd1 _8123_/Q sky130_fd_sc_hd__dfxtp_1
X_6384_ _7741_/A _7970_/Q _6352_/X _6364_/X vssd1 vssd1 vccd1 vccd1 _6384_/X sky130_fd_sc_hd__a31o_1
X_5335_ _5335_/A vssd1 vssd1 vccd1 vccd1 _7680_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8054_ _8054_/CLK _8054_/D vssd1 vssd1 vccd1 vccd1 _8054_/Q sky130_fd_sc_hd__dfxtp_1
X_5266_ _8238_/Q _8254_/Q _5281_/S vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3450_ clkbuf_0__3450_/X vssd1 vssd1 vccd1 vccd1 _7054__497/A sky130_fd_sc_hd__clkbuf_4
X_6883__380 _6883__380/A vssd1 vssd1 vccd1 vccd1 _8094_/CLK sky130_fd_sc_hd__inv_2
X_4217_ _4217_/A _4217_/B _4931_/B vssd1 vssd1 vccd1 vccd1 _5859_/A sky130_fd_sc_hd__or3_4
X_5197_ _5197_/A vssd1 vssd1 vccd1 vccd1 _5319_/B sky130_fd_sc_hd__clkbuf_2
X_4148_ _4170_/S vssd1 vssd1 vccd1 vccd1 _4161_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _4094_/S vssd1 vssd1 vccd1 vccd1 _4088_/S sky130_fd_sc_hd__buf_2
XFILLER_71_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7907_ _7907_/CLK _7907_/D vssd1 vssd1 vccd1 vccd1 _7907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7838_ _7838_/CLK _7838_/D vssd1 vssd1 vccd1 vccd1 _7838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7769_ _7769_/CLK _7769_/D vssd1 vssd1 vccd1 vccd1 _7769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3648_ clkbuf_0__3648_/X vssd1 vssd1 vccd1 vccd1 _7450__165/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6717__320 _6717__320/A vssd1 vssd1 vccd1 vccd1 _8030_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5120_ _5079_/X _5119_/X _5235_/A vssd1 vssd1 vccd1 vccd1 _5120_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7150__74 _7151__75/A vssd1 vssd1 vccd1 vccd1 _8301_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5051_ _5070_/B _5063_/B vssd1 vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__nor2_1
X_4002_ _3911_/X _8443_/Q _4002_/S vssd1 vssd1 vccd1 vccd1 _4003_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _5953_/A vssd1 vssd1 vccd1 vccd1 _5953_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5884_ _6465_/A _5890_/B vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__and2_1
X_4904_ _4638_/A _4900_/Y _4903_/Y _4670_/X vssd1 vssd1 vccd1 vccd1 _4904_/X sky130_fd_sc_hd__a31o_1
X_4835_ _7824_/Q _4791_/X _4809_/A _4834_/X vssd1 vssd1 vccd1 vccd1 _4835_/X sky130_fd_sc_hd__o22a_1
X_7623_ _8484_/Q _7614_/X vssd1 vssd1 vccd1 vccd1 _7623_/X sky130_fd_sc_hd__or2b_1
XFILLER_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4766_ _4767_/A _4766_/B vssd1 vssd1 vccd1 vccd1 _4768_/A sky130_fd_sc_hd__nand2_2
X_7554_ _8463_/Q vssd1 vssd1 vccd1 vccd1 _7554_/Y sky130_fd_sc_hd__inv_2
X_6505_ _8009_/Q _7894_/Q _6509_/S vssd1 vssd1 vccd1 vccd1 _6506_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4697_ _8219_/Q _8203_/Q _8165_/Q _8235_/Q _4810_/S _4649_/X vssd1 vssd1 vccd1 vccd1
+ _4697_/X sky130_fd_sc_hd__mux4_1
X_6436_ _7867_/Q _6424_/X _6415_/X _6434_/X _6435_/X vssd1 vssd1 vccd1 vccd1 _7867_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6367_ _6367_/A vssd1 vssd1 vccd1 vccd1 _6367_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5318_ _7830_/Q _8427_/Q _5318_/S vssd1 vssd1 vccd1 vccd1 _5318_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8106_ _8480_/CLK _8106_/D vssd1 vssd1 vccd1 vccd1 _8106_/Q sky130_fd_sc_hd__dfxtp_4
X_6298_ _6310_/A vssd1 vssd1 vccd1 vccd1 _6298_/X sky130_fd_sc_hd__buf_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8037_ _8037_/CLK _8037_/D vssd1 vssd1 vccd1 vccd1 _8037_/Q sky130_fd_sc_hd__dfxtp_1
X_5249_ _8498_/Q _5232_/X _5198_/X _8514_/Q vssd1 vssd1 vccd1 vccd1 _5249_/X sky130_fd_sc_hd__o22a_1
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _8551_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3433_ clkbuf_0__3433_/X vssd1 vssd1 vccd1 vccd1 _6968__430/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _8189_/Q _4196_/X _4620_/S vssd1 vssd1 vccd1 vccd1 _4621_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7444__160 _7444__160/A vssd1 vssd1 vccd1 vccd1 _8417_/CLK sky130_fd_sc_hd__inv_2
X_4551_ _4418_/X _8220_/Q _4559_/S vssd1 vssd1 vccd1 vccd1 _4552_/A sky130_fd_sc_hd__mux2_1
X_4482_ _8247_/Q _4481_/X _4488_/S vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__mux2_1
X_7270_ _7270_/A vssd1 vssd1 vccd1 vccd1 _8333_/D sky130_fd_sc_hd__clkbuf_1
X_6221_ _6239_/A vssd1 vssd1 vccd1 vccd1 _6221_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6152_ _7810_/Q _7633_/A _6139_/A _6151_/X _6063_/A vssd1 vssd1 vccd1 vccd1 _6152_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5103_ _8118_/Q _5103_/B vssd1 vssd1 vccd1 vccd1 _5177_/A sky130_fd_sc_hd__xnor2_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _7633_/C vssd1 vssd1 vccd1 vccd1 _6083_/X sky130_fd_sc_hd__clkbuf_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5034_/A _5034_/B _5034_/C _5034_/D vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__and4_1
XFILLER_93_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6956__421 _6957__422/A vssd1 vssd1 vccd1 vccd1 _8145_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5936_ _5936_/A vssd1 vssd1 vccd1 vccd1 _5936_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5867_ _4157_/X _7767_/Q _5869_/S vssd1 vssd1 vccd1 vccd1 _5868_/A sky130_fd_sc_hd__mux2_1
X_7606_ _7609_/A _7606_/B _7606_/C vssd1 vssd1 vccd1 vccd1 _7606_/X sky130_fd_sc_hd__or3_1
X_5798_ _5798_/A vssd1 vssd1 vccd1 vccd1 _7841_/D sky130_fd_sc_hd__clkbuf_1
X_4818_ _7913_/Q _8085_/Q _4880_/S vssd1 vssd1 vccd1 vccd1 _4818_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4749_ _4953_/B _4746_/X _4748_/X vssd1 vssd1 vccd1 vccd1 _4749_/X sky130_fd_sc_hd__a21o_1
X_7537_ _7504_/X _7575_/A _7550_/C vssd1 vssd1 vccd1 vccd1 _7539_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6419_ _8063_/Q vssd1 vssd1 vccd1 vccd1 _6431_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput103 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _6654_/A sky130_fd_sc_hd__buf_6
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8595__242 vssd1 vssd1 vccd1 vccd1 _8595__242/HI partID[7] sky130_fd_sc_hd__conb_1
XFILLER_72_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7387__114 _7388__115/A vssd1 vssd1 vccd1 vccd1 _8371_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3982_ _8451_/Q _3981_/X _3982_/S vssd1 vssd1 vccd1 vccd1 _3983_/A sky130_fd_sc_hd__mux2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5721_ _7923_/Q _5647_/X _5725_/S vssd1 vssd1 vccd1 vccd1 _5722_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8440_ _8440_/CLK _8440_/D vssd1 vssd1 vccd1 vccd1 _8440_/Q sky130_fd_sc_hd__dfxtp_1
X_5652_ _5652_/A vssd1 vssd1 vccd1 vccd1 _7954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8371_ _8371_/CLK _8371_/D vssd1 vssd1 vccd1 vccd1 _8371_/Q sky130_fd_sc_hd__dfxtp_1
X_4603_ _4603_/A vssd1 vssd1 vccd1 vccd1 _8197_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3450_ _7052_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3450_/X sky130_fd_sc_hd__clkbuf_16
X_5583_ _8112_/Q vssd1 vssd1 vccd1 vccd1 _5583_/X sky130_fd_sc_hd__buf_4
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4534_ _4534_/A vssd1 vssd1 vccd1 vccd1 _8228_/D sky130_fd_sc_hd__clkbuf_1
X_7322_ _7360_/B vssd1 vssd1 vccd1 vccd1 _7336_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7253_ _7210_/A _7210_/B _7197_/D _7220_/A _7252_/Y vssd1 vssd1 vccd1 vccd1 _7254_/B
+ sky130_fd_sc_hd__a32o_1
X_4465_ _8113_/Q vssd1 vssd1 vccd1 vccd1 _4465_/X sky130_fd_sc_hd__buf_4
XFILLER_116_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7184_ _7395_/A vssd1 vssd1 vccd1 vccd1 _7184_/X sky130_fd_sc_hd__buf_1
X_4396_ _4396_/A vssd1 vssd1 vccd1 vccd1 _8278_/D sky130_fd_sc_hd__clkbuf_1
X_6204_ _6213_/A vssd1 vssd1 vccd1 vccd1 _6204_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6135_ _6135_/A _6140_/B vssd1 vssd1 vccd1 vccd1 _6135_/X sky130_fd_sc_hd__and2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6066_ _7785_/Q _6066_/B vssd1 vssd1 vccd1 vccd1 _6066_/X sky130_fd_sc_hd__or2_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _4418_/X _8142_/Q _5025_/S vssd1 vssd1 vccd1 vccd1 _5018_/A sky130_fd_sc_hd__mux2_1
X_8579__226 vssd1 vssd1 vccd1 vccd1 _8579__226/HI core1Index[6] sky130_fd_sc_hd__conb_1
XFILLER_54_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5919_ _5919_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5920_/A sky130_fd_sc_hd__or2_1
XFILLER_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6899_ _6899_/A vssd1 vssd1 vccd1 vccd1 _8106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3648_ _7445_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3648_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_108_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7496__26 _7650__29/A vssd1 vssd1 vccd1 vccd1 _8458_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4250_ _8337_/Q _4163_/X _4254_/S vssd1 vssd1 vccd1 vccd1 _4251_/A sky130_fd_sc_hd__mux2_1
X_4181_ _8493_/Q vssd1 vssd1 vccd1 vccd1 _4181_/X sky130_fd_sc_hd__buf_2
X_7940_ _7940_/CLK _7940_/D vssd1 vssd1 vccd1 vccd1 _7940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7871_ _8548_/CLK _7871_/D vssd1 vssd1 vccd1 vccd1 _7871_/Q sky130_fd_sc_hd__dfxtp_1
X_6822_ _7571_/A _7571_/B _8545_/Q vssd1 vssd1 vccd1 vccd1 _6822_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3965_ _3965_/A vssd1 vssd1 vccd1 vccd1 _8457_/D sky130_fd_sc_hd__clkbuf_1
X_5704_ _5704_/A vssd1 vssd1 vccd1 vccd1 _7931_/D sky130_fd_sc_hd__clkbuf_1
X_7053__496 _7054__497/A vssd1 vssd1 vccd1 vccd1 _8223_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3465_ clkbuf_0__3465_/X vssd1 vssd1 vccd1 vccd1 _7124__52/A sky130_fd_sc_hd__clkbuf_4
X_3896_ _8493_/Q vssd1 vssd1 vccd1 vccd1 _3896_/X sky130_fd_sc_hd__buf_4
X_6684_ _5948_/A _8011_/Q _6688_/S vssd1 vssd1 vccd1 vccd1 _6685_/A sky130_fd_sc_hd__mux2_1
X_5635_ _5569_/X _7960_/Q _5639_/S vssd1 vssd1 vccd1 vccd1 _5636_/A sky130_fd_sc_hd__mux2_1
X_8423_ _8423_/CLK _8423_/D vssd1 vssd1 vccd1 vccd1 _8423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3433_ _6963_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3433_/X sky130_fd_sc_hd__clkbuf_16
X_5566_ _5566_/A vssd1 vssd1 vccd1 vccd1 _5566_/X sky130_fd_sc_hd__buf_2
X_8354_ _8355_/CLK _8354_/D vssd1 vssd1 vccd1 vccd1 _8354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5497_ _5497_/A vssd1 vssd1 vccd1 vccd1 _8047_/D sky130_fd_sc_hd__clkbuf_1
X_8285_ _8285_/CLK _8285_/D vssd1 vssd1 vccd1 vccd1 _8285_/Q sky130_fd_sc_hd__dfxtp_1
X_7305_ _7360_/B vssd1 vssd1 vccd1 vccd1 _7321_/A sky130_fd_sc_hd__clkbuf_2
X_4517_ _8111_/Q vssd1 vssd1 vccd1 vccd1 _4517_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_104_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4448_ _4463_/S vssd1 vssd1 vccd1 vccd1 _4457_/S sky130_fd_sc_hd__clkbuf_2
X_7236_ _7236_/A _7236_/B vssd1 vssd1 vccd1 vccd1 _7237_/B sky130_fd_sc_hd__xnor2_1
X_6290__195 _6290__195/A vssd1 vssd1 vccd1 vccd1 _7825_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4379_ _8494_/Q vssd1 vssd1 vccd1 vccd1 _4379_/X sky130_fd_sc_hd__buf_2
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _7874_/Q input15/X _6153_/B vssd1 vssd1 vccd1 vccd1 _6118_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6049_ _7856_/Q input25/X _6123_/B vssd1 vssd1 vccd1 vccd1 _6049_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6711__315 _6711__315/A vssd1 vssd1 vccd1 vccd1 _8025_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3250_ clkbuf_0__3250_/X vssd1 vssd1 vccd1 vccd1 _6571_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5420_ _5375_/X _8085_/Q _5420_/S vssd1 vssd1 vccd1 vccd1 _5421_/A sky130_fd_sc_hd__mux2_1
X_5351_ _8118_/Q _5348_/X _5350_/Y _5339_/X vssd1 vssd1 vccd1 vccd1 _8118_/D sky130_fd_sc_hd__o211a_1
Xoutput204 _6064_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_114_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8070_ _8070_/CLK _8070_/D vssd1 vssd1 vccd1 vccd1 _8070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5282_ _8412_/Q _5270_/X _5239_/X _8404_/Q _5205_/S vssd1 vssd1 vccd1 vccd1 _5282_/X
+ sky130_fd_sc_hd__o221a_1
X_4302_ _4531_/A _4356_/B vssd1 vssd1 vccd1 vccd1 _4318_/S sky130_fd_sc_hd__or2_2
X_4233_ _8372_/Q _4166_/X _4235_/S vssd1 vssd1 vccd1 vccd1 _4234_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7021_ _7021_/A vssd1 vssd1 vccd1 vccd1 _7021_/X sky130_fd_sc_hd__buf_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4164_ _8397_/Q _4163_/X _4170_/S vssd1 vssd1 vccd1 vccd1 _4165_/A sky130_fd_sc_hd__mux2_1
X_4095_ _4095_/A vssd1 vssd1 vccd1 vccd1 _8411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7923_ _7923_/CLK _7923_/D vssd1 vssd1 vccd1 vccd1 _7923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7854_ _8370_/CLK _7854_/D vssd1 vssd1 vccd1 vccd1 _7854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6805_ _8469_/Q _6830_/A _6824_/B _8470_/Q vssd1 vssd1 vccd1 vccd1 _6806_/B sky130_fd_sc_hd__a31o_1
X_7785_ _8543_/CLK _7785_/D vssd1 vssd1 vccd1 vccd1 _7785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4997_ _5012_/S vssd1 vssd1 vccd1 vccd1 _5006_/S sky130_fd_sc_hd__buf_2
X_3948_ _3905_/X _8498_/Q _3952_/S vssd1 vssd1 vccd1 vccd1 _3949_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3448_ clkbuf_0__3448_/X vssd1 vssd1 vccd1 vccd1 _7043__488/A sky130_fd_sc_hd__clkbuf_4
X_6667_ _6667_/A vssd1 vssd1 vccd1 vccd1 _8003_/D sky130_fd_sc_hd__clkbuf_1
X_3879_ _7900_/Q _7899_/Q vssd1 vssd1 vccd1 vccd1 _7696_/A sky130_fd_sc_hd__nor2_2
X_8406_ _8406_/CLK _8406_/D vssd1 vssd1 vccd1 vccd1 _8406_/Q sky130_fd_sc_hd__dfxtp_1
X_5618_ _5572_/X _7975_/Q _5620_/S vssd1 vssd1 vccd1 vccd1 _5619_/A sky130_fd_sc_hd__mux2_1
X_8337_ _8337_/CLK _8337_/D vssd1 vssd1 vccd1 vccd1 _8337_/Q sky130_fd_sc_hd__dfxtp_1
X_5549_ _5549_/A vssd1 vssd1 vccd1 vccd1 _8024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8268_ _8268_/CLK _8268_/D vssd1 vssd1 vccd1 vccd1 _8268_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8199_ _8199_/CLK _8199_/D vssd1 vssd1 vccd1 vccd1 _8199_/Q sky130_fd_sc_hd__dfxtp_1
X_7219_ _7210_/A _7210_/B _7218_/D _8353_/Q vssd1 vssd1 vccd1 vccd1 _7220_/B sky130_fd_sc_hd__a31o_1
XFILLER_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6570__260 _6570__260/A vssd1 vssd1 vccd1 vccd1 _7938_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7162__83 _7163__84/A vssd1 vssd1 vccd1 vccd1 _8310_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ _4920_/A _4920_/B vssd1 vssd1 vccd1 vccd1 _4920_/Y sky130_fd_sc_hd__nand2_2
X_4851_ _8153_/Q _4784_/A _4850_/X _4786_/A vssd1 vssd1 vccd1 vccd1 _4851_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4782_ _4782_/A vssd1 vssd1 vccd1 vccd1 _4782_/X sky130_fd_sc_hd__clkbuf_2
X_6950__416 _6952__418/A vssd1 vssd1 vccd1 vccd1 _8140_/CLK sky130_fd_sc_hd__inv_2
X_7570_ _7588_/A vssd1 vssd1 vccd1 vccd1 _7570_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6521_ _6521_/A _6521_/B _6521_/C vssd1 vssd1 vccd1 vccd1 _6522_/C sky130_fd_sc_hd__or3_1
X_6452_ _8533_/Q _6452_/B _6454_/C vssd1 vssd1 vccd1 vccd1 _6452_/X sky130_fd_sc_hd__and3_1
X_5403_ _5403_/A vssd1 vssd1 vccd1 vccd1 _8093_/D sky130_fd_sc_hd__clkbuf_1
X_6317__216 _6318__217/A vssd1 vssd1 vccd1 vccd1 _7846_/CLK sky130_fd_sc_hd__inv_2
X_6383_ _8547_/Q _6362_/X _6410_/C _6343_/X vssd1 vssd1 vccd1 vccd1 _6383_/X sky130_fd_sc_hd__a31o_1
X_8122_ _8122_/CLK _8122_/D vssd1 vssd1 vccd1 vccd1 _8122_/Q sky130_fd_sc_hd__dfxtp_1
X_5334_ _5334_/A _5334_/B _5334_/C vssd1 vssd1 vccd1 vccd1 _5337_/B sky130_fd_sc_hd__nand3_1
X_8053_ _8053_/CLK _8053_/D vssd1 vssd1 vccd1 vccd1 _8053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5265_ _5305_/S vssd1 vssd1 vccd1 vccd1 _5281_/S sky130_fd_sc_hd__buf_4
X_4216_ _4216_/A vssd1 vssd1 vccd1 vccd1 _8379_/D sky130_fd_sc_hd__clkbuf_1
X_5196_ _5227_/A vssd1 vssd1 vccd1 vccd1 _5196_/X sky130_fd_sc_hd__buf_2
XFILLER_87_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4147_ _5602_/A _5641_/A vssd1 vssd1 vccd1 vccd1 _4170_/S sky130_fd_sc_hd__nor2_2
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4078_ _4531_/A _4199_/B vssd1 vssd1 vccd1 vccd1 _4094_/S sky130_fd_sc_hd__or2_2
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7906_ _7906_/CLK _7906_/D vssd1 vssd1 vccd1 vccd1 _7906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7837_ _7837_/CLK _7837_/D vssd1 vssd1 vccd1 vccd1 _7837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7768_ _7768_/CLK _7768_/D vssd1 vssd1 vccd1 vccd1 _7768_/Q sky130_fd_sc_hd__dfxtp_1
X_7699_ _8064_/Q _7747_/B vssd1 vssd1 vccd1 vccd1 _7700_/A sky130_fd_sc_hd__and2_1
XFILLER_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3647_ clkbuf_0__3647_/X vssd1 vssd1 vccd1 vccd1 _7441__157/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8559__257 vssd1 vssd1 vccd1 vccd1 partID[11] _8559__257/LO sky130_fd_sc_hd__conb_1
XFILLER_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7135__61 _7136__62/A vssd1 vssd1 vccd1 vccd1 _8288_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _5181_/A _5182_/B _8116_/Q vssd1 vssd1 vccd1 vccd1 _5063_/B sky130_fd_sc_hd__a21oi_4
X_4001_ _4001_/A vssd1 vssd1 vccd1 vccd1 _8444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5952_ _5952_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _5953_/A sky130_fd_sc_hd__or2_4
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4903_ _4803_/X _4901_/X _4902_/X vssd1 vssd1 vccd1 vccd1 _4903_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5883_ _6021_/A vssd1 vssd1 vccd1 vccd1 _5890_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4834_ _7960_/Q _7944_/Q _4866_/S vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__mux2_1
X_7622_ _8484_/Q _7613_/X _7621_/X _7552_/X vssd1 vssd1 vccd1 vccd1 _8483_/D sky130_fd_sc_hd__o211a_1
X_7553_ _7550_/X _7551_/X _7552_/X vssd1 vssd1 vccd1 vccd1 _8462_/D sky130_fd_sc_hd__o21a_1
X_4765_ _4712_/X _4763_/X _4764_/X _4690_/X vssd1 vssd1 vccd1 vccd1 _8183_/D sky130_fd_sc_hd__o211a_1
X_6504_ _6504_/A vssd1 vssd1 vccd1 vccd1 _7893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4696_ _4714_/A _4692_/X _4695_/X vssd1 vssd1 vccd1 vccd1 _4696_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6435_ _6435_/A vssd1 vssd1 vccd1 vccd1 _6435_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6366_ _8526_/Q _6356_/X _6365_/X _6350_/X _6358_/X vssd1 vssd1 vccd1 vccd1 _6366_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5317_ _5193_/X _5315_/X _5316_/X vssd1 vssd1 vccd1 vccd1 _5317_/X sky130_fd_sc_hd__o21a_1
X_8105_ _8105_/CLK _8105_/D vssd1 vssd1 vccd1 vccd1 _8105_/Q sky130_fd_sc_hd__dfxtp_1
X_6297_ _6297_/A vssd1 vssd1 vccd1 vccd1 _6297_/X sky130_fd_sc_hd__buf_1
X_8036_ _8036_/CLK _8036_/D vssd1 vssd1 vccd1 vccd1 _8036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5248_ _8040_/Q _8067_/Q _5312_/S vssd1 vssd1 vccd1 vccd1 _5248_/X sky130_fd_sc_hd__mux2_1
X_5179_ _5227_/A vssd1 vssd1 vccd1 vccd1 _5232_/A sky130_fd_sc_hd__inv_2
XFILLER_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3432_ clkbuf_0__3432_/X vssd1 vssd1 vccd1 vccd1 _6987_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7116__547 _7118__549/A vssd1 vssd1 vccd1 vccd1 _8274_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4550_ _4565_/S vssd1 vssd1 vccd1 vccd1 _4559_/S sky130_fd_sc_hd__buf_2
X_4481_ _8108_/Q vssd1 vssd1 vccd1 vccd1 _4481_/X sky130_fd_sc_hd__buf_2
XFILLER_7_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6220_ _6217_/X _8004_/Q _6219_/X _6213_/X _7793_/Q vssd1 vssd1 vccd1 vccd1 _7793_/D
+ sky130_fd_sc_hd__o32a_1
X_6151_ _6151_/A _6151_/B vssd1 vssd1 vccd1 vccd1 _6151_/X sky130_fd_sc_hd__and2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5102_ _5258_/A vssd1 vssd1 vccd1 vccd1 _5206_/A sky130_fd_sc_hd__clkbuf_2
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6082_/A vssd1 vssd1 vccd1 vccd1 _7633_/C sky130_fd_sc_hd__buf_4
XFILLER_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _8133_/Q vssd1 vssd1 vccd1 vccd1 _5106_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5935_ _5935_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__or2_1
X_5866_ _5866_/A vssd1 vssd1 vccd1 vccd1 _7768_/D sky130_fd_sc_hd__clkbuf_1
X_7017__467 _7020__470/A vssd1 vssd1 vccd1 vccd1 _8194_/CLK sky130_fd_sc_hd__inv_2
X_4817_ _4803_/A _4815_/X _4816_/X vssd1 vssd1 vccd1 vccd1 _4821_/B sky130_fd_sc_hd__o21a_1
X_7605_ _8478_/Q _8477_/Q vssd1 vssd1 vccd1 vccd1 _7606_/C sky130_fd_sc_hd__nor2_1
X_5797_ _7841_/Q _4289_/A _5797_/S vssd1 vssd1 vccd1 vccd1 _5798_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4748_ _4664_/X _4747_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _4748_/X sky130_fd_sc_hd__a21o_1
X_7536_ _6860_/X _7609_/A _7505_/Y _7535_/X vssd1 vssd1 vccd1 vccd1 _7575_/A sky130_fd_sc_hd__o22a_1
XFILLER_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4679_ _7829_/Q _7949_/Q _7965_/Q _7933_/Q _4876_/A _4649_/A vssd1 vssd1 vccd1 vccd1
+ _4679_/X sky130_fd_sc_hd__mux4_1
X_6418_ _6456_/B vssd1 vssd1 vccd1 vccd1 _6434_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_1_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6349_ _6461_/B _6461_/C _6341_/A _6461_/D _6355_/B vssd1 vssd1 vccd1 vccd1 _6397_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput104 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _6672_/A sky130_fd_sc_hd__buf_6
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8019_ _8486_/CLK _8019_/D vssd1 vssd1 vccd1 vccd1 _8019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7671__46 _7672__47/A vssd1 vssd1 vccd1 vccd1 _8515_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ _8488_/Q vssd1 vssd1 vccd1 vccd1 _3981_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5720_ _5720_/A vssd1 vssd1 vccd1 vccd1 _7924_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5651_ _7954_/Q _5650_/X _5653_/S vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5582_ _5582_/A vssd1 vssd1 vccd1 vccd1 _7989_/D sky130_fd_sc_hd__clkbuf_1
X_4602_ _4444_/X _8197_/Q _4602_/S vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__mux2_1
X_8370_ _8370_/CLK _8370_/D vssd1 vssd1 vccd1 vccd1 _8370_/Q sky130_fd_sc_hd__dfxtp_1
X_4533_ _4374_/X _8228_/Q _4541_/S vssd1 vssd1 vccd1 vccd1 _4534_/A sky130_fd_sc_hd__mux2_1
X_7321_ _7321_/A _7321_/B vssd1 vssd1 vccd1 vccd1 _8348_/D sky130_fd_sc_hd__nor2_1
XFILLER_117_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7252_ _8354_/Q vssd1 vssd1 vccd1 vccd1 _7252_/Y sky130_fd_sc_hd__inv_2
X_4464_ _4464_/A vssd1 vssd1 vccd1 vccd1 _8253_/D sky130_fd_sc_hd__clkbuf_1
X_6203_ _6200_/X _7815_/Q _6202_/X _6195_/X _7783_/Q vssd1 vssd1 vccd1 vccd1 _7783_/D
+ sky130_fd_sc_hd__o32a_1
X_7183_ _7432_/A vssd1 vssd1 vccd1 vccd1 _7183_/X sky130_fd_sc_hd__buf_1
XFILLER_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4395_ _4394_/X _8278_/Q _4398_/S vssd1 vssd1 vccd1 vccd1 _4396_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6134_ _7803_/Q _6122_/X _6126_/X _6133_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6134_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6065_ _7860_/Q input31/X _6072_/S vssd1 vssd1 vccd1 vccd1 _6065_/X sky130_fd_sc_hd__mux2_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5016_ _5031_/S vssd1 vssd1 vccd1 vccd1 _5025_/S sky130_fd_sc_hd__clkbuf_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5918_ _5918_/A vssd1 vssd1 vccd1 vccd1 _5918_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6776__362 _6777__363/A vssd1 vssd1 vccd1 vccd1 _8075_/CLK sky130_fd_sc_hd__inv_2
X_6898_ _8480_/Q _6900_/B vssd1 vssd1 vccd1 vccd1 _6899_/A sky130_fd_sc_hd__and2_1
X_5849_ _5611_/X _7775_/Q _5851_/S vssd1 vssd1 vccd1 vccd1 _5850_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3647_ _7439_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3647_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7519_ _7519_/A _7519_/B _7519_/C _6842_/B vssd1 vssd1 vccd1 vccd1 _7523_/A sky130_fd_sc_hd__or4b_1
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8499_ _8499_/CLK _8499_/D vssd1 vssd1 vccd1 vccd1 _8499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__3275_ clkbuf_0__3275_/X vssd1 vssd1 vccd1 vccd1 _6653__311/A sky130_fd_sc_hd__clkbuf_16
X_7169__89 _7169__89/A vssd1 vssd1 vccd1 vccd1 _8316_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4180_ _4180_/A vssd1 vssd1 vccd1 vccd1 _8393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7870_ _8537_/CLK _7870_/D vssd1 vssd1 vccd1 vccd1 _7870_/Q sky130_fd_sc_hd__dfxtp_1
X_6821_ _6849_/B _6830_/B _8467_/Q vssd1 vssd1 vccd1 vccd1 _7571_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3964_ _8457_/Q _3963_/X _3973_/S vssd1 vssd1 vccd1 vccd1 _3965_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5703_ _7931_/Q _5647_/X _5707_/S vssd1 vssd1 vccd1 vccd1 _5704_/A sky130_fd_sc_hd__mux2_1
X_3895_ _3895_/A vssd1 vssd1 vccd1 vccd1 _8518_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3464_ clkbuf_0__3464_/X vssd1 vssd1 vccd1 vccd1 _7122_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6683_ _6683_/A vssd1 vssd1 vccd1 vccd1 _8010_/D sky130_fd_sc_hd__clkbuf_1
X_5634_ _5634_/A vssd1 vssd1 vccd1 vccd1 _7961_/D sky130_fd_sc_hd__clkbuf_1
X_8422_ _8422_/CLK _8422_/D vssd1 vssd1 vccd1 vccd1 _8422_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3432_ _6962_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3432_/X sky130_fd_sc_hd__clkbuf_16
X_8353_ _8355_/CLK _8353_/D vssd1 vssd1 vccd1 vccd1 _8353_/Q sky130_fd_sc_hd__dfxtp_1
X_5565_ _5565_/A vssd1 vssd1 vccd1 vccd1 _7994_/D sky130_fd_sc_hd__clkbuf_1
X_7304_ _7301_/X _7302_/Y _7303_/Y _7302_/A _7286_/X vssd1 vssd1 vccd1 vccd1 _8343_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5496_ _8047_/Q _4295_/A _5498_/S vssd1 vssd1 vccd1 vccd1 _5497_/A sky130_fd_sc_hd__mux2_1
X_8284_ _8284_/CLK _8284_/D vssd1 vssd1 vccd1 vccd1 _8284_/Q sky130_fd_sc_hd__dfxtp_1
X_4516_ _4516_/A vssd1 vssd1 vccd1 vccd1 _8235_/D sky130_fd_sc_hd__clkbuf_1
X_4447_ _4490_/A _5464_/A vssd1 vssd1 vccd1 vccd1 _4463_/S sky130_fd_sc_hd__or2_2
X_7235_ _8543_/Q _7329_/A _7329_/B vssd1 vssd1 vccd1 vccd1 _7235_/X sky130_fd_sc_hd__and3_1
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4378_ _4378_/A vssd1 vssd1 vccd1 vccd1 _8284_/D sky130_fd_sc_hd__clkbuf_1
X_6117_ _6075_/A _6115_/X _6116_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6117_/X sky130_fd_sc_hd__o211a_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6048_ _6034_/X _6046_/X _6047_/X _6044_/X vssd1 vssd1 vccd1 vccd1 _6048_/X sky130_fd_sc_hd__o211a_1
XFILLER_27_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7999_ _8540_/CLK _7999_/D vssd1 vssd1 vccd1 vccd1 _7999_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6976__436 _6979__439/A vssd1 vssd1 vccd1 vccd1 _8160_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5350_ _5356_/A _5350_/B vssd1 vssd1 vccd1 vccd1 _5350_/Y sky130_fd_sc_hd__nand2_1
Xoutput205 _6067_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[6] sky130_fd_sc_hd__buf_2
X_5281_ _8380_/Q _8388_/Q _5281_/S vssd1 vssd1 vccd1 vccd1 _5281_/X sky130_fd_sc_hd__mux2_2
X_4301_ _4301_/A _4301_/B _4256_/C vssd1 vssd1 vccd1 vccd1 _4356_/B sky130_fd_sc_hd__or3b_1
X_4232_ _4232_/A vssd1 vssd1 vccd1 vccd1 _8373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7296__112 _7297__113/A vssd1 vssd1 vccd1 vccd1 _8341_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4163_ _8108_/Q vssd1 vssd1 vccd1 vccd1 _4163_/X sky130_fd_sc_hd__buf_2
X_4094_ _4035_/X _8411_/Q _4094_/S vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7922_ _7922_/CLK _7922_/D vssd1 vssd1 vccd1 vccd1 _7922_/Q sky130_fd_sc_hd__dfxtp_1
X_7853_ _7853_/CLK _7853_/D vssd1 vssd1 vccd1 vccd1 _7853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4996_ _5823_/A _5555_/A vssd1 vssd1 vccd1 vccd1 _5012_/S sky130_fd_sc_hd__nor2_2
X_7784_ _8543_/CLK _7784_/D vssd1 vssd1 vccd1 vccd1 _7784_/Q sky130_fd_sc_hd__dfxtp_1
X_6804_ _6804_/A _6830_/A _6824_/B vssd1 vssd1 vccd1 vccd1 _6816_/B sky130_fd_sc_hd__nand3_2
X_3947_ _3947_/A vssd1 vssd1 vccd1 vccd1 _8499_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3447_ clkbuf_0__3447_/X vssd1 vssd1 vccd1 vccd1 _7038__484/A sky130_fd_sc_hd__clkbuf_4
X_6666_ _5930_/A _8003_/Q _6670_/S vssd1 vssd1 vccd1 vccd1 _6667_/A sky130_fd_sc_hd__mux2_1
X_3878_ _6355_/A _6337_/A vssd1 vssd1 vccd1 vccd1 _6398_/A sky130_fd_sc_hd__or2_2
X_5617_ _5617_/A vssd1 vssd1 vccd1 vccd1 _7976_/D sky130_fd_sc_hd__clkbuf_1
X_8405_ _8405_/CLK _8405_/D vssd1 vssd1 vccd1 vccd1 _8405_/Q sky130_fd_sc_hd__dfxtp_1
X_8336_ _8336_/CLK _8336_/D vssd1 vssd1 vccd1 vccd1 _8336_/Q sky130_fd_sc_hd__dfxtp_1
X_5548_ _5379_/X _8024_/Q _5552_/S vssd1 vssd1 vccd1 vccd1 _5549_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_opt_3_0_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8267_ _8267_/CLK _8267_/D vssd1 vssd1 vccd1 vccd1 _8267_/Q sky130_fd_sc_hd__dfxtp_1
X_5479_ _5479_/A vssd1 vssd1 vccd1 vccd1 _8055_/D sky130_fd_sc_hd__clkbuf_1
X_7218_ _8353_/Q _7232_/B _7232_/C _7218_/D vssd1 vssd1 vccd1 vccd1 _7220_/A sky130_fd_sc_hd__nand4_2
XFILLER_59_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8198_ _8198_/CLK _8198_/D vssd1 vssd1 vccd1 vccd1 _8198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4850_ _7912_/Q _8084_/Q _4880_/S vssd1 vssd1 vccd1 vccd1 _4850_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4781_ _4781_/A vssd1 vssd1 vccd1 vccd1 _4781_/X sky130_fd_sc_hd__clkbuf_2
X_6520_ _6388_/X _6517_/Y _6522_/B vssd1 vssd1 vccd1 vccd1 _7899_/D sky130_fd_sc_hd__o21a_1
XFILLER_119_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6451_ _7871_/Q _6442_/X _6437_/X _6450_/X _6435_/X vssd1 vssd1 vccd1 vccd1 _7871_/D
+ sky130_fd_sc_hd__a221o_1
X_5402_ _5375_/X _8093_/Q _5402_/S vssd1 vssd1 vccd1 vccd1 _5403_/A sky130_fd_sc_hd__mux2_1
X_6382_ _6382_/A vssd1 vssd1 vccd1 vccd1 _6410_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5333_ _5343_/B _5787_/B _5332_/X _5262_/X vssd1 vssd1 vccd1 vccd1 _8123_/D sky130_fd_sc_hd__o211a_1
X_8121_ _8121_/CLK _8121_/D vssd1 vssd1 vccd1 vccd1 _8121_/Q sky130_fd_sc_hd__dfxtp_1
X_8052_ _8052_/CLK _8052_/D vssd1 vssd1 vccd1 vccd1 _8052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5264_ _5264_/A vssd1 vssd1 vccd1 vccd1 _5356_/B sky130_fd_sc_hd__clkbuf_2
X_4215_ _8379_/Q _4196_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__mux2_1
X_5195_ _8454_/Q _8192_/Q _5315_/S vssd1 vssd1 vccd1 vccd1 _5195_/X sky130_fd_sc_hd__mux2_1
X_4146_ _5751_/A vssd1 vssd1 vccd1 vccd1 _5641_/A sky130_fd_sc_hd__buf_4
X_6547__241 _6549__243/A vssd1 vssd1 vccd1 vccd1 _7919_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7415__136 _7416__137/A vssd1 vssd1 vccd1 vccd1 _8393_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4301_/B _5334_/B _4256_/A vssd1 vssd1 vccd1 vccd1 _4199_/B sky130_fd_sc_hd__nand3b_4
X_7905_ _7905_/CLK _7905_/D vssd1 vssd1 vccd1 vccd1 _7905_/Q sky130_fd_sc_hd__dfxtp_1
X_7836_ _7836_/CLK _7836_/D vssd1 vssd1 vccd1 vccd1 _7836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7767_ _7767_/CLK _7767_/D vssd1 vssd1 vccd1 vccd1 _7767_/Q sky130_fd_sc_hd__dfxtp_1
X_4979_ _4994_/S vssd1 vssd1 vccd1 vccd1 _4988_/S sky130_fd_sc_hd__buf_2
X_6718_ _6718_/A vssd1 vssd1 vccd1 vccd1 _6718_/X sky130_fd_sc_hd__buf_1
X_7698_ _7742_/B _7742_/C _7698_/C _7698_/D vssd1 vssd1 vccd1 vccd1 _7747_/B sky130_fd_sc_hd__nor4_4
XFILLER_105_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8319_ _8319_/CLK _8319_/D vssd1 vssd1 vccd1 vccd1 _8319_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3646_ clkbuf_0__3646_/X vssd1 vssd1 vccd1 vccd1 _7438__155/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4000_ _3908_/X _8444_/Q _4002_/S vssd1 vssd1 vccd1 vccd1 _4001_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5951_ _5951_/A vssd1 vssd1 vccd1 vccd1 _5951_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4902_ _8229_/Q _4775_/X _4781_/A _8213_/Q _4733_/A vssd1 vssd1 vccd1 vccd1 _4902_/X
+ sky130_fd_sc_hd__o221a_1
X_6323__221 _6325__223/A vssd1 vssd1 vccd1 vccd1 _7851_/CLK sky130_fd_sc_hd__inv_2
X_5882_ _5898_/A vssd1 vssd1 vccd1 vccd1 _6021_/A sky130_fd_sc_hd__inv_6
X_4833_ _7928_/Q _4658_/B _4784_/X vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7621_ _8483_/Q _7614_/X vssd1 vssd1 vccd1 vccd1 _7621_/X sky130_fd_sc_hd__or2b_1
XFILLER_33_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7552_ _7552_/A vssd1 vssd1 vccd1 vccd1 _7552_/X sky130_fd_sc_hd__clkbuf_2
X_4764_ _5399_/A _4764_/B vssd1 vssd1 vccd1 vccd1 _4764_/X sky130_fd_sc_hd__or2_1
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6770__357 _6772__359/A vssd1 vssd1 vccd1 vccd1 _8070_/CLK sky130_fd_sc_hd__inv_2
X_6503_ _8008_/Q _7893_/Q _6509_/S vssd1 vssd1 vccd1 vccd1 _6504_/A sky130_fd_sc_hd__mux2_1
X_4695_ _4654_/X _4693_/X _4694_/X vssd1 vssd1 vccd1 vccd1 _4695_/X sky130_fd_sc_hd__a21o_1
X_6434_ _7528_/A _6434_/B _6444_/C vssd1 vssd1 vccd1 vccd1 _6434_/X sky130_fd_sc_hd__and3_1
X_6365_ _6362_/A _7967_/Q _6382_/A _6364_/X vssd1 vssd1 vccd1 vccd1 _6365_/X sky130_fd_sc_hd__a31o_1
X_6176__184 _6177__185/A vssd1 vssd1 vccd1 vccd1 _7771_/CLK sky130_fd_sc_hd__inv_2
X_5316_ _5196_/X _8073_/Q _7838_/Q _5198_/X _5092_/A vssd1 vssd1 vccd1 vccd1 _5316_/X
+ sky130_fd_sc_hd__o221a_1
X_8104_ _8104_/CLK _8104_/D vssd1 vssd1 vccd1 vccd1 _8104_/Q sky130_fd_sc_hd__dfxtp_1
X_8035_ _8035_/CLK _8035_/D vssd1 vssd1 vccd1 vccd1 _8035_/Q sky130_fd_sc_hd__dfxtp_1
X_5247_ _5306_/A _5245_/X _5246_/X vssd1 vssd1 vccd1 vccd1 _5247_/X sky130_fd_sc_hd__o21a_1
X_5178_ _8116_/Q vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0__3431_ clkbuf_0__3431_/X vssd1 vssd1 vccd1 vccd1 _7089_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4129_ _8175_/Q _8170_/Q vssd1 vssd1 vccd1 vccd1 _4622_/A sky130_fd_sc_hd__xor2_1
XFILLER_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7819_ _8355_/CLK _7819_/D vssd1 vssd1 vccd1 vccd1 _7819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6730__330 _6730__330/A vssd1 vssd1 vccd1 vccd1 _8040_/CLK sky130_fd_sc_hd__inv_2
X_4480_ _4480_/A vssd1 vssd1 vccd1 vccd1 _8248_/D sky130_fd_sc_hd__clkbuf_1
X_6150_ _7809_/Q _6138_/X _6139_/X _6149_/X _6063_/A vssd1 vssd1 vccd1 vccd1 _6150_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5096_/X _5099_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _5101_/X sky130_fd_sc_hd__mux2_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _7789_/Q _6086_/B vssd1 vssd1 vccd1 vccd1 _6081_/X sky130_fd_sc_hd__or2_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5032_ _5032_/A vssd1 vssd1 vccd1 vccd1 _8135_/D sky130_fd_sc_hd__clkbuf_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8520_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5934_ _5956_/A vssd1 vssd1 vccd1 vccd1 _5943_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5865_ _4154_/X _7768_/Q _5869_/S vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__mux2_1
X_4816_ _4805_/A _7905_/Q _4806_/A _8138_/Q _4663_/A vssd1 vssd1 vccd1 vccd1 _4816_/X
+ sky130_fd_sc_hd__o221a_1
X_7604_ _6865_/B _7602_/Y _7603_/X _7568_/A vssd1 vssd1 vccd1 vccd1 _8477_/D sky130_fd_sc_hd__a211oi_1
X_5796_ _5796_/A vssd1 vssd1 vccd1 vccd1 _7842_/D sky130_fd_sc_hd__clkbuf_1
X_4747_ _8217_/Q _8201_/Q _8163_/Q _8233_/Q _4655_/X _4656_/X vssd1 vssd1 vccd1 vccd1
+ _4747_/X sky130_fd_sc_hd__mux4_1
X_7535_ _7524_/X _7535_/B _7535_/C _7535_/D vssd1 vssd1 vccd1 vccd1 _7535_/X sky130_fd_sc_hd__and4b_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4678_ _7770_/Q _7778_/Q _7853_/Q _7957_/Q _4666_/X _4667_/X vssd1 vssd1 vccd1 vccd1
+ _4678_/X sky130_fd_sc_hd__mux4_2
XFILLER_110_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6417_ _6417_/A vssd1 vssd1 vccd1 vccd1 _6456_/B sky130_fd_sc_hd__buf_2
X_6348_ _7742_/C _6348_/B _6348_/C _6348_/D vssd1 vssd1 vccd1 vccd1 _6355_/B sky130_fd_sc_hd__or4_1
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput105 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _6690_/A sky130_fd_sc_hd__buf_6
X_6279_ _8362_/Q _8363_/Q _8364_/Q _8365_/Q _8359_/Q _8360_/Q vssd1 vssd1 vccd1 vccd1
+ _6280_/B sky130_fd_sc_hd__mux4_1
XFILLER_102_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8018_ _8486_/CLK _8018_/D vssd1 vssd1 vccd1 vccd1 _8018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7290__107 _7290__107/A vssd1 vssd1 vccd1 vccd1 _8336_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3980_ _3980_/A vssd1 vssd1 vccd1 vccd1 _8452_/D sky130_fd_sc_hd__clkbuf_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5650_ _8110_/Q vssd1 vssd1 vccd1 vccd1 _5650_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4601_ _4601_/A vssd1 vssd1 vccd1 vccd1 _8198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5581_ _7989_/Q _5578_/X _5591_/S vssd1 vssd1 vccd1 vccd1 _5582_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4532_ _4547_/S vssd1 vssd1 vccd1 vccd1 _4541_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7320_ _7227_/A _7318_/X _7310_/X _7319_/Y vssd1 vssd1 vccd1 vccd1 _7321_/B sky130_fd_sc_hd__o2bb2a_1
X_4463_ _4397_/X _8253_/Q _4463_/S vssd1 vssd1 vccd1 vccd1 _4464_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7251_ _7251_/A _7251_/B _7251_/C _7251_/D vssd1 vssd1 vccd1 vccd1 _7263_/C sky130_fd_sc_hd__and4_1
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6202_ _6202_/A vssd1 vssd1 vccd1 vccd1 _6202_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4394_ _8489_/Q vssd1 vssd1 vccd1 vccd1 _4394_/X sky130_fd_sc_hd__clkbuf_2
X_6133_ _6133_/A _6140_/B vssd1 vssd1 vccd1 vccd1 _6133_/X sky130_fd_sc_hd__and2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6064_ _6056_/X _6061_/X _6062_/X _6063_/X vssd1 vssd1 vccd1 vccd1 _6064_/X sky130_fd_sc_hd__o211a_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7023__472 _7023__472/A vssd1 vssd1 vccd1 vccd1 _8199_/CLK sky130_fd_sc_hd__inv_2
X_5015_ _5859_/A _5751_/B vssd1 vssd1 vccd1 vccd1 _5031_/S sky130_fd_sc_hd__or2_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5917_ _7646_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__or2_1
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5848_ _5848_/A vssd1 vssd1 vccd1 vccd1 _7776_/D sky130_fd_sc_hd__clkbuf_1
X_6930__404 _6930__404/A vssd1 vssd1 vccd1 vccd1 _8126_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3646_ _7433_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3646_/X sky130_fd_sc_hd__clkbuf_16
X_5779_ _5566_/X _7849_/Q _5779_/S vssd1 vssd1 vccd1 vccd1 _5780_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7518_ _8548_/Q _7518_/B _7556_/B vssd1 vssd1 vccd1 vccd1 _7519_/C sky130_fd_sc_hd__and3b_1
X_8498_ _8498_/CLK _8498_/D vssd1 vssd1 vccd1 vccd1 _8498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3259_ clkbuf_0__3259_/X vssd1 vssd1 vccd1 vccd1 _6625__290/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6820_ _8467_/Q _6849_/B _6830_/B vssd1 vssd1 vccd1 vccd1 _7571_/A sky130_fd_sc_hd__nand3_2
X_6541__236 _6544__239/A vssd1 vssd1 vccd1 vccd1 _7914_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3963_ _8494_/Q vssd1 vssd1 vccd1 vccd1 _3963_/X sky130_fd_sc_hd__buf_4
X_5702_ _5702_/A vssd1 vssd1 vccd1 vccd1 _7932_/D sky130_fd_sc_hd__clkbuf_1
X_3894_ _3893_/X _8518_/Q _3903_/S vssd1 vssd1 vccd1 vccd1 _3895_/A sky130_fd_sc_hd__mux2_1
X_6682_ _5946_/A _8010_/Q _6682_/S vssd1 vssd1 vccd1 vccd1 _6683_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_5633_ _5566_/X _7961_/Q _5633_/S vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__mux2_1
X_8421_ _8421_/CLK _8421_/D vssd1 vssd1 vccd1 vccd1 _8421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5564_ _5399_/X _7994_/Q _5567_/S vssd1 vssd1 vccd1 vccd1 _5565_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3431_ _6961_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3431_/X sky130_fd_sc_hd__clkbuf_16
X_8352_ _8355_/CLK _8352_/D vssd1 vssd1 vccd1 vccd1 _8352_/Q sky130_fd_sc_hd__dfxtp_1
X_7303_ _7303_/A _7303_/B vssd1 vssd1 vccd1 vccd1 _7303_/Y sky130_fd_sc_hd__nor2_1
X_4515_ _8235_/Q _4471_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5495_ _5495_/A vssd1 vssd1 vccd1 vccd1 _8048_/D sky130_fd_sc_hd__clkbuf_1
X_8585__232 vssd1 vssd1 vccd1 vccd1 _8585__232/HI manufacturerID[4] sky130_fd_sc_hd__conb_1
X_8283_ _8283_/CLK _8283_/D vssd1 vssd1 vccd1 vccd1 _8283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4446_ _4446_/A vssd1 vssd1 vccd1 vccd1 _8261_/D sky130_fd_sc_hd__clkbuf_1
X_7234_ _7329_/A _7329_/B _8543_/Q vssd1 vssd1 vccd1 vccd1 _7234_/Y sky130_fd_sc_hd__a21oi_1
X_7165_ _7165_/A vssd1 vssd1 vccd1 vccd1 _7165_/X sky130_fd_sc_hd__buf_1
X_4377_ _4374_/X _8284_/Q _4389_/S vssd1 vssd1 vccd1 vccd1 _4378_/A sky130_fd_sc_hd__mux2_1
X_6116_ _7798_/Q _6122_/A vssd1 vssd1 vccd1 vccd1 _6116_/X sky130_fd_sc_hd__or2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7096_ _7108_/A vssd1 vssd1 vccd1 vccd1 _7096_/X sky130_fd_sc_hd__buf_1
XFILLER_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6047_ _7780_/Q _7633_/A vssd1 vssd1 vccd1 vccd1 _6047_/X sky130_fd_sc_hd__or2_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7998_ _8540_/CLK _7998_/D vssd1 vssd1 vccd1 vccd1 _7998_/Q sky130_fd_sc_hd__dfxtp_1
X_6949_ _6955_/A vssd1 vssd1 vccd1 vccd1 _6949_/X sky130_fd_sc_hd__buf_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7174__93 _7176__95/A vssd1 vssd1 vccd1 vccd1 _8320_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8569__216 vssd1 vssd1 vccd1 vccd1 _8569__216/HI core0Index[3] sky130_fd_sc_hd__conb_1
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput206 _6071_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_114_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5280_ _5206_/A _5268_/Y _5272_/Y _5279_/X vssd1 vssd1 vccd1 vccd1 _5295_/A sky130_fd_sc_hd__a31o_1
X_4300_ _4300_/A vssd1 vssd1 vccd1 vccd1 _8317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4231_ _8373_/Q _4163_/X _4235_/S vssd1 vssd1 vccd1 vccd1 _4232_/A sky130_fd_sc_hd__mux2_1
X_4162_ _4162_/A vssd1 vssd1 vccd1 vccd1 _8398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6170__179 _6170__179/A vssd1 vssd1 vccd1 vccd1 _7766_/CLK sky130_fd_sc_hd__inv_2
X_4093_ _4093_/A vssd1 vssd1 vccd1 vccd1 _8412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7921_ _7921_/CLK _7921_/D vssd1 vssd1 vccd1 vccd1 _7921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7852_ _7852_/CLK _7852_/D vssd1 vssd1 vccd1 vccd1 _7852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4995_ _4995_/A vssd1 vssd1 vccd1 vccd1 _8151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6803_ _8539_/Q _7528_/B vssd1 vssd1 vccd1 vccd1 _6808_/C sky130_fd_sc_hd__xor2_1
X_7783_ _8543_/CLK _7783_/D vssd1 vssd1 vccd1 vccd1 _7783_/Q sky130_fd_sc_hd__dfxtp_1
X_3946_ _3902_/X _8499_/Q _3946_/S vssd1 vssd1 vccd1 vccd1 _3947_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3446_ clkbuf_0__3446_/X vssd1 vssd1 vccd1 vccd1 _7033__480/A sky130_fd_sc_hd__clkbuf_4
X_8404_ _8404_/CLK _8404_/D vssd1 vssd1 vccd1 vccd1 _8404_/Q sky130_fd_sc_hd__dfxtp_1
X_6665_ _6665_/A vssd1 vssd1 vccd1 vccd1 _8002_/D sky130_fd_sc_hd__clkbuf_1
X_3877_ _7879_/Q _7880_/Q _6345_/B vssd1 vssd1 vccd1 vccd1 _6337_/A sky130_fd_sc_hd__or3_1
X_6596_ _6632_/A vssd1 vssd1 vccd1 vccd1 _6596_/X sky130_fd_sc_hd__buf_1
X_5616_ _5569_/X _7976_/Q _5620_/S vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8335_ _8335_/CLK _8335_/D vssd1 vssd1 vccd1 vccd1 _8335_/Q sky130_fd_sc_hd__dfxtp_1
X_5547_ _5547_/A vssd1 vssd1 vccd1 vccd1 _8025_/D sky130_fd_sc_hd__clkbuf_1
X_8266_ _8266_/CLK _8266_/D vssd1 vssd1 vccd1 vccd1 _8266_/Q sky130_fd_sc_hd__dfxtp_1
X_5478_ _3978_/X _8055_/Q _5480_/S vssd1 vssd1 vccd1 vccd1 _5479_/A sky130_fd_sc_hd__mux2_1
X_4429_ _4428_/X _8266_/Q _4436_/S vssd1 vssd1 vccd1 vccd1 _4430_/A sky130_fd_sc_hd__mux2_1
X_7217_ _8352_/Q _8351_/Q vssd1 vssd1 vccd1 vccd1 _7218_/D sky130_fd_sc_hd__and2_1
X_8197_ _8197_/CLK _8197_/D vssd1 vssd1 vccd1 vccd1 _8197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7036__482 _7039__485/A vssd1 vssd1 vccd1 vccd1 _8209_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3027_ clkbuf_0__3027_/X vssd1 vssd1 vccd1 vccd1 _6290__195/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7147__71 _7149__73/A vssd1 vssd1 vccd1 vccd1 _8298_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6982__441 _6983__442/A vssd1 vssd1 vccd1 vccd1 _8165_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7078__516 _7079__517/A vssd1 vssd1 vccd1 vccd1 _8243_/CLK sky130_fd_sc_hd__inv_2
X_7004__459 _7005__460/A vssd1 vssd1 vccd1 vccd1 _8184_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4780_ _4797_/A vssd1 vssd1 vccd1 vccd1 _4781_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6450_ _7008_/A _6452_/B _6454_/C vssd1 vssd1 vccd1 vccd1 _6450_/X sky130_fd_sc_hd__and3_1
X_6381_ _7857_/Q _6328_/X _6380_/X vssd1 vssd1 vccd1 vccd1 _7857_/D sky130_fd_sc_hd__a21o_1
X_5401_ _5401_/A vssd1 vssd1 vccd1 vccd1 _8094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5332_ _5334_/A _5334_/B _5334_/C _4256_/A vssd1 vssd1 vccd1 vccd1 _5332_/X sky130_fd_sc_hd__a31o_1
X_8120_ _8120_/CLK _8120_/D vssd1 vssd1 vccd1 vccd1 _8120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8051_ _8051_/CLK _8051_/D vssd1 vssd1 vccd1 vccd1 _8051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5263_ _3905_/X _5038_/A _5261_/X _5262_/X vssd1 vssd1 vccd1 vccd1 _8127_/D sky130_fd_sc_hd__o211a_1
X_5194_ _5321_/S vssd1 vssd1 vccd1 vccd1 _5315_/S sky130_fd_sc_hd__clkbuf_4
X_4214_ _4214_/A vssd1 vssd1 vccd1 vccd1 _8380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4145_ _4217_/A _4944_/A _4931_/B vssd1 vssd1 vccd1 vccd1 _5751_/A sky130_fd_sc_hd__or3_4
XFILLER_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4076_ _4076_/A vssd1 vssd1 vccd1 vccd1 _5334_/B sky130_fd_sc_hd__clkbuf_2
X_7904_ _7904_/CLK _7904_/D vssd1 vssd1 vccd1 vccd1 _7904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7835_ _7835_/CLK _7835_/D vssd1 vssd1 vccd1 vccd1 _7835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7766_ _7766_/CLK _7766_/D vssd1 vssd1 vccd1 vccd1 _7766_/Q sky130_fd_sc_hd__dfxtp_1
X_4978_ _5641_/A _5733_/B vssd1 vssd1 vccd1 vccd1 _4994_/S sky130_fd_sc_hd__nor2_2
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3929_ _3905_/X _8506_/Q _3933_/S vssd1 vssd1 vccd1 vccd1 _3930_/A sky130_fd_sc_hd__mux2_1
X_7697_ _7878_/Q _6348_/C _6352_/A vssd1 vssd1 vccd1 vccd1 _7698_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_1_1_0__3429_ clkbuf_0__3429_/X vssd1 vssd1 vccd1 vccd1 _6954__420/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8318_ _8318_/CLK _8318_/D vssd1 vssd1 vccd1 vccd1 _8318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8249_ _8249_/CLK _8249_/D vssd1 vssd1 vccd1 vccd1 _8249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3259_ _6602_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3259_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3645_ clkbuf_0__3645_/X vssd1 vssd1 vccd1 vccd1 _7457_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _5950_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _5951_/A sky130_fd_sc_hd__or2_4
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4901_ _8159_/Q _8197_/Q _4901_/S vssd1 vssd1 vccd1 vccd1 _4901_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5881_ _5881_/A _6161_/C vssd1 vssd1 vccd1 vccd1 _5898_/A sky130_fd_sc_hd__or2_2
X_7620_ _8483_/Q _7613_/X _7619_/X _7552_/X vssd1 vssd1 vccd1 vccd1 _8482_/D sky130_fd_sc_hd__o211a_1
X_4832_ _8247_/Q _4781_/X _4755_/A _4831_/X vssd1 vssd1 vccd1 vccd1 _4832_/X sky130_fd_sc_hd__o211a_1
XFILLER_119_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7551_ _7547_/X _7551_/B vssd1 vssd1 vccd1 vccd1 _7551_/X sky130_fd_sc_hd__and2b_1
X_4763_ _4713_/X _8183_/Q _4947_/A _4762_/X vssd1 vssd1 vccd1 vccd1 _4763_/X sky130_fd_sc_hd__a22o_1
X_7482_ _7482_/A vssd1 vssd1 vccd1 vccd1 _7482_/X sky130_fd_sc_hd__buf_1
X_4694_ _4694_/A vssd1 vssd1 vccd1 vccd1 _4694_/X sky130_fd_sc_hd__buf_2
X_6502_ _6502_/A vssd1 vssd1 vccd1 vccd1 _7892_/D sky130_fd_sc_hd__clkbuf_1
X_6989__447 _6989__447/A vssd1 vssd1 vccd1 vccd1 _8172_/CLK sky130_fd_sc_hd__inv_2
X_6433_ _8538_/Q vssd1 vssd1 vccd1 vccd1 _7528_/A sky130_fd_sc_hd__buf_2
X_7472__7 _7472__7/A vssd1 vssd1 vccd1 vccd1 _8439_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7421__141 _7422__142/A vssd1 vssd1 vccd1 vccd1 _8398_/CLK sky130_fd_sc_hd__inv_2
X_6364_ _6395_/A vssd1 vssd1 vccd1 vccd1 _6364_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5315_ _8325_/Q _8046_/Q _5315_/S vssd1 vssd1 vccd1 vccd1 _5315_/X sky130_fd_sc_hd__mux2_1
X_8103_ _8103_/CLK _8103_/D vssd1 vssd1 vccd1 vccd1 _8103_/Q sky130_fd_sc_hd__dfxtp_1
X_7141__66 _7145__70/A vssd1 vssd1 vccd1 vccd1 _8293_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5246_ _5196_/X _8075_/Q _7840_/Q _5207_/A _5092_/A vssd1 vssd1 vccd1 vccd1 _5246_/X
+ sky130_fd_sc_hd__o221a_1
X_8034_ _8034_/CLK _8034_/D vssd1 vssd1 vccd1 vccd1 _8034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3430_ clkbuf_0__3430_/X vssd1 vssd1 vccd1 vccd1 _6957__422/A sky130_fd_sc_hd__clkbuf_4
X_5177_ _5177_/A vssd1 vssd1 vccd1 vccd1 _5350_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4128_ _8174_/Q vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__inv_2
X_4059_ _4074_/S vssd1 vssd1 vccd1 vccd1 _4068_/S sky130_fd_sc_hd__buf_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7818_ _8543_/CLK _7818_/D vssd1 vssd1 vccd1 vccd1 _7818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7749_ _8545_/Q _7747_/Y _7748_/X vssd1 vssd1 vccd1 vccd1 _8545_/D sky130_fd_sc_hd__a21o_1
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6643__303 _6643__303/A vssd1 vssd1 vccd1 vccd1 _7989_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5100_ _5100_/A vssd1 vssd1 vccd1 vccd1 _5101_/S sky130_fd_sc_hd__buf_2
X_6080_ _7864_/Q input4/X _6092_/S vssd1 vssd1 vccd1 vccd1 _6080_/X sky130_fd_sc_hd__mux2_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _4444_/X _8135_/Q _5031_/S vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__mux2_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6995__451 _6998__454/A vssd1 vssd1 vccd1 vccd1 _8176_/CLK sky130_fd_sc_hd__inv_2
X_5933_ _5933_/A vssd1 vssd1 vccd1 vccd1 _5933_/X sky130_fd_sc_hd__clkbuf_1
X_5864_ _5864_/A vssd1 vssd1 vccd1 vccd1 _7769_/D sky130_fd_sc_hd__clkbuf_1
X_7189__105 _7189__105/A vssd1 vssd1 vccd1 vccd1 _8332_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4815_ _7921_/Q _8025_/Q _4883_/S vssd1 vssd1 vccd1 vccd1 _4815_/X sky130_fd_sc_hd__mux2_1
X_7603_ _8477_/Q _7505_/A _7614_/A _6867_/C _7597_/X vssd1 vssd1 vccd1 vccd1 _7603_/X
+ sky130_fd_sc_hd__o221a_1
X_5795_ _7842_/Q _4286_/A _5797_/S vssd1 vssd1 vccd1 vccd1 _5796_/A sky130_fd_sc_hd__mux2_1
X_7534_ _6440_/A _6793_/B _7531_/Y _7532_/X _7533_/Y vssd1 vssd1 vccd1 vccd1 _7535_/D
+ sky130_fd_sc_hd__o221a_1
X_4746_ _8375_/Q _8265_/Q _7978_/Q _8399_/Q _4646_/X _4716_/X vssd1 vssd1 vccd1 vccd1
+ _4746_/X sky130_fd_sc_hd__mux4_2
X_4677_ _4675_/X _4676_/X _4677_/S vssd1 vssd1 vccd1 vccd1 _4677_/X sky130_fd_sc_hd__mux2_1
X_6416_ _8542_/Q vssd1 vssd1 vccd1 vccd1 _7514_/A sky130_fd_sc_hd__clkbuf_4
X_6347_ _7878_/Q _6521_/B vssd1 vssd1 vccd1 vccd1 _6348_/D sky130_fd_sc_hd__nand2_1
XFILLER_115_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6631__295 _6631__295/A vssd1 vssd1 vccd1 vccd1 _7981_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput106 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _6465_/A sky130_fd_sc_hd__buf_6
X_6278_ _8366_/Q _8367_/Q _8368_/Q _8369_/Q _7356_/B _8360_/Q vssd1 vssd1 vccd1 vccd1
+ _6278_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5229_ _5264_/A _5226_/X _5228_/X vssd1 vssd1 vccd1 vccd1 _5235_/B sky130_fd_sc_hd__o21a_1
XFILLER_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8017_ _8486_/CLK _8017_/D vssd1 vssd1 vccd1 vccd1 _8017_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3027_ _6184_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3027_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7428__147 _7429__148/A vssd1 vssd1 vccd1 vccd1 _8404_/CLK sky130_fd_sc_hd__inv_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7656__34 _7656__34/A vssd1 vssd1 vccd1 vccd1 _8503_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4600_ _4441_/X _8198_/Q _4602_/S vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__mux2_1
X_5580_ _5600_/S vssd1 vssd1 vccd1 vccd1 _5591_/S sky130_fd_sc_hd__buf_2
XFILLER_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4531_ _4531_/A _4604_/A vssd1 vssd1 vccd1 vccd1 _4547_/S sky130_fd_sc_hd__or2_2
XFILLER_7_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4462_ _4462_/A vssd1 vssd1 vccd1 vccd1 _8254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7250_ _7234_/Y _7235_/X _7281_/C _7280_/C _7281_/D vssd1 vssd1 vccd1 vccd1 _7251_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_116_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6201_ _6200_/X _7814_/Q _6191_/X _6195_/X _7782_/Q vssd1 vssd1 vccd1 vccd1 _7782_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4393_ _4393_/A vssd1 vssd1 vccd1 vccd1 _8279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6132_ _7802_/Q _6122_/X _6126_/X _6131_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6132_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6063_ _6063_/A vssd1 vssd1 vccd1 vccd1 _6063_/X sky130_fd_sc_hd__clkbuf_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5014_ _5014_/A _5014_/B _5014_/C vssd1 vssd1 vccd1 vccd1 _5751_/B sky130_fd_sc_hd__nand3_4
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5916_ _5916_/A vssd1 vssd1 vccd1 vccd1 _5916_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6896_ _6919_/A vssd1 vssd1 vccd1 vccd1 _6896_/X sky130_fd_sc_hd__buf_1
X_5847_ _5608_/X _7776_/Q _5851_/S vssd1 vssd1 vccd1 vccd1 _5848_/A sky130_fd_sc_hd__mux2_1
X_5778_ _5778_/A vssd1 vssd1 vccd1 vccd1 _7850_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3645_ _7432_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3645_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4729_ _4880_/S vssd1 vssd1 vccd1 vccd1 _4729_/X sky130_fd_sc_hd__buf_4
X_8497_ _8497_/CLK _8497_/D vssd1 vssd1 vccd1 vccd1 _8497_/Q sky130_fd_sc_hd__dfxtp_1
X_7517_ _7556_/A _7556_/B _7754_/A vssd1 vssd1 vccd1 vccd1 _7519_/B sky130_fd_sc_hd__a21boi_1
X_7030__477 _7030__477/A vssd1 vssd1 vccd1 vccd1 _8204_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7379_ _8367_/Q _7383_/B vssd1 vssd1 vccd1 vccd1 _7379_/X sky130_fd_sc_hd__or2_1
XFILLER_115_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7434__151 _7436__153/A vssd1 vssd1 vccd1 vccd1 _8408_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__3411_ clkbuf_0__3411_/X vssd1 vssd1 vccd1 vccd1 _6897__391/A sky130_fd_sc_hd__clkbuf_16
XFILLER_17_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3258_ clkbuf_0__3258_/X vssd1 vssd1 vccd1 vccd1 _6600__284/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5701_ _7932_/Q _5583_/X _5707_/S vssd1 vssd1 vccd1 vccd1 _5702_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3962_ _3962_/A vssd1 vssd1 vccd1 vccd1 _8458_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3462_ clkbuf_0__3462_/X vssd1 vssd1 vccd1 vccd1 _7119__550/A sky130_fd_sc_hd__clkbuf_4
X_3893_ _8494_/Q vssd1 vssd1 vccd1 vccd1 _3893_/X sky130_fd_sc_hd__buf_4
X_6681_ _6681_/A vssd1 vssd1 vccd1 vccd1 _8009_/D sky130_fd_sc_hd__clkbuf_1
X_5632_ _5632_/A vssd1 vssd1 vccd1 vccd1 _7962_/D sky130_fd_sc_hd__clkbuf_1
X_8420_ _8420_/CLK _8420_/D vssd1 vssd1 vccd1 vccd1 _8420_/Q sky130_fd_sc_hd__dfxtp_1
X_5563_ _5563_/A vssd1 vssd1 vccd1 vccd1 _7995_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3430_ _6955_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3430_/X sky130_fd_sc_hd__clkbuf_16
X_8351_ _8358_/CLK _8351_/D vssd1 vssd1 vccd1 vccd1 _8351_/Q sky130_fd_sc_hd__dfxtp_1
X_4514_ _4514_/A vssd1 vssd1 vccd1 vccd1 _8236_/D sky130_fd_sc_hd__clkbuf_1
X_7302_ _7302_/A _7308_/A vssd1 vssd1 vccd1 vccd1 _7302_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5494_ _8048_/Q _4292_/A _5498_/S vssd1 vssd1 vccd1 vccd1 _5495_/A sky130_fd_sc_hd__mux2_1
X_8282_ _8282_/CLK _8282_/D vssd1 vssd1 vccd1 vccd1 _8282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4445_ _4444_/X _8261_/Q _4445_/S vssd1 vssd1 vccd1 vccd1 _4446_/A sky130_fd_sc_hd__mux2_1
X_7233_ _7236_/B _7232_/C _8351_/Q vssd1 vssd1 vccd1 vccd1 _7329_/B sky130_fd_sc_hd__a21o_1
X_4376_ _4398_/S vssd1 vssd1 vccd1 vccd1 _4389_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _7873_/Q input13/X _6153_/B vssd1 vssd1 vccd1 vccd1 _6115_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7650__29 _7650__29/A vssd1 vssd1 vccd1 vccd1 _8498_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _7855_/Q input14/X _6123_/B vssd1 vssd1 vccd1 vccd1 _6046_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7997_ _7997_/CLK _7997_/D vssd1 vssd1 vccd1 vccd1 _7997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8549_ _8551_/CLK _8549_/D vssd1 vssd1 vccd1 vccd1 _8549_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput207 _6074_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[8] sky130_fd_sc_hd__buf_2
X_4230_ _4230_/A vssd1 vssd1 vccd1 vccd1 _8374_/D sky130_fd_sc_hd__clkbuf_1
X_4161_ _8398_/Q _4160_/X _4161_/S vssd1 vssd1 vccd1 vccd1 _4162_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4092_ _4031_/X _8412_/Q _4094_/S vssd1 vssd1 vccd1 vccd1 _4093_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7920_ _7920_/CLK _7920_/D vssd1 vssd1 vccd1 vccd1 _7920_/Q sky130_fd_sc_hd__dfxtp_1
X_7851_ _7851_/CLK _7851_/D vssd1 vssd1 vccd1 vccd1 _7851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6802_ _6802_/A _6802_/B vssd1 vssd1 vccd1 vccd1 _7528_/B sky130_fd_sc_hd__xnor2_4
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4994_ _8151_/Q _4487_/X _4994_/S vssd1 vssd1 vccd1 vccd1 _4995_/A sky130_fd_sc_hd__mux2_1
X_7782_ _8543_/CLK _7782_/D vssd1 vssd1 vccd1 vccd1 _7782_/Q sky130_fd_sc_hd__dfxtp_1
X_3945_ _3945_/A vssd1 vssd1 vccd1 vccd1 _8500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3445_ clkbuf_0__3445_/X vssd1 vssd1 vccd1 vccd1 _7040_/A sky130_fd_sc_hd__clkbuf_4
X_6664_ _7728_/A _8002_/Q _6664_/S vssd1 vssd1 vccd1 vccd1 _6665_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5615_ _5615_/A vssd1 vssd1 vccd1 vccd1 _7977_/D sky130_fd_sc_hd__clkbuf_1
X_8403_ _8403_/CLK _8403_/D vssd1 vssd1 vccd1 vccd1 _8403_/Q sky130_fd_sc_hd__dfxtp_1
X_3876_ _7881_/Q _7882_/Q _7883_/Q _7884_/Q vssd1 vssd1 vccd1 vccd1 _6345_/B sky130_fd_sc_hd__or4_1
X_5546_ _5375_/X _8025_/Q _5546_/S vssd1 vssd1 vccd1 vccd1 _5547_/A sky130_fd_sc_hd__mux2_1
X_8334_ _8370_/CLK _8334_/D vssd1 vssd1 vccd1 vccd1 _8334_/Q sky130_fd_sc_hd__dfxtp_1
X_8265_ _8265_/CLK _8265_/D vssd1 vssd1 vccd1 vccd1 _8265_/Q sky130_fd_sc_hd__dfxtp_1
X_5477_ _5477_/A vssd1 vssd1 vccd1 vccd1 _8056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4428_ _5396_/A vssd1 vssd1 vccd1 vccd1 _4428_/X sky130_fd_sc_hd__buf_4
X_7216_ _7216_/A _7216_/B vssd1 vssd1 vccd1 vccd1 _7251_/A sky130_fd_sc_hd__xor2_1
Xclkbuf_0__3275_ _6652_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3275_/X sky130_fd_sc_hd__clkbuf_16
X_8196_ _8196_/CLK _8196_/D vssd1 vssd1 vccd1 vccd1 _8196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4359_ _4359_/A vssd1 vssd1 vccd1 vccd1 _8292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _6029_/A vssd1 vssd1 vccd1 vccd1 _6029_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3026_ clkbuf_0__3026_/X vssd1 vssd1 vccd1 vccd1 _6180__187/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_90 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5400_ _5399_/X _8094_/Q _5402_/S vssd1 vssd1 vccd1 vccd1 _5401_/A sky130_fd_sc_hd__mux2_1
X_6380_ _6331_/A _6377_/X _6379_/X _6367_/X vssd1 vssd1 vccd1 vccd1 _6380_/X sky130_fd_sc_hd__a31o_1
XFILLER_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3092_ clkbuf_0__3092_/X vssd1 vssd1 vccd1 vccd1 _6325__223/A sky130_fd_sc_hd__clkbuf_4
X_5331_ _5334_/C vssd1 vssd1 vccd1 vccd1 _5343_/B sky130_fd_sc_hd__inv_2
XFILLER_114_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8050_ _8050_/CLK _8050_/D vssd1 vssd1 vccd1 vccd1 _8050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5262_ _5343_/A vssd1 vssd1 vccd1 vccd1 _5262_/X sky130_fd_sc_hd__clkbuf_2
X_5193_ _5244_/A vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__buf_2
X_4213_ _8380_/Q _4193_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4214_/A sky130_fd_sc_hd__mux2_1
X_4144_ _6902_/A _4944_/B vssd1 vssd1 vccd1 vccd1 _4931_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4075_ _4075_/A vssd1 vssd1 vccd1 vccd1 _8419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7903_ _7903_/CLK _7903_/D vssd1 vssd1 vccd1 vccd1 _7903_/Q sky130_fd_sc_hd__dfxtp_1
X_7834_ _7834_/CLK _7834_/D vssd1 vssd1 vccd1 vccd1 _7834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7765_ _7765_/CLK _7765_/D vssd1 vssd1 vccd1 vccd1 _7765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4977_ _4933_/C _5014_/B _5014_/A vssd1 vssd1 vccd1 vccd1 _5733_/B sky130_fd_sc_hd__nand3b_4
XFILLER_11_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3928_ _3928_/A vssd1 vssd1 vccd1 vccd1 _8507_/D sky130_fd_sc_hd__clkbuf_1
X_7696_ _7696_/A _7696_/B _7696_/C _7696_/D vssd1 vssd1 vccd1 vccd1 _7698_/C sky130_fd_sc_hd__or4_1
XFILLER_109_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3428_ clkbuf_0__3428_/X vssd1 vssd1 vccd1 vccd1 _6948__415/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3859_ _8120_/Q _4038_/A _5034_/A _3858_/Y vssd1 vssd1 vccd1 vccd1 _3860_/D sky130_fd_sc_hd__a31o_1
X_6554__247 _6554__247/A vssd1 vssd1 vccd1 vccd1 _7925_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5529_ _5529_/A vssd1 vssd1 vccd1 vccd1 _8033_/D sky130_fd_sc_hd__clkbuf_1
X_8317_ _8317_/CLK _8317_/D vssd1 vssd1 vccd1 vccd1 _8317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8248_ _8248_/CLK _8248_/D vssd1 vssd1 vccd1 vccd1 _8248_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3258_ _6596_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3258_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3644_ clkbuf_0__3644_/X vssd1 vssd1 vccd1 vccd1 _7429__148/A sky130_fd_sc_hd__clkbuf_4
X_8179_ _8179_/CLK _8179_/D vssd1 vssd1 vccd1 vccd1 _8179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3575_ clkbuf_0__3575_/X vssd1 vssd1 vccd1 vccd1 _7297__113/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7182__100 _7181__99/A vssd1 vssd1 vccd1 vccd1 _8327_/CLK sky130_fd_sc_hd__inv_2
X_7084__521 _7088__525/A vssd1 vssd1 vccd1 vccd1 _8248_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4900_ _4803_/X _4898_/X _4899_/X vssd1 vssd1 vccd1 vccd1 _4900_/Y sky130_fd_sc_hd__o21ai_1
X_5880_ _6035_/A _5878_/B _5879_/X _7762_/Q vssd1 vssd1 vccd1 vccd1 _6161_/C sky130_fd_sc_hd__a31o_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4831_ _7936_/Q _4784_/X _4830_/X _4787_/X vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4762_ _4638_/X _4749_/X _4753_/X _4761_/X vssd1 vssd1 vccd1 vccd1 _4762_/X sky130_fd_sc_hd__a31o_1
X_7550_ _7550_/A _8460_/Q _7550_/C vssd1 vssd1 vccd1 vccd1 _7550_/X sky130_fd_sc_hd__and3_1
XFILLER_119_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4693_ _8141_/Q _8028_/Q _7924_/Q _7908_/Q _4655_/X _4656_/X vssd1 vssd1 vccd1 vccd1
+ _4693_/X sky130_fd_sc_hd__mux4_1
X_6501_ _8007_/Q _7892_/Q _6509_/S vssd1 vssd1 vccd1 vccd1 _6502_/A sky130_fd_sc_hd__mux2_1
X_6432_ _7866_/Q _6424_/X _6415_/X _6431_/X _6422_/X vssd1 vssd1 vccd1 vccd1 _7866_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8102_ _8102_/CLK _8102_/D vssd1 vssd1 vccd1 vccd1 _8102_/Q sky130_fd_sc_hd__dfxtp_1
X_6363_ _8550_/Q _6362_/X _6336_/X _6343_/X vssd1 vssd1 vccd1 vccd1 _6363_/X sky130_fd_sc_hd__a31o_1
XFILLER_115_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5314_ _5230_/X _5312_/X _5313_/X _5169_/A vssd1 vssd1 vccd1 vccd1 _5314_/X sky130_fd_sc_hd__o211a_1
XFILLER_114_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5245_ _8327_/Q _8048_/Q _5308_/S vssd1 vssd1 vccd1 vccd1 _5245_/X sky130_fd_sc_hd__mux2_1
X_8033_ _8033_/CLK _8033_/D vssd1 vssd1 vccd1 vccd1 _8033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5176_ _5176_/A vssd1 vssd1 vccd1 vccd1 _5349_/A sky130_fd_sc_hd__clkbuf_2
X_4127_ _4217_/B _8168_/Q vssd1 vssd1 vccd1 vccd1 _4627_/C sky130_fd_sc_hd__or2_1
X_4058_ _5787_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _4074_/S sky130_fd_sc_hd__or2_2
X_6560__251 _6564__255/A vssd1 vssd1 vccd1 vccd1 _7929_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7817_ _8543_/CLK _7817_/D vssd1 vssd1 vccd1 vccd1 _7817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7748_ _7644_/A _7646_/B _7743_/X _7729_/A vssd1 vssd1 vccd1 vccd1 _7748_/X sky130_fd_sc_hd__a31o_1
X_7679_ _7680_/A _7679_/B vssd1 vssd1 vccd1 vccd1 _8522_/D sky130_fd_sc_hd__nor2_1
XFILLER_118_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6873__372 _6873__372/A vssd1 vssd1 vccd1 vccd1 _8086_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7049__493 _7049__493/A vssd1 vssd1 vccd1 vccd1 _8220_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5030_ _5030_/A vssd1 vssd1 vccd1 vccd1 _8136_/D sky130_fd_sc_hd__clkbuf_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6981_ _6987_/A vssd1 vssd1 vccd1 vccd1 _6981_/X sky130_fd_sc_hd__buf_1
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5932_ _5932_/A _5932_/B vssd1 vssd1 vccd1 vccd1 _5933_/A sky130_fd_sc_hd__or2_4
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5863_ _4151_/X _7769_/Q _5869_/S vssd1 vssd1 vccd1 vccd1 _5864_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5794_ _5794_/A vssd1 vssd1 vccd1 vccd1 _7843_/D sky130_fd_sc_hd__clkbuf_1
X_4814_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4883_/S sky130_fd_sc_hd__clkbuf_2
X_7602_ _7601_/X _6867_/C _7597_/X vssd1 vssd1 vccd1 vccd1 _7602_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7533_ _6440_/A _6793_/B _6800_/B _7727_/B vssd1 vssd1 vccd1 vccd1 _7533_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4745_ _4712_/X _4743_/X _4744_/X _4690_/X vssd1 vssd1 vccd1 vccd1 _8184_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7464_ _7482_/A vssd1 vssd1 vccd1 vccd1 _7464_/X sky130_fd_sc_hd__buf_1
X_4676_ _8252_/Q _8037_/Q _7989_/Q _7941_/Q _4646_/A _4649_/A vssd1 vssd1 vccd1 vccd1
+ _4676_/X sky130_fd_sc_hd__mux4_1
X_7395_ _7395_/A vssd1 vssd1 vccd1 vccd1 _7395_/X sky130_fd_sc_hd__buf_1
X_6415_ _6437_/A vssd1 vssd1 vccd1 vccd1 _6415_/X sky130_fd_sc_hd__clkbuf_2
X_6346_ _6517_/A _6417_/A vssd1 vssd1 vccd1 vccd1 _6521_/B sky130_fd_sc_hd__and2b_1
XFILLER_103_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput107 wbs_we_i vssd1 vssd1 vccd1 vccd1 _6269_/C sky130_fd_sc_hd__buf_6
X_8016_ _8531_/CLK _8016_/D vssd1 vssd1 vccd1 vccd1 _8016_/Q sky130_fd_sc_hd__dfxtp_1
X_6277_ _8359_/Q vssd1 vssd1 vccd1 vccd1 _7356_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5228_ _8223_/Q _5270_/A _5214_/X _8207_/Q _5092_/A vssd1 vssd1 vccd1 vccd1 _5228_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__3026_ _6178_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3026_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_111_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5159_ _5079_/X _5158_/X _5083_/X vssd1 vssd1 vccd1 vccd1 _5159_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3274_ clkbuf_0__3274_/X vssd1 vssd1 vccd1 vccd1 _6649__308/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6567__257 _6568__258/A vssd1 vssd1 vccd1 vccd1 _7935_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4530_ _4530_/A vssd1 vssd1 vccd1 vccd1 _8229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4461_ _4394_/X _8254_/Q _4463_/S vssd1 vssd1 vccd1 vccd1 _4462_/A sky130_fd_sc_hd__mux2_1
X_6200_ _6235_/A vssd1 vssd1 vccd1 vccd1 _6200_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4392_ _4391_/X _8279_/Q _4398_/S vssd1 vssd1 vccd1 vccd1 _4393_/A sky130_fd_sc_hd__mux2_1
X_6131_ _6131_/A _6140_/B vssd1 vssd1 vccd1 vccd1 _6131_/X sky130_fd_sc_hd__and2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6062_ _7784_/Q _6066_/B vssd1 vssd1 vccd1 vccd1 _6062_/X sky130_fd_sc_hd__or2_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5013_ _5013_/A vssd1 vssd1 vccd1 vccd1 _8143_/D sky130_fd_sc_hd__clkbuf_1
X_7097__531 _7099__533/A vssd1 vssd1 vccd1 vccd1 _8258_/CLK sky130_fd_sc_hd__inv_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5915_ _7644_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__or2_1
XFILLER_81_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5846_ _5846_/A vssd1 vssd1 vccd1 vccd1 _7777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5777_ _5611_/X _7850_/Q _5779_/S vssd1 vssd1 vccd1 vccd1 _5778_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3644_ _7426_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3644_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__3575_ _7294_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3575_/X sky130_fd_sc_hd__clkbuf_16
X_8496_ _8496_/CLK _8496_/D vssd1 vssd1 vccd1 vccd1 _8496_/Q sky130_fd_sc_hd__dfxtp_1
X_4728_ _4766_/B vssd1 vssd1 vccd1 vccd1 _4880_/S sky130_fd_sc_hd__buf_2
X_7516_ _8549_/Q _7551_/B vssd1 vssd1 vccd1 vccd1 _7519_/A sky130_fd_sc_hd__xor2_1
X_4659_ _4683_/B _4669_/B vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__or2_2
X_7378_ _8129_/Q _7364_/A _7366_/X _7377_/X _7371_/X vssd1 vssd1 vccd1 vccd1 _8366_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6329_ _6329_/A vssd1 vssd1 vccd1 vccd1 _7742_/B sky130_fd_sc_hd__buf_2
XFILLER_107_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3257_ clkbuf_0__3257_/X vssd1 vssd1 vccd1 vccd1 _6595__280/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6946__413 _6946__413/A vssd1 vssd1 vccd1 vccd1 _8137_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3961_ _8458_/Q _3954_/X _3973_/S vssd1 vssd1 vccd1 vccd1 _3962_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5700_ _5700_/A vssd1 vssd1 vccd1 vccd1 _7933_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3461_ clkbuf_0__3461_/X vssd1 vssd1 vccd1 vccd1 _7109__541/A sky130_fd_sc_hd__clkbuf_4
X_3892_ _3892_/A vssd1 vssd1 vccd1 vccd1 _8519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6680_ _5943_/A _8009_/Q _6682_/S vssd1 vssd1 vccd1 vccd1 _6681_/A sky130_fd_sc_hd__mux2_1
X_5631_ _5611_/X _7962_/Q _5633_/S vssd1 vssd1 vccd1 vccd1 _5632_/A sky130_fd_sc_hd__mux2_1
X_5562_ _5396_/X _7995_/Q _5567_/S vssd1 vssd1 vccd1 vccd1 _5563_/A sky130_fd_sc_hd__mux2_1
X_8350_ _8358_/CLK _8350_/D vssd1 vssd1 vccd1 vccd1 _8350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8281_ _8281_/CLK _8281_/D vssd1 vssd1 vccd1 vccd1 _8281_/Q sky130_fd_sc_hd__dfxtp_1
X_4513_ _8236_/Q _4465_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4514_/A sky130_fd_sc_hd__mux2_1
X_7301_ _7334_/A vssd1 vssd1 vccd1 vccd1 _7301_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5493_ _5493_/A vssd1 vssd1 vccd1 vccd1 _8049_/D sky130_fd_sc_hd__clkbuf_1
X_7232_ _8351_/Q _7232_/B _7232_/C vssd1 vssd1 vccd1 vccd1 _7329_/A sky130_fd_sc_hd__nand3_2
X_4444_ _8106_/Q vssd1 vssd1 vccd1 vccd1 _4444_/X sky130_fd_sc_hd__buf_2
X_4375_ _4490_/A _5428_/A vssd1 vssd1 vccd1 vccd1 _4398_/S sky130_fd_sc_hd__or2_2
X_6886__382 _6887__383/A vssd1 vssd1 vccd1 vccd1 _8096_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6114_/A vssd1 vssd1 vccd1 vccd1 _6153_/B sky130_fd_sc_hd__clkbuf_4
X_6045_ _6034_/X _6039_/X _6042_/X _6044_/X vssd1 vssd1 vccd1 vccd1 _6045_/X sky130_fd_sc_hd__o211a_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7996_ _7996_/CLK _7996_/D vssd1 vssd1 vccd1 vccd1 _7996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6878_ _6890_/A vssd1 vssd1 vccd1 vccd1 _6878_/X sky130_fd_sc_hd__buf_1
X_5829_ _7827_/Q _5396_/A _5833_/S vssd1 vssd1 vccd1 vccd1 _5830_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8548_ _8548_/CLK _8548_/D vssd1 vssd1 vccd1 vccd1 _8548_/Q sky130_fd_sc_hd__dfxtp_1
X_6750__346 _6754__350/A vssd1 vssd1 vccd1 vccd1 _8056_/CLK sky130_fd_sc_hd__inv_2
X_8479_ _8479_/CLK _8479_/D vssd1 vssd1 vccd1 vccd1 _8479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3309_ clkbuf_0__3309_/X vssd1 vssd1 vccd1 vccd1 _6730__330/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput208 _6079_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_114_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7180__98 _7181__99/A vssd1 vssd1 vccd1 vccd1 _8325_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4160_ _8109_/Q vssd1 vssd1 vccd1 vccd1 _4160_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4091_ _4091_/A vssd1 vssd1 vccd1 vccd1 _8413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7850_ _7850_/CLK _7850_/D vssd1 vssd1 vccd1 vccd1 _7850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6801_ _8473_/Q vssd1 vssd1 vccd1 vccd1 _6802_/A sky130_fd_sc_hd__clkinv_2
XFILLER_63_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ _4993_/A vssd1 vssd1 vccd1 vccd1 _8152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7781_ _8355_/CLK _7781_/D vssd1 vssd1 vccd1 vccd1 _7781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3944_ _3899_/X _8500_/Q _3946_/S vssd1 vssd1 vccd1 vccd1 _3945_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3444_ clkbuf_0__3444_/X vssd1 vssd1 vccd1 vccd1 _7023__472/A sky130_fd_sc_hd__clkbuf_4
X_6663_ _6663_/A vssd1 vssd1 vccd1 vccd1 _8001_/D sky130_fd_sc_hd__clkbuf_1
X_3875_ _8062_/Q _6352_/A vssd1 vssd1 vccd1 vccd1 _6355_/A sky130_fd_sc_hd__nand2_1
X_8402_ _8402_/CLK _8402_/D vssd1 vssd1 vccd1 vccd1 _8402_/Q sky130_fd_sc_hd__dfxtp_1
X_5614_ _5566_/X _7977_/Q _5614_/S vssd1 vssd1 vccd1 vccd1 _5615_/A sky130_fd_sc_hd__mux2_1
X_8333_ _8370_/CLK _8333_/D vssd1 vssd1 vccd1 vccd1 _8333_/Q sky130_fd_sc_hd__dfxtp_2
X_5545_ _5545_/A vssd1 vssd1 vccd1 vccd1 _8026_/D sky130_fd_sc_hd__clkbuf_1
X_5476_ _3975_/X _8056_/Q _5480_/S vssd1 vssd1 vccd1 vccd1 _5477_/A sky130_fd_sc_hd__mux2_1
X_8264_ _8264_/CLK _8264_/D vssd1 vssd1 vccd1 vccd1 _8264_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3274_ _6646_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3274_/X sky130_fd_sc_hd__clkbuf_16
X_8195_ _8195_/CLK _8195_/D vssd1 vssd1 vccd1 vccd1 _8195_/Q sky130_fd_sc_hd__dfxtp_1
X_7215_ _7272_/B _7272_/C vssd1 vssd1 vccd1 vccd1 _7216_/B sky130_fd_sc_hd__nand2_1
X_4427_ _8111_/Q vssd1 vssd1 vccd1 vccd1 _5396_/A sky130_fd_sc_hd__buf_6
X_7146_ _7146_/A vssd1 vssd1 vccd1 vccd1 _7146_/X sky130_fd_sc_hd__buf_1
XFILLER_113_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4358_ _4275_/X _8292_/Q _4366_/S vssd1 vssd1 vccd1 vccd1 _4359_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4289_ _4289_/A vssd1 vssd1 vccd1 vccd1 _4289_/X sky130_fd_sc_hd__clkbuf_2
X_7077_ _7077_/A vssd1 vssd1 vccd1 vccd1 _7077_/X sky130_fd_sc_hd__buf_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6028_ _8016_/Q _6030_/B vssd1 vssd1 vccd1 vccd1 _6029_/A sky130_fd_sc_hd__and2_2
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7979_ _7979_/CLK _7979_/D vssd1 vssd1 vccd1 vccd1 _7979_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3025_ clkbuf_0__3025_/X vssd1 vssd1 vccd1 vccd1 _6177__185/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7043__488 _7043__488/A vssd1 vssd1 vccd1 vccd1 _8215_/CLK sky130_fd_sc_hd__inv_2
X_7480__14 _7481__15/A vssd1 vssd1 vccd1 vccd1 _8446_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_80 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_91 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8575__222 vssd1 vssd1 vccd1 vccd1 _8575__222/HI core1Index[2] sky130_fd_sc_hd__conb_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7447__162 _7447__162/A vssd1 vssd1 vccd1 vccd1 _8419_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3091_ clkbuf_0__3091_/X vssd1 vssd1 vccd1 vccd1 _6321__220/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5330_ _5330_/A vssd1 vssd1 vccd1 vccd1 _5334_/C sky130_fd_sc_hd__clkbuf_2
X_5261_ _8127_/Q _5041_/A _5349_/A _5260_/X _5107_/A vssd1 vssd1 vccd1 vccd1 _5261_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4212_ _4212_/A vssd1 vssd1 vccd1 vccd1 _8381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7000_ _7006_/A vssd1 vssd1 vccd1 vccd1 _7000_/X sky130_fd_sc_hd__buf_1
X_5192_ _5192_/A vssd1 vssd1 vccd1 vccd1 _5244_/A sky130_fd_sc_hd__clkbuf_2
X_4143_ _8187_/Q _7676_/B vssd1 vssd1 vccd1 vccd1 _4944_/B sky130_fd_sc_hd__and2_1
XFILLER_110_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4074_ _4035_/X _8419_/Q _4074_/S vssd1 vssd1 vccd1 vccd1 _4075_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7902_ _7902_/CLK _7902_/D vssd1 vssd1 vccd1 vccd1 _7902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7833_ _7833_/CLK _7833_/D vssd1 vssd1 vccd1 vccd1 _7833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7764_ _7764_/CLK _7764_/D vssd1 vssd1 vccd1 vccd1 _7764_/Q sky130_fd_sc_hd__dfxtp_1
X_4976_ _4976_/A vssd1 vssd1 vccd1 vccd1 _8159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6300__202 _6303__205/A vssd1 vssd1 vccd1 vccd1 _7832_/CLK sky130_fd_sc_hd__inv_2
X_7695_ _7695_/A vssd1 vssd1 vccd1 vccd1 _8530_/D sky130_fd_sc_hd__clkbuf_1
X_3927_ _3902_/X _8507_/Q _3927_/S vssd1 vssd1 vccd1 vccd1 _3928_/A sky130_fd_sc_hd__mux2_1
X_6646_ _6652_/A vssd1 vssd1 vccd1 vccd1 _6646_/X sky130_fd_sc_hd__buf_1
X_3858_ _5035_/B _3849_/B _3846_/Y vssd1 vssd1 vccd1 vccd1 _3858_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6577_ _6583_/A vssd1 vssd1 vccd1 vccd1 _6577_/X sky130_fd_sc_hd__buf_1
XFILLER_118_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5528_ _5375_/X _8033_/Q _5528_/S vssd1 vssd1 vccd1 vccd1 _5529_/A sky130_fd_sc_hd__mux2_1
X_8316_ _8316_/CLK _8316_/D vssd1 vssd1 vccd1 vccd1 _8316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5459_ _5459_/A vssd1 vssd1 vccd1 vccd1 _8067_/D sky130_fd_sc_hd__clkbuf_1
X_8247_ _8247_/CLK _8247_/D vssd1 vssd1 vccd1 vccd1 _8247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3257_ _6590_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3257_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3643_ clkbuf_0__3643_/X vssd1 vssd1 vccd1 vccd1 _7422__142/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8178_ _8178_/CLK _8178_/D vssd1 vssd1 vccd1 vccd1 _8178_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3574_ clkbuf_0__3574_/X vssd1 vssd1 vccd1 vccd1 _7290__107/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7091__526 _7093__528/A vssd1 vssd1 vccd1 vccd1 _8253_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_2_0_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_4830_ _7984_/Q _8032_/Q _4883_/S vssd1 vssd1 vccd1 vccd1 _4830_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _4755_/X _4757_/X _4760_/X _4740_/X _4684_/X vssd1 vssd1 vccd1 vccd1 _4761_/X
+ sky130_fd_sc_hd__o221a_2
X_6500_ _6511_/A vssd1 vssd1 vccd1 vccd1 _6509_/S sky130_fd_sc_hd__clkbuf_2
X_4692_ _8096_/Q _8088_/Q _7916_/Q _8157_/Q _4810_/S _4649_/X vssd1 vssd1 vccd1 vccd1
+ _4692_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6431_ _7727_/B _6434_/B _6431_/C vssd1 vssd1 vccd1 vccd1 _6431_/X sky130_fd_sc_hd__and3_1
X_7126__54 _7127__55/A vssd1 vssd1 vccd1 vccd1 _8281_/CLK sky130_fd_sc_hd__inv_2
X_6362_ _6362_/A vssd1 vssd1 vccd1 vccd1 _6362_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5313_ _8496_/Q _5232_/X _5207_/A _8512_/Q vssd1 vssd1 vccd1 vccd1 _5313_/X sky130_fd_sc_hd__o22a_1
X_8101_ _8101_/CLK _8101_/D vssd1 vssd1 vccd1 vccd1 _8101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5244_ _5244_/A vssd1 vssd1 vccd1 vccd1 _5306_/A sky130_fd_sc_hd__buf_2
X_8032_ _8032_/CLK _8032_/D vssd1 vssd1 vccd1 vccd1 _8032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5175_ _3899_/X _5038_/X _5174_/X _5111_/X vssd1 vssd1 vccd1 vccd1 _8129_/D sky130_fd_sc_hd__o211a_1
XFILLER_96_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4126_ _8173_/Q vssd1 vssd1 vccd1 vccd1 _4217_/B sky130_fd_sc_hd__inv_2
XFILLER_29_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4057_ _4301_/A _4057_/B _4256_/C vssd1 vssd1 vccd1 vccd1 _5464_/B sky130_fd_sc_hd__or3_2
XFILLER_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7816_ _8543_/CLK _7816_/D vssd1 vssd1 vccd1 vccd1 _7816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ _4959_/A _5733_/A vssd1 vssd1 vccd1 vccd1 _4975_/S sky130_fd_sc_hd__nor2_2
X_7747_ _7747_/A _7747_/B vssd1 vssd1 vccd1 vccd1 _7747_/Y sky130_fd_sc_hd__nand2_2
X_7678_ _7678_/A vssd1 vssd1 vccd1 vccd1 _8521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7668__44 _7669__45/A vssd1 vssd1 vccd1 vccd1 _8513_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3309_ _6725_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3309_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6307__208 _6309__210/A vssd1 vssd1 vccd1 vccd1 _7838_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6650__309 _6651__310/A vssd1 vssd1 vccd1 vccd1 _7995_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6880__377 _6881__378/A vssd1 vssd1 vccd1 vccd1 _8091_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5931_ _5931_/A vssd1 vssd1 vccd1 vccd1 _5931_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5862_ _5862_/A vssd1 vssd1 vccd1 vccd1 _7770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5793_ _7843_/Q _4283_/A _5797_/S vssd1 vssd1 vccd1 vccd1 _5794_/A sky130_fd_sc_hd__mux2_1
X_4813_ _4955_/B _4810_/X _4812_/X vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__o21a_1
X_7601_ _7614_/A vssd1 vssd1 vccd1 vccd1 _7601_/X sky130_fd_sc_hd__clkbuf_2
X_7532_ _8536_/Q _7532_/B _7532_/C vssd1 vssd1 vccd1 vccd1 _7532_/X sky130_fd_sc_hd__and3_1
X_4744_ _5396_/A _4764_/B vssd1 vssd1 vccd1 vccd1 _4744_/X sky130_fd_sc_hd__or2_1
XFILLER_107_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4675_ _8150_/Q _8105_/Q _7997_/Q _8342_/Q _4646_/A _4674_/X vssd1 vssd1 vccd1 vccd1
+ _4675_/X sky130_fd_sc_hd__mux4_1
X_7463_ _7494_/A vssd1 vssd1 vccd1 vccd1 _7463_/X sky130_fd_sc_hd__buf_1
X_6414_ _6331_/X _6412_/X _6413_/X vssd1 vssd1 vccd1 vccd1 _7862_/D sky130_fd_sc_hd__a21o_1
X_6345_ _7880_/Q _6345_/B _7879_/Q vssd1 vssd1 vccd1 vccd1 _6461_/D sky130_fd_sc_hd__or3b_2
X_6293__197 _6294__198/A vssd1 vssd1 vccd1 vccd1 _7827_/CLK sky130_fd_sc_hd__inv_2
X_6276_ _7298_/A vssd1 vssd1 vccd1 vccd1 _7359_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5227_ _5227_/A vssd1 vssd1 vccd1 vccd1 _5270_/A sky130_fd_sc_hd__clkbuf_2
X_8015_ _8531_/CLK _8015_/D vssd1 vssd1 vccd1 vccd1 _8015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3025_ _6172_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3025_/X sky130_fd_sc_hd__clkbuf_16
X_5158_ _8439_/Q _8431_/Q _7834_/Q _8447_/Q _5066_/X _5080_/X vssd1 vssd1 vccd1 vccd1
+ _5158_/X sky130_fd_sc_hd__mux4_2
XFILLER_96_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4109_ _4109_/A vssd1 vssd1 vccd1 vccd1 _8405_/D sky130_fd_sc_hd__clkbuf_1
X_5089_ _8511_/Q _8260_/Q _8244_/Q _8284_/Q _5087_/X _5088_/X vssd1 vssd1 vccd1 vccd1
+ _5090_/B sky130_fd_sc_hd__mux4_2
XFILLER_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3273_ clkbuf_0__3273_/X vssd1 vssd1 vccd1 vccd1 _6645__305/A sky130_fd_sc_hd__clkbuf_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6714__317 _6716__319/A vssd1 vssd1 vccd1 vccd1 _8027_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _4460_/A vssd1 vssd1 vccd1 vccd1 _8255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4391_ _8490_/Q vssd1 vssd1 vccd1 vccd1 _4391_/X sky130_fd_sc_hd__clkbuf_2
X_6130_ _7801_/Q _6122_/X _6126_/X _6129_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6130_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _7859_/Q input30/X _6072_/S vssd1 vssd1 vccd1 vccd1 _6061_/X sky130_fd_sc_hd__mux2_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _8143_/Q _4487_/X _5012_/S vssd1 vssd1 vccd1 vccd1 _5013_/A sky130_fd_sc_hd__mux2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7662__39 _7663__40/A vssd1 vssd1 vccd1 vccd1 _8508_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6963_ _6975_/A vssd1 vssd1 vccd1 vccd1 _6963_/X sky130_fd_sc_hd__buf_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5914_ _5914_/A vssd1 vssd1 vccd1 vccd1 _5914_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5845_ _4151_/X _7777_/Q _5851_/S vssd1 vssd1 vccd1 vccd1 _5846_/A sky130_fd_sc_hd__mux2_1
X_8555__253 vssd1 vssd1 vccd1 vccd1 partID[4] _8555__253/LO sky130_fd_sc_hd__conb_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5776_ _5776_/A vssd1 vssd1 vccd1 vccd1 _7851_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3643_ _7420_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3643_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__3574_ _7288_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3574_/X sky130_fd_sc_hd__clkbuf_16
X_4727_ _4782_/A vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__clkbuf_2
X_7515_ _7550_/A _7548_/S vssd1 vssd1 vccd1 vccd1 _7551_/B sky130_fd_sc_hd__xor2_2
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8495_ _8527_/CLK _8495_/D vssd1 vssd1 vccd1 vccd1 _8495_/Q sky130_fd_sc_hd__dfxtp_2
X_4658_ _8171_/Q _4658_/B vssd1 vssd1 vccd1 vccd1 _4669_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput90 wbs_data_i[28] vssd1 vssd1 vccd1 vccd1 _5963_/A sky130_fd_sc_hd__buf_4
XFILLER_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7377_ _8366_/Q _7377_/B vssd1 vssd1 vccd1 vccd1 _7377_/X sky130_fd_sc_hd__or2_1
X_4589_ _4589_/A vssd1 vssd1 vccd1 vccd1 _8204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7106__539 _7106__539/A vssd1 vssd1 vccd1 vccd1 _8266_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6328_ _6328_/A vssd1 vssd1 vccd1 vccd1 _6328_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6259_ _6259_/A vssd1 vssd1 vccd1 vccd1 _7815_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3256_ clkbuf_0__3256_/X vssd1 vssd1 vccd1 vccd1 _6626_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6573__262 _6574__263/A vssd1 vssd1 vccd1 vccd1 _7940_/CLK sky130_fd_sc_hd__inv_2
X_7441__157 _7441__157/A vssd1 vssd1 vccd1 vccd1 _8414_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3960_ _3982_/S vssd1 vssd1 vccd1 vccd1 _3973_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_63_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3460_ clkbuf_0__3460_/X vssd1 vssd1 vccd1 vccd1 _7106__539/A sky130_fd_sc_hd__clkbuf_4
X_3891_ _3831_/X _8519_/Q _3903_/S vssd1 vssd1 vccd1 vccd1 _3892_/A sky130_fd_sc_hd__mux2_1
X_5630_ _5630_/A vssd1 vssd1 vccd1 vccd1 _7963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5561_ _5561_/A vssd1 vssd1 vccd1 vccd1 _7996_/D sky130_fd_sc_hd__clkbuf_1
X_5492_ _8049_/Q _4289_/A _5492_/S vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__mux2_1
X_4512_ _4529_/S vssd1 vssd1 vccd1 vccd1 _4523_/S sky130_fd_sc_hd__buf_2
X_8280_ _8280_/CLK _8280_/D vssd1 vssd1 vccd1 vccd1 _8280_/Q sky130_fd_sc_hd__dfxtp_1
X_7300_ _7298_/A _7285_/B _7303_/B vssd1 vssd1 vccd1 vccd1 _7334_/A sky130_fd_sc_hd__a21o_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7231_ _7280_/A _7281_/A _7280_/B _7281_/B vssd1 vssd1 vccd1 vccd1 _7251_/C sky130_fd_sc_hd__and4_1
XFILLER_104_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4443_ _4443_/A vssd1 vssd1 vccd1 vccd1 _8262_/D sky130_fd_sc_hd__clkbuf_1
X_4374_ _8495_/Q vssd1 vssd1 vccd1 vccd1 _4374_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6113_ _6095_/X _6111_/X _6112_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6113_/X sky130_fd_sc_hd__o211a_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6044_ _6063_/A vssd1 vssd1 vccd1 vccd1 _6044_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7995_ _7995_/CLK _7995_/D vssd1 vssd1 vccd1 vccd1 _7995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8592__239 vssd1 vssd1 vccd1 vccd1 _8592__239/HI partID[1] sky130_fd_sc_hd__conb_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3658_ clkbuf_0__3658_/X vssd1 vssd1 vccd1 vccd1 _7651__30/A sky130_fd_sc_hd__clkbuf_4
X_6877_ _6925_/A vssd1 vssd1 vccd1 vccd1 _6877_/X sky130_fd_sc_hd__buf_1
XFILLER_22_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5828_ _5828_/A vssd1 vssd1 vccd1 vccd1 _7828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5759_ _7906_/Q _5399_/A _5761_/S vssd1 vssd1 vccd1 vccd1 _5760_/A sky130_fd_sc_hd__mux2_1
X_8547_ _8550_/CLK _8547_/D vssd1 vssd1 vccd1 vccd1 _8547_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8478_ _8479_/CLK _8478_/D vssd1 vssd1 vccd1 vccd1 _8478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3308_ clkbuf_0__3308_/X vssd1 vssd1 vccd1 vccd1 _6749_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6766__354 _6766__354/A vssd1 vssd1 vccd1 vccd1 _8067_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6727__327 _6727__327/A vssd1 vssd1 vccd1 vccd1 _8037_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4090_ _4027_/X _8413_/Q _4094_/S vssd1 vssd1 vccd1 vccd1 _4091_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ _8540_/Q _6800_/B vssd1 vssd1 vccd1 vccd1 _6808_/B sky130_fd_sc_hd__xor2_1
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4992_ _8152_/Q _4484_/X _4994_/S vssd1 vssd1 vccd1 vccd1 _4993_/A sky130_fd_sc_hd__mux2_1
X_7780_ _8355_/CLK _7780_/D vssd1 vssd1 vccd1 vccd1 _7780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3943_ _3943_/A vssd1 vssd1 vccd1 vccd1 _8501_/D sky130_fd_sc_hd__clkbuf_1
X_6731_ _6737_/A vssd1 vssd1 vccd1 vccd1 _6731_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3443_ clkbuf_0__3443_/X vssd1 vssd1 vccd1 vccd1 _7019__469/A sky130_fd_sc_hd__clkbuf_4
X_6662_ _5926_/A _8001_/Q _6664_/S vssd1 vssd1 vccd1 vccd1 _6663_/A sky130_fd_sc_hd__mux2_1
X_3874_ _7900_/Q _7899_/Q vssd1 vssd1 vccd1 vccd1 _6352_/A sky130_fd_sc_hd__or2_1
X_8401_ _8401_/CLK _8401_/D vssd1 vssd1 vccd1 vccd1 _8401_/Q sky130_fd_sc_hd__dfxtp_1
X_5613_ _5613_/A vssd1 vssd1 vccd1 vccd1 _7978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8332_ _8332_/CLK _8332_/D vssd1 vssd1 vccd1 vccd1 _8332_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3411_ _6896_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3411_/X sky130_fd_sc_hd__clkbuf_16
X_5544_ _5399_/X _8026_/Q _5546_/S vssd1 vssd1 vccd1 vccd1 _5545_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5475_ _5475_/A vssd1 vssd1 vccd1 vccd1 _8057_/D sky130_fd_sc_hd__clkbuf_1
X_8263_ _8263_/CLK _8263_/D vssd1 vssd1 vccd1 vccd1 _8263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3273_ _6640_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3273_/X sky130_fd_sc_hd__clkbuf_16
X_4426_ _4426_/A vssd1 vssd1 vccd1 vccd1 _8267_/D sky130_fd_sc_hd__clkbuf_1
X_8194_ _8194_/CLK _8194_/D vssd1 vssd1 vccd1 vccd1 _8194_/Q sky130_fd_sc_hd__dfxtp_1
X_7214_ _8349_/Q _7227_/A _7236_/A _7232_/B _8350_/Q vssd1 vssd1 vccd1 vccd1 _7272_/C
+ sky130_fd_sc_hd__a41o_1
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4357_ _4372_/S vssd1 vssd1 vccd1 vccd1 _4366_/S sky130_fd_sc_hd__buf_2
XFILLER_59_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4288_ _4288_/A vssd1 vssd1 vccd1 vccd1 _8321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _6027_/A vssd1 vssd1 vccd1 vccd1 _6027_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7978_ _7978_/CLK _7978_/D vssd1 vssd1 vccd1 vccd1 _7978_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3024_ clkbuf_0__3024_/X vssd1 vssd1 vccd1 vccd1 _6170__179/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6163_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_70 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_92 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_81 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3090_ clkbuf_0__3090_/X vssd1 vssd1 vccd1 vccd1 _6315__215/A sky130_fd_sc_hd__clkbuf_4
X_5260_ _5350_/B _5235_/X _5243_/X _5259_/X vssd1 vssd1 vccd1 vccd1 _5260_/X sky130_fd_sc_hd__a31o_2
XFILLER_114_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4211_ _8381_/Q _4190_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5191_ _8280_/Q _5180_/X _5264_/A _5187_/X _5190_/X vssd1 vssd1 vccd1 vccd1 _5191_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4142_ _4125_/X _4131_/X _4138_/Y _4141_/X vssd1 vssd1 vccd1 vccd1 _7676_/B sky130_fd_sc_hd__a211o_1
XFILLER_95_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4073_ _4073_/A vssd1 vssd1 vccd1 vccd1 _8420_/D sky130_fd_sc_hd__clkbuf_1
X_6959__424 _6960__425/A vssd1 vssd1 vccd1 vccd1 _8148_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7901_ _8543_/CLK _7901_/D vssd1 vssd1 vccd1 vccd1 _7901_/Q sky130_fd_sc_hd__dfxtp_1
X_6627__291 _6628__292/A vssd1 vssd1 vccd1 vccd1 _7977_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8487_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7832_ _7832_/CLK _7832_/D vssd1 vssd1 vccd1 vccd1 _7832_/Q sky130_fd_sc_hd__dfxtp_1
X_7763_ _7763_/CLK _7763_/D vssd1 vssd1 vccd1 vccd1 _7763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4975_ _8159_/Q _4487_/X _4975_/S vssd1 vssd1 vccd1 vccd1 _4976_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3926_ _3926_/A vssd1 vssd1 vccd1 vccd1 _8508_/D sky130_fd_sc_hd__clkbuf_1
X_7694_ _7719_/A _8524_/Q vssd1 vssd1 vccd1 vccd1 _7695_/A sky130_fd_sc_hd__and2_1
XFILLER_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3857_ _8119_/Q vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5527_ _5527_/A vssd1 vssd1 vccd1 vccd1 _8034_/D sky130_fd_sc_hd__clkbuf_1
X_6966__428 _6968__430/A vssd1 vssd1 vccd1 vccd1 _8152_/CLK sky130_fd_sc_hd__inv_2
X_8315_ _8315_/CLK _8315_/D vssd1 vssd1 vccd1 vccd1 _8315_/Q sky130_fd_sc_hd__dfxtp_1
X_8246_ _8246_/CLK _8246_/D vssd1 vssd1 vccd1 vccd1 _8246_/Q sky130_fd_sc_hd__dfxtp_1
X_5458_ _8067_/Q _4190_/X _5462_/S vssd1 vssd1 vccd1 vccd1 _5459_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3256_ _6589_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3256_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3642_ clkbuf_0__3642_/X vssd1 vssd1 vccd1 vccd1 _7419__140/A sky130_fd_sc_hd__clkbuf_4
X_5389_ _5389_/A vssd1 vssd1 vccd1 vccd1 _8098_/D sky130_fd_sc_hd__clkbuf_1
X_4409_ _4409_/A vssd1 vssd1 vccd1 vccd1 _8273_/D sky130_fd_sc_hd__clkbuf_1
X_8177_ _8177_/CLK _8177_/D vssd1 vssd1 vccd1 vccd1 _8177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7128_ _7146_/A vssd1 vssd1 vccd1 vccd1 _7128_/X sky130_fd_sc_hd__buf_1
XFILLER_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7059_ _7083_/A vssd1 vssd1 vccd1 vccd1 _7059_/X sky130_fd_sc_hd__buf_1
XFILLER_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8598__245 vssd1 vssd1 vccd1 vccd1 _8598__245/HI partID[13] sky130_fd_sc_hd__conb_1
XFILLER_27_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3022_ clkbuf_0__3022_/X vssd1 vssd1 vccd1 vccd1 _6589_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4758_/X _4759_/X _4760_/S vssd1 vssd1 vccd1 vccd1 _4760_/X sky130_fd_sc_hd__mux2_1
X_4691_ _4418_/X _4629_/X _4688_/X _4690_/X vssd1 vssd1 vccd1 vccd1 _8186_/D sky130_fd_sc_hd__o211a_1
X_6430_ _8539_/Q vssd1 vssd1 vccd1 vccd1 _7727_/B sky130_fd_sc_hd__clkbuf_4
X_6361_ _7854_/Q _6328_/X _6360_/X vssd1 vssd1 vccd1 vccd1 _7854_/D sky130_fd_sc_hd__a21o_1
X_5312_ _8038_/Q _8065_/Q _5312_/S vssd1 vssd1 vccd1 vccd1 _5312_/X sky130_fd_sc_hd__mux2_1
X_8100_ _8100_/CLK _8100_/D vssd1 vssd1 vccd1 vccd1 _8100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5243_ _5293_/A _5243_/B _5243_/C vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__or3_1
X_8031_ _8031_/CLK _8031_/D vssd1 vssd1 vccd1 vccd1 _8031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5174_ _8129_/Q _5040_/X _5348_/A _5173_/X _5107_/X vssd1 vssd1 vccd1 vccd1 _5174_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4125_ _4125_/A _4944_/A _8168_/Q vssd1 vssd1 vccd1 vccd1 _4125_/X sky130_fd_sc_hd__or3b_1
XFILLER_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4056_ _4056_/A vssd1 vssd1 vccd1 vccd1 _8427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7815_ _8543_/CLK _7815_/D vssd1 vssd1 vccd1 vccd1 _7815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7746_ _7216_/A _7743_/X _7745_/X _7737_/X vssd1 vssd1 vccd1 vccd1 _8544_/D sky130_fd_sc_hd__o211a_1
X_4958_ _4909_/S _4947_/X _4957_/Y vssd1 vssd1 vccd1 vccd1 _8168_/D sky130_fd_sc_hd__a21oi_1
X_3909_ _3908_/X _8513_/Q _3912_/S vssd1 vssd1 vccd1 vccd1 _3910_/A sky130_fd_sc_hd__mux2_1
X_4889_ _4713_/X _8180_/Q _4712_/X _4888_/X vssd1 vssd1 vccd1 vccd1 _4889_/X sky130_fd_sc_hd__a211o_1
X_7677_ _8178_/Q _7737_/A vssd1 vssd1 vccd1 vccd1 _7678_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3409_ clkbuf_0__3409_/X vssd1 vssd1 vccd1 vccd1 _6889__385/A sky130_fd_sc_hd__clkbuf_4
XFILLER_117_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6559_ _6571_/A vssd1 vssd1 vccd1 vccd1 _6559_/X sky130_fd_sc_hd__buf_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7396__121 _7400__125/A vssd1 vssd1 vccd1 vccd1 _8378_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3308_ _6724_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3308_/X sky130_fd_sc_hd__clkbuf_16
X_8229_ _8229_/CLK _8229_/D vssd1 vssd1 vccd1 vccd1 _8229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6537__233 _6538__234/A vssd1 vssd1 vccd1 vccd1 _7911_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7405__128 _7405__128/A vssd1 vssd1 vccd1 vccd1 _8385_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6921__397 _6924__400/A vssd1 vssd1 vccd1 vccd1 _8119_/CLK sky130_fd_sc_hd__inv_2
X_5930_ _5930_/A _5932_/B vssd1 vssd1 vccd1 vccd1 _5931_/A sky130_fd_sc_hd__or2_4
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5861_ _4114_/X _7770_/Q _5869_/S vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__mux2_1
X_7056__499 _7057__500/A vssd1 vssd1 vccd1 vccd1 _8226_/CLK sky130_fd_sc_hd__inv_2
X_7600_ _7600_/A _7600_/B vssd1 vssd1 vccd1 vccd1 _8476_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5792_ _5792_/A vssd1 vssd1 vccd1 vccd1 _7844_/D sky130_fd_sc_hd__clkbuf_1
X_4812_ _8232_/Q _4811_/X _4806_/X _8216_/Q _4760_/S vssd1 vssd1 vccd1 vccd1 _4812_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7531_ _7532_/B _7532_/C _7201_/A vssd1 vssd1 vccd1 vccd1 _7531_/Y sky130_fd_sc_hd__a21oi_1
X_4743_ _4713_/X _8184_/Q _4947_/A _4742_/X vssd1 vssd1 vccd1 vccd1 _4743_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4674_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4674_/X sky130_fd_sc_hd__buf_2
X_6413_ _7862_/Q _6328_/A _6233_/X vssd1 vssd1 vccd1 vccd1 _6413_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6344_ _7247_/A _7747_/A _6336_/X _6343_/X vssd1 vssd1 vccd1 vccd1 _6344_/X sky130_fd_sc_hd__a31o_1
XFILLER_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6275_ _8334_/Q vssd1 vssd1 vccd1 vccd1 _7298_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5226_ _8453_/Q _8191_/Q _5312_/S vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__mux2_1
X_8014_ _8531_/CLK _8014_/D vssd1 vssd1 vccd1 vccd1 _8014_/Q sky130_fd_sc_hd__dfxtp_1
X_5157_ _8407_/Q _8391_/Q _8383_/Q _8415_/Q _5284_/S _5061_/X vssd1 vssd1 vccd1 vccd1
+ _5157_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_0__3024_ _6166_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3024_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3410_ clkbuf_0__3410_/X vssd1 vssd1 vccd1 vccd1 _6892__387/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ _4027_/X _8405_/Q _4112_/S vssd1 vssd1 vccd1 vccd1 _4109_/A sky130_fd_sc_hd__mux2_1
X_5088_ _5181_/A vssd1 vssd1 vccd1 vccd1 _5088_/X sky130_fd_sc_hd__clkbuf_4
X_4039_ _5805_/B _5464_/A vssd1 vssd1 vccd1 vccd1 _4055_/S sky130_fd_sc_hd__or2_2
Xclkbuf_1_0_0__3272_ clkbuf_0__3272_/X vssd1 vssd1 vccd1 vccd1 _6652_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7729_ _7729_/A _7729_/B _7729_/C vssd1 vssd1 vccd1 vccd1 _7730_/A sky130_fd_sc_hd__or3_1
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6313__213 _6315__215/A vssd1 vssd1 vccd1 vccd1 _7843_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4390_ _4390_/A vssd1 vssd1 vccd1 vccd1 _8280_/D sky130_fd_sc_hd__clkbuf_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6060_ _6056_/X _6058_/X _6059_/X _6044_/X vssd1 vssd1 vccd1 vccd1 _6060_/X sky130_fd_sc_hd__o211a_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5011_ _5011_/A vssd1 vssd1 vccd1 vccd1 _8144_/D sky130_fd_sc_hd__clkbuf_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6962_ _7089_/A vssd1 vssd1 vccd1 vccd1 _6962_/X sky130_fd_sc_hd__buf_1
X_5913_ _7642_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__or2_1
X_5844_ _5844_/A vssd1 vssd1 vccd1 vccd1 _7778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3642_ _7414_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3642_/X sky130_fd_sc_hd__clkbuf_16
X_5775_ _5608_/X _7851_/Q _5779_/S vssd1 vssd1 vccd1 vccd1 _5776_/A sky130_fd_sc_hd__mux2_1
X_7514_ _7514_/A _7514_/B vssd1 vssd1 vccd1 vccd1 _7524_/C sky130_fd_sc_hd__nor2_1
X_4726_ _4726_/A vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__clkbuf_2
X_8494_ _8530_/CLK _8494_/D vssd1 vssd1 vccd1 vccd1 _8494_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7445_ _7457_/A vssd1 vssd1 vccd1 vccd1 _7445_/X sky130_fd_sc_hd__buf_1
X_4657_ _8142_/Q _8029_/Q _7925_/Q _7909_/Q _4655_/X _4656_/X vssd1 vssd1 vccd1 vccd1
+ _4657_/X sky130_fd_sc_hd__mux4_1
Xinput80 wbs_data_i[19] vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__buf_4
Xinput91 wbs_data_i[29] vssd1 vssd1 vccd1 vccd1 _5965_/A sky130_fd_sc_hd__buf_4
X_7376_ _8128_/Q _7679_/B _7366_/X _7375_/X _7371_/X vssd1 vssd1 vccd1 vccd1 _8365_/D
+ sky130_fd_sc_hd__o311a_1
X_6327_ _6521_/A vssd1 vssd1 vccd1 vccd1 _6328_/A sky130_fd_sc_hd__buf_2
X_4588_ _4418_/X _8204_/Q _4596_/S vssd1 vssd1 vccd1 vccd1 _4589_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6258_ _7640_/A _7815_/Q _6258_/S vssd1 vssd1 vccd1 vccd1 _6259_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5209_ _8446_/Q _5063_/B _5208_/X _5244_/A vssd1 vssd1 vccd1 vccd1 _5209_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6189_ _7819_/Q _7820_/Q vssd1 vssd1 vccd1 vccd1 _6210_/A sky130_fd_sc_hd__or2b_1
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6720__322 _6720__322/A vssd1 vssd1 vccd1 vccd1 _8032_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3255_ clkbuf_0__3255_/X vssd1 vssd1 vccd1 vccd1 _6588__275/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6953__419 _6954__420/A vssd1 vssd1 vccd1 vccd1 _8143_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3890_ _3912_/S vssd1 vssd1 vccd1 vccd1 _3903_/S sky130_fd_sc_hd__buf_2
XFILLER_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _5559_/X _7996_/Q _5567_/S vssd1 vssd1 vccd1 vccd1 _5561_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5491_ _5491_/A vssd1 vssd1 vccd1 vccd1 _8050_/D sky130_fd_sc_hd__clkbuf_1
X_4511_ _5641_/A _4959_/A vssd1 vssd1 vccd1 vccd1 _4529_/S sky130_fd_sc_hd__nor2_2
XFILLER_8_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4442_ _4441_/X _8262_/Q _4445_/S vssd1 vssd1 vccd1 vccd1 _4443_/A sky130_fd_sc_hd__mux2_1
X_7230_ _8546_/Q _7319_/A _7319_/B vssd1 vssd1 vccd1 vccd1 _7281_/B sky130_fd_sc_hd__nand3b_1
X_4373_ _4373_/A vssd1 vssd1 vccd1 vccd1 _8285_/D sky130_fd_sc_hd__clkbuf_1
X_6112_ _7797_/Q _6122_/A vssd1 vssd1 vccd1 vccd1 _6112_/X sky130_fd_sc_hd__or2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6043_ _6082_/A vssd1 vssd1 vccd1 vccd1 _6063_/A sky130_fd_sc_hd__buf_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7994_ _7994_/CLK _7994_/D vssd1 vssd1 vccd1 vccd1 _7994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3657_ clkbuf_0__3657_/X vssd1 vssd1 vccd1 vccd1 _7670_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6893__388 _6895__390/A vssd1 vssd1 vccd1 vccd1 _8102_/CLK sky130_fd_sc_hd__inv_2
X_5827_ _7828_/Q _5559_/A _5833_/S vssd1 vssd1 vccd1 vccd1 _5828_/A sky130_fd_sc_hd__mux2_1
X_7112__544 _7113__545/A vssd1 vssd1 vccd1 vccd1 _8271_/CLK sky130_fd_sc_hd__inv_2
X_8546_ _8550_/CLK _8546_/D vssd1 vssd1 vccd1 vccd1 _8546_/Q sky130_fd_sc_hd__dfxtp_2
X_5758_ _5758_/A vssd1 vssd1 vccd1 vccd1 _7907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4709_ _4638_/X _4696_/X _4700_/X _4708_/X vssd1 vssd1 vccd1 vccd1 _4709_/X sky130_fd_sc_hd__a31o_1
X_8477_ _8479_/CLK _8477_/D vssd1 vssd1 vccd1 vccd1 _8477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5689_ _7937_/Q _5590_/X _5689_/S vssd1 vssd1 vccd1 vccd1 _5690_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7359_ _7359_/A _7359_/B vssd1 vssd1 vccd1 vccd1 _7360_/C sky130_fd_sc_hd__nand2_1
XFILLER_89_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7492__24 _7493__25/A vssd1 vssd1 vccd1 vccd1 _8456_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3307_ clkbuf_0__3307_/X vssd1 vssd1 vccd1 vccd1 _6720__322/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7013__464 _7014__465/A vssd1 vssd1 vccd1 vccd1 _8191_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _4991_/A vssd1 vssd1 vccd1 vccd1 _8153_/D sky130_fd_sc_hd__clkbuf_1
X_3942_ _3896_/X _8501_/Q _3946_/S vssd1 vssd1 vccd1 vccd1 _3943_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6661_ _6661_/A vssd1 vssd1 vccd1 vccd1 _8000_/D sky130_fd_sc_hd__clkbuf_1
X_3873_ _7637_/A _6326_/A _6035_/A vssd1 vssd1 vccd1 vccd1 _3873_/X sky130_fd_sc_hd__and3_1
X_8400_ _8400_/CLK _8400_/D vssd1 vssd1 vccd1 vccd1 _8400_/Q sky130_fd_sc_hd__dfxtp_1
X_5612_ _5611_/X _7978_/Q _5614_/S vssd1 vssd1 vccd1 vccd1 _5613_/A sky130_fd_sc_hd__mux2_1
X_8331_ _8331_/CLK _8331_/D vssd1 vssd1 vccd1 vccd1 _8331_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3410_ _6890_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3410_/X sky130_fd_sc_hd__clkbuf_16
X_5543_ _5543_/A vssd1 vssd1 vccd1 vccd1 _8027_/D sky130_fd_sc_hd__clkbuf_1
X_6179__186 _6180__187/A vssd1 vssd1 vccd1 vccd1 _7773_/CLK sky130_fd_sc_hd__inv_2
X_5474_ _3972_/X _8057_/Q _5474_/S vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__mux2_1
X_8262_ _8262_/CLK _8262_/D vssd1 vssd1 vccd1 vccd1 _8262_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3272_ _6639_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3272_/X sky130_fd_sc_hd__clkbuf_16
X_4425_ _4424_/X _8267_/Q _4436_/S vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__mux2_1
X_8193_ _8193_/CLK _8193_/D vssd1 vssd1 vccd1 vccd1 _8193_/Q sky130_fd_sc_hd__dfxtp_1
X_7213_ _7213_/A vssd1 vssd1 vccd1 vccd1 _7232_/B sky130_fd_sc_hd__clkbuf_2
X_4356_ _5805_/A _4356_/B vssd1 vssd1 vccd1 vccd1 _4372_/S sky130_fd_sc_hd__or2_2
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _4286_/X _8321_/Q _4290_/S vssd1 vssd1 vccd1 vccd1 _4288_/A sky130_fd_sc_hd__mux2_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7390__116 _7392__118/A vssd1 vssd1 vccd1 vccd1 _8373_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _8015_/Q _6030_/B vssd1 vssd1 vccd1 vccd1 _6027_/A sky130_fd_sc_hd__and2_2
X_8600__247 vssd1 vssd1 vccd1 vccd1 _8600__247/HI versionID[1] sky130_fd_sc_hd__conb_1
XFILLER_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7977_ _7977_/CLK _7977_/D vssd1 vssd1 vccd1 vccd1 _7977_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3023_ clkbuf_0__3023_/X vssd1 vssd1 vccd1 vccd1 _6291_/A sky130_fd_sc_hd__clkbuf_4
X_6859_ _7201_/A _7598_/A vssd1 vssd1 vccd1 vccd1 _6860_/D sky130_fd_sc_hd__xor2_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8529_ _8530_/CLK _8529_/D vssd1 vssd1 vccd1 vccd1 _8529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6531__228 _6533__230/A vssd1 vssd1 vccd1 vccd1 _7906_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_60 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_71 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_93 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_82 _5973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6733__332 _6733__332/A vssd1 vssd1 vccd1 vccd1 _8042_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7138__64 _7139__65/A vssd1 vssd1 vccd1 vccd1 _8291_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4210_ _4210_/A vssd1 vssd1 vccd1 vccd1 _8382_/D sky130_fd_sc_hd__clkbuf_1
X_7061__502 _7063__504/A vssd1 vssd1 vccd1 vccd1 _8229_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5190_ _8507_/Q _5207_/A vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__or2_1
XFILLER_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4141_ _4141_/A _4141_/B vssd1 vssd1 vccd1 vccd1 _4141_/X sky130_fd_sc_hd__and2_1
X_4072_ _4031_/X _8420_/Q _4074_/S vssd1 vssd1 vccd1 vccd1 _4073_/A sky130_fd_sc_hd__mux2_1
X_6586__273 _6588__275/A vssd1 vssd1 vccd1 vccd1 _7951_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7454__168 _7456__170/A vssd1 vssd1 vccd1 vccd1 _8425_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7900_ _8551_/CLK _7900_/D vssd1 vssd1 vccd1 vccd1 _7900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7831_ _7831_/CLK _7831_/D vssd1 vssd1 vccd1 vccd1 _7831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4974_ _4974_/A vssd1 vssd1 vccd1 vccd1 _8160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7762_ _8550_/CLK _7762_/D vssd1 vssd1 vccd1 vccd1 _7762_/Q sky130_fd_sc_hd__dfxtp_1
X_7693_ _7693_/A vssd1 vssd1 vccd1 vccd1 _8529_/D sky130_fd_sc_hd__clkbuf_1
X_3925_ _3899_/X _8508_/Q _3927_/S vssd1 vssd1 vccd1 vccd1 _3926_/A sky130_fd_sc_hd__mux2_1
X_3856_ _3853_/Y _3855_/X _3849_/B vssd1 vssd1 vccd1 vccd1 _3860_/C sky130_fd_sc_hd__a21oi_1
XFILLER_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5526_ _5399_/X _8034_/Q _5528_/S vssd1 vssd1 vccd1 vccd1 _5527_/A sky130_fd_sc_hd__mux2_1
X_8314_ _8314_/CLK _8314_/D vssd1 vssd1 vccd1 vccd1 _8314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5457_ _5457_/A vssd1 vssd1 vccd1 vccd1 _8068_/D sky130_fd_sc_hd__clkbuf_1
X_8245_ _8245_/CLK _8245_/D vssd1 vssd1 vccd1 vccd1 _8245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4408_ _4385_/X _8273_/Q _4410_/S vssd1 vssd1 vccd1 vccd1 _4409_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3641_ clkbuf_0__3641_/X vssd1 vssd1 vccd1 vccd1 _7411__133/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3255_ _6583_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3255_/X sky130_fd_sc_hd__clkbuf_16
X_5388_ _5387_/X _8098_/Q _5388_/S vssd1 vssd1 vccd1 vccd1 _5389_/A sky130_fd_sc_hd__mux2_1
X_8176_ _8176_/CLK _8176_/D vssd1 vssd1 vccd1 vccd1 _8176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4339_ _4354_/S vssd1 vssd1 vccd1 vccd1 _4348_/S sky130_fd_sc_hd__buf_2
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7058_ _7058_/A vssd1 vssd1 vccd1 vccd1 _7058_/X sky130_fd_sc_hd__buf_1
X_6009_ _6009_/A vssd1 vssd1 vccd1 vccd1 _6009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4690_ _6900_/B vssd1 vssd1 vccd1 vccd1 _4690_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6360_ _6331_/X _6344_/X _6359_/X _6233_/X vssd1 vssd1 vccd1 vccd1 _6360_/X sky130_fd_sc_hd__a31o_1
XFILLER_115_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5311_ _5306_/X _5307_/X _5206_/A _5310_/X vssd1 vssd1 vccd1 vccd1 _5311_/X sky130_fd_sc_hd__a211o_1
XFILLER_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6291_ _6291_/A vssd1 vssd1 vccd1 vccd1 _6291_/X sky130_fd_sc_hd__buf_1
X_8030_ _8030_/CLK _8030_/D vssd1 vssd1 vccd1 vccd1 _8030_/Q sky130_fd_sc_hd__dfxtp_1
X_5242_ _8421_/Q _5239_/X _5101_/S _5241_/X vssd1 vssd1 vccd1 vccd1 _5243_/C sky130_fd_sc_hd__o211a_1
X_5173_ _5047_/X _5160_/X _5164_/X _5172_/X vssd1 vssd1 vccd1 vccd1 _5173_/X sky130_fd_sc_hd__a31o_2
XFILLER_68_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4124_ _4217_/A _8169_/Q vssd1 vssd1 vccd1 vccd1 _4125_/A sky130_fd_sc_hd__xor2_1
XFILLER_29_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput1 caravel_uart_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4055_ _4035_/X _8427_/Q _4055_/S vssd1 vssd1 vccd1 vccd1 _4056_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6779__365 _6779__365/A vssd1 vssd1 vccd1 vccd1 _8078_/CLK sky130_fd_sc_hd__inv_2
X_7814_ _8355_/CLK _7814_/D vssd1 vssd1 vccd1 vccd1 _7814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6972__433 _6973__434/A vssd1 vssd1 vccd1 vccd1 _8157_/CLK sky130_fd_sc_hd__inv_2
X_7745_ _7646_/A _7731_/X _7744_/X vssd1 vssd1 vccd1 vccd1 _7745_/X sky130_fd_sc_hd__a21bo_1
X_4957_ _4909_/S _4955_/A _6900_/B vssd1 vssd1 vccd1 vccd1 _4957_/Y sky130_fd_sc_hd__o21ai_1
X_6933__406 _6936__409/A vssd1 vssd1 vccd1 vccd1 _8128_/CLK sky130_fd_sc_hd__inv_2
X_4888_ _4872_/X _4887_/X _4948_/A vssd1 vssd1 vccd1 vccd1 _4888_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7676_ _7680_/A _7676_/B vssd1 vssd1 vccd1 vccd1 _8520_/D sky130_fd_sc_hd__nor2_1
X_3908_ _8489_/Q vssd1 vssd1 vccd1 vccd1 _3908_/X sky130_fd_sc_hd__buf_4
Xclkbuf_1_1_0__3408_ clkbuf_0__3408_/X vssd1 vssd1 vccd1 vccd1 _6881__378/A sky130_fd_sc_hd__clkbuf_4
X_7068__508 _7069__509/A vssd1 vssd1 vccd1 vccd1 _8235_/CLK sky130_fd_sc_hd__inv_2
X_3839_ _8120_/Q vssd1 vssd1 vccd1 vccd1 _3956_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6558_ _6589_/A vssd1 vssd1 vccd1 vccd1 _6558_/X sky130_fd_sc_hd__buf_1
XFILLER_4_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8565__212 vssd1 vssd1 vccd1 vccd1 _8565__212/HI caravel_irq[3] sky130_fd_sc_hd__conb_1
XFILLER_105_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5509_ _5509_/A vssd1 vssd1 vccd1 vccd1 _8042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6489_ _6511_/A vssd1 vssd1 vccd1 vccd1 _6498_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3307_ _6718_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3307_/X sky130_fd_sc_hd__clkbuf_16
X_7132__59 _7133__60/A vssd1 vssd1 vccd1 vccd1 _8286_/CLK sky130_fd_sc_hd__inv_2
X_8228_ _8228_/CLK _8228_/D vssd1 vssd1 vccd1 vccd1 _8228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8159_ _8159_/CLK _8159_/D vssd1 vssd1 vccd1 vccd1 _8159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7674__49 _7675__50/A vssd1 vssd1 vccd1 vccd1 _8518_/CLK sky130_fd_sc_hd__inv_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5860_ _5875_/S vssd1 vssd1 vccd1 vccd1 _5869_/S sky130_fd_sc_hd__buf_2
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _4811_/A vssd1 vssd1 vccd1 vccd1 _4811_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5791_ _7844_/Q _4280_/A _5797_/S vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4742_ _4638_/X _4721_/X _4725_/X _4741_/X vssd1 vssd1 vccd1 vccd1 _4742_/X sky130_fd_sc_hd__a31o_1
X_7530_ _7598_/A _7530_/B _7530_/C _7530_/D vssd1 vssd1 vccd1 vccd1 _7535_/C sky130_fd_sc_hd__and4_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4673_ _4740_/A vssd1 vssd1 vccd1 vccd1 _4673_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6412_ _6397_/X _6408_/X _6410_/X _6437_/A vssd1 vssd1 vccd1 vccd1 _6412_/X sky130_fd_sc_hd__a22o_1
X_6343_ _6397_/A vssd1 vssd1 vccd1 vccd1 _6343_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6274_ _6274_/A vssd1 vssd1 vccd1 vccd1 _7820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8013_ _8531_/CLK _8013_/D vssd1 vssd1 vccd1 vccd1 _8013_/Q sky130_fd_sc_hd__dfxtp_1
X_5225_ _3902_/X _5038_/X _5224_/X _5111_/X vssd1 vssd1 vccd1 vccd1 _8128_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_0__3023_ _6165_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3023_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_102_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5156_ _3896_/X _5038_/X _5155_/X _5111_/X vssd1 vssd1 vccd1 vccd1 _8130_/D sky130_fd_sc_hd__o211a_1
X_4107_ _4107_/A vssd1 vssd1 vccd1 vccd1 _8406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5087_ _5215_/S vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3271_ clkbuf_0__3271_/X vssd1 vssd1 vccd1 vccd1 _6925_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4038_ _4038_/A _5345_/B _5109_/A _3956_/B vssd1 vssd1 vccd1 vccd1 _5464_/A sky130_fd_sc_hd__or4bb_4
XFILLER_25_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5989_ _5989_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5990_/A sky130_fd_sc_hd__and2_1
X_6599__283 _6601__285/A vssd1 vssd1 vccd1 vccd1 _7961_/CLK sky130_fd_sc_hd__inv_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7728_ _7728_/A _7731_/A _7728_/C vssd1 vssd1 vccd1 vccd1 _7729_/C sky130_fd_sc_hd__and3_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput190 _6127_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_87_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6979__439 _6979__439/A vssd1 vssd1 vccd1 vccd1 _8163_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3469_ clkbuf_0__3469_/X vssd1 vssd1 vccd1 vccd1 _7149__73/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7411__133 _7411__133/A vssd1 vssd1 vccd1 vccd1 _8390_/CLK sky130_fd_sc_hd__inv_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5010_ _8144_/Q _4484_/X _5012_/S vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__mux2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6961_ _6961_/A vssd1 vssd1 vccd1 vccd1 _6961_/X sky130_fd_sc_hd__buf_1
X_5912_ _5969_/B vssd1 vssd1 vccd1 vccd1 _5921_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5843_ _4114_/X _7778_/Q _5851_/S vssd1 vssd1 vccd1 vccd1 _5844_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3641_ _7408_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3641_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5774_ _5774_/A vssd1 vssd1 vccd1 vccd1 _7852_/D sky130_fd_sc_hd__clkbuf_1
X_7513_ _7513_/A _7513_/B _7513_/C _7513_/D vssd1 vssd1 vccd1 vccd1 _7524_/B sky130_fd_sc_hd__or4_1
X_4725_ _4953_/B _4722_/X _4724_/X vssd1 vssd1 vccd1 vccd1 _4725_/X sky130_fd_sc_hd__a21o_1
X_8493_ _8527_/CLK _8493_/D vssd1 vssd1 vccd1 vccd1 _8493_/Q sky130_fd_sc_hd__dfxtp_2
X_4656_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4656_/X sky130_fd_sc_hd__buf_2
X_4587_ _4602_/S vssd1 vssd1 vccd1 vccd1 _4596_/S sky130_fd_sc_hd__buf_2
Xinput70 wbs_data_i[0] vssd1 vssd1 vccd1 vccd1 _7631_/A sky130_fd_sc_hd__buf_8
Xinput81 wbs_data_i[1] vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__clkbuf_2
X_7375_ _8365_/Q _7377_/B vssd1 vssd1 vccd1 vccd1 _7375_/X sky130_fd_sc_hd__or2_1
Xinput92 wbs_data_i[2] vssd1 vssd1 vccd1 vccd1 _7635_/A sky130_fd_sc_hd__buf_8
X_6326_ _6326_/A vssd1 vssd1 vccd1 vccd1 _6521_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6257_ _6257_/A vssd1 vssd1 vccd1 vccd1 _7814_/D sky130_fd_sc_hd__clkbuf_1
X_5208_ _7833_/Q _8430_/Q _5318_/S vssd1 vssd1 vccd1 vccd1 _5208_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6188_ _6367_/A vssd1 vssd1 vccd1 vccd1 _6188_/X sky130_fd_sc_hd__buf_4
X_5139_ _5354_/B _5138_/X _5083_/X vssd1 vssd1 vccd1 vccd1 _5139_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3254_ clkbuf_0__3254_/X vssd1 vssd1 vccd1 vccd1 _6579__267/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6580__268 _6582__270/A vssd1 vssd1 vccd1 vccd1 _7946_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5490_ _8050_/Q _4286_/A _5492_/S vssd1 vssd1 vccd1 vccd1 _5491_/A sky130_fd_sc_hd__mux2_1
X_4510_ _4466_/B _5014_/C _5014_/A vssd1 vssd1 vccd1 vccd1 _4959_/A sky130_fd_sc_hd__nand3b_2
X_4441_ _8107_/Q vssd1 vssd1 vccd1 vccd1 _4441_/X sky130_fd_sc_hd__buf_2
XFILLER_8_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4372_ _4298_/X _8285_/Q _4372_/S vssd1 vssd1 vccd1 vccd1 _4373_/A sky130_fd_sc_hd__mux2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _7872_/Q input12/X _6111_/S vssd1 vssd1 vccd1 vccd1 _6111_/X sky130_fd_sc_hd__mux2_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6042_ _7779_/Q _7633_/A vssd1 vssd1 vccd1 vccd1 _6042_/X sky130_fd_sc_hd__or2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7418__139 _7419__140/A vssd1 vssd1 vccd1 vccd1 _8396_/CLK sky130_fd_sc_hd__inv_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7993_ _7993_/CLK _7993_/D vssd1 vssd1 vccd1 vccd1 _7993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3656_ clkbuf_0__3656_/X vssd1 vssd1 vccd1 vccd1 _7490__22/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5826_ _5826_/A vssd1 vssd1 vccd1 vccd1 _7829_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8545_ _8550_/CLK _8545_/D vssd1 vssd1 vccd1 vccd1 _8545_/Q sky130_fd_sc_hd__dfxtp_4
X_5757_ _7907_/Q _5396_/A _5761_/S vssd1 vssd1 vccd1 vccd1 _5758_/A sky130_fd_sc_hd__mux2_1
X_4708_ _4673_/X _4703_/X _4707_/X _4684_/X vssd1 vssd1 vccd1 vccd1 _4708_/X sky130_fd_sc_hd__o211a_1
X_8476_ _8479_/CLK _8476_/D vssd1 vssd1 vccd1 vccd1 _8476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5688_ _5688_/A vssd1 vssd1 vccd1 vccd1 _7938_/D sky130_fd_sc_hd__clkbuf_1
X_7477__11 _7479__13/A vssd1 vssd1 vccd1 vccd1 _8443_/CLK sky130_fd_sc_hd__inv_2
X_4639_ _4651_/A vssd1 vssd1 vccd1 vccd1 _4658_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7358_ _8360_/Q _7354_/Y _7357_/X _7286_/X vssd1 vssd1 vccd1 vccd1 _8360_/D sky130_fd_sc_hd__o211a_1
XFILLER_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3306_ clkbuf_0__3306_/X vssd1 vssd1 vccd1 vccd1 _6716__319/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3321_ clkbuf_0__3321_/X vssd1 vssd1 vccd1 vccd1 _6870__370/A sky130_fd_sc_hd__clkbuf_16
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7185__101 _7186__102/A vssd1 vssd1 vccd1 vccd1 _8328_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _8153_/Q _4481_/X _4994_/S vssd1 vssd1 vccd1 vccd1 _4991_/A sky130_fd_sc_hd__mux2_1
X_3941_ _3941_/A vssd1 vssd1 vccd1 vccd1 _8502_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3441_ clkbuf_0__3441_/X vssd1 vssd1 vccd1 vccd1 _7014__465/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3872_ _6108_/A _6082_/A vssd1 vssd1 vccd1 vccd1 _6035_/A sky130_fd_sc_hd__and2_2
X_6660_ _5924_/A _8000_/Q _6664_/S vssd1 vssd1 vccd1 vccd1 _6661_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5611_ _8110_/Q vssd1 vssd1 vccd1 vccd1 _5611_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8330_ _8330_/CLK _8330_/D vssd1 vssd1 vccd1 vccd1 _8330_/Q sky130_fd_sc_hd__dfxtp_1
X_5542_ _5396_/X _8027_/Q _5546_/S vssd1 vssd1 vccd1 vccd1 _5543_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5473_ _5473_/A vssd1 vssd1 vccd1 vccd1 _8058_/D sky130_fd_sc_hd__clkbuf_1
X_8261_ _8261_/CLK _8261_/D vssd1 vssd1 vccd1 vccd1 _8261_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3271_ _6638_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3271_/X sky130_fd_sc_hd__clkbuf_16
X_8192_ _8192_/CLK _8192_/D vssd1 vssd1 vccd1 vccd1 _8192_/Q sky130_fd_sc_hd__dfxtp_1
X_7212_ _8347_/Q vssd1 vssd1 vccd1 vccd1 _7236_/A sky130_fd_sc_hd__clkbuf_2
X_4424_ _8112_/Q vssd1 vssd1 vccd1 vccd1 _4424_/X sky130_fd_sc_hd__clkbuf_4
X_4355_ _4355_/A vssd1 vssd1 vccd1 vccd1 _8293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _4286_/A vssd1 vssd1 vccd1 vccd1 _4286_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6025_/A vssd1 vssd1 vccd1 vccd1 _6025_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7976_ _7976_/CLK _7976_/D vssd1 vssd1 vccd1 vccd1 _7976_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0__3639_ clkbuf_0__3639_/X vssd1 vssd1 vccd1 vccd1 _7420_/A sky130_fd_sc_hd__clkbuf_4
X_6858_ _8476_/Q _7532_/C _6857_/X vssd1 vssd1 vccd1 vccd1 _7598_/A sky130_fd_sc_hd__a21oi_2
X_5809_ _3963_/X _7836_/Q _5815_/S vssd1 vssd1 vccd1 vccd1 _5810_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6789_ _8464_/Q _8463_/Q _8462_/Q _8461_/Q vssd1 vssd1 vccd1 vccd1 _6818_/A sky130_fd_sc_hd__and4_1
X_8528_ _8530_/CLK _8528_/D vssd1 vssd1 vccd1 vccd1 _8528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8459_ _8479_/CLK _8459_/D vssd1 vssd1 vccd1 vccd1 _8459_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3469_ _7146_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3469_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7170__90 _7170__90/A vssd1 vssd1 vccd1 vccd1 _8317_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_50 _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_61 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_94 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_83 _5973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_72 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8582__229 vssd1 vssd1 vccd1 vccd1 _8582__229/HI manufacturerID[1] sky130_fd_sc_hd__conb_1
X_4140_ _4622_/A _4931_/A _4622_/B _4622_/C vssd1 vssd1 vccd1 vccd1 _4141_/B sky130_fd_sc_hd__a211o_1
XFILLER_95_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4071_ _4071_/A vssd1 vssd1 vccd1 vccd1 _8421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7830_ _7830_/CLK _7830_/D vssd1 vssd1 vccd1 vccd1 _7830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _8160_/Q _4484_/X _4975_/S vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__mux2_1
X_7761_ _7247_/A _7747_/Y _7760_/X vssd1 vssd1 vccd1 vccd1 _8551_/D sky130_fd_sc_hd__a21o_1
X_6185__191 _6185__191/A vssd1 vssd1 vccd1 vccd1 _7778_/CLK sky130_fd_sc_hd__inv_2
X_6712_ _6718_/A vssd1 vssd1 vccd1 vccd1 _6712_/X sky130_fd_sc_hd__buf_1
X_3924_ _3924_/A vssd1 vssd1 vccd1 vccd1 _8509_/D sky130_fd_sc_hd__clkbuf_1
X_7692_ _7719_/A _8523_/Q vssd1 vssd1 vccd1 vccd1 _7693_/A sky130_fd_sc_hd__and2_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3424_ clkbuf_0__3424_/X vssd1 vssd1 vccd1 vccd1 _6936__409/A sky130_fd_sc_hd__clkbuf_4
X_3855_ _8120_/Q _8119_/Q _5034_/A vssd1 vssd1 vccd1 vccd1 _3855_/X sky130_fd_sc_hd__a21o_1
X_6593__278 _6594__279/A vssd1 vssd1 vccd1 vccd1 _7956_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5525_ _5525_/A vssd1 vssd1 vccd1 vccd1 _8035_/D sky130_fd_sc_hd__clkbuf_1
X_8313_ _8313_/CLK _8313_/D vssd1 vssd1 vccd1 vccd1 _8313_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_opt_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8355_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5456_ _8068_/Q _4187_/X _5456_/S vssd1 vssd1 vccd1 vccd1 _5457_/A sky130_fd_sc_hd__mux2_1
X_6634__297 _6635__298/A vssd1 vssd1 vccd1 vccd1 _7983_/CLK sky130_fd_sc_hd__inv_2
X_8244_ _8244_/CLK _8244_/D vssd1 vssd1 vccd1 vccd1 _8244_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3254_ _6577_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3254_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3640_ clkbuf_0__3640_/X vssd1 vssd1 vccd1 vccd1 _7407__130/A sky130_fd_sc_hd__clkbuf_4
X_4407_ _4407_/A vssd1 vssd1 vccd1 vccd1 _8274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5387_ _5575_/A vssd1 vssd1 vccd1 vccd1 _5387_/X sky130_fd_sc_hd__clkbuf_2
X_8175_ _8175_/CLK _8175_/D vssd1 vssd1 vccd1 vccd1 _8175_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4338_ _5482_/A _4356_/B vssd1 vssd1 vccd1 vccd1 _4354_/S sky130_fd_sc_hd__or2_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4269_ _8327_/Q _4190_/X _4273_/S vssd1 vssd1 vccd1 vccd1 _4270_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6008_ _8007_/Q _6008_/B vssd1 vssd1 vccd1 vccd1 _6009_/A sky130_fd_sc_hd__and2_1
XFILLER_101_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7959_ _7959_/CLK _7959_/D vssd1 vssd1 vccd1 vccd1 _7959_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5310_ _5306_/A _5308_/X _5309_/X _5250_/X vssd1 vssd1 vccd1 vccd1 _5310_/X sky130_fd_sc_hd__o211a_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7460__173 _7460__173/A vssd1 vssd1 vccd1 vccd1 _8430_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5241_ _8271_/Q _5063_/B _5240_/X _5230_/A vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5172_ _5293_/A _5167_/X _5169_/X _5171_/X _5177_/A vssd1 vssd1 vccd1 vccd1 _5172_/X
+ sky130_fd_sc_hd__o221a_1
X_7026__475 _7026__475/A vssd1 vssd1 vccd1 vccd1 _8202_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4123_ _7635_/A _6035_/A _4122_/Y _6247_/A vssd1 vssd1 vccd1 vccd1 _6902_/A sky130_fd_sc_hd__a31oi_4
Xinput2 caravel_wb_ack_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4054_ _4054_/A vssd1 vssd1 vccd1 vccd1 _8428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7813_ _8355_/CLK _7813_/D vssd1 vssd1 vccd1 vccd1 _7813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7744_ _7754_/B vssd1 vssd1 vccd1 vccd1 _7744_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4956_ _4716_/X _4947_/X _4955_/Y _4924_/X vssd1 vssd1 vccd1 vccd1 _8169_/D sky130_fd_sc_hd__o211a_1
X_6601__285 _6601__285/A vssd1 vssd1 vccd1 vccd1 _7963_/CLK sky130_fd_sc_hd__inv_2
X_3907_ _3907_/A vssd1 vssd1 vccd1 vccd1 _8514_/D sky130_fd_sc_hd__clkbuf_1
X_4887_ _4740_/X _4875_/X _4879_/X _4886_/X _4638_/A vssd1 vssd1 vccd1 vccd1 _4887_/X
+ sky130_fd_sc_hd__o311a_1
X_6626_ _6626_/A vssd1 vssd1 vccd1 vccd1 _6626_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3407_ clkbuf_0__3407_/X vssd1 vssd1 vccd1 vccd1 _6890_/A sky130_fd_sc_hd__clkbuf_4
X_3838_ _4256_/C _5334_/A _4256_/A vssd1 vssd1 vccd1 vccd1 _5500_/A sky130_fd_sc_hd__nand3b_4
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3269_ clkbuf_0__3269_/X vssd1 vssd1 vccd1 vccd1 _6631__295/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5508_ _8042_/Q _4286_/A _5510_/S vssd1 vssd1 vccd1 vccd1 _5509_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6488_ _6488_/A vssd1 vssd1 vccd1 vccd1 _7886_/D sky130_fd_sc_hd__clkbuf_1
X_5439_ _5439_/A vssd1 vssd1 vccd1 vccd1 _8076_/D sky130_fd_sc_hd__clkbuf_1
X_8227_ _8227_/CLK _8227_/D vssd1 vssd1 vccd1 vccd1 _8227_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3306_ _6712_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3306_/X sky130_fd_sc_hd__clkbuf_16
X_8158_ _8158_/CLK _8158_/D vssd1 vssd1 vccd1 vccd1 _8158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8089_ _8089_/CLK _8089_/D vssd1 vssd1 vccd1 vccd1 _8089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7659__36 _7660__37/A vssd1 vssd1 vccd1 vccd1 _8505_/CLK sky130_fd_sc_hd__inv_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6544__239 _6544__239/A vssd1 vssd1 vccd1 vccd1 _7917_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _8162_/Q _8200_/Q _4810_/S vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5790_ _5790_/A vssd1 vssd1 vccd1 vccd1 _7845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4731_/X _4735_/X _4739_/X _4740_/X _4684_/X vssd1 vssd1 vccd1 vccd1 _4741_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4672_ _4664_/X _4665_/X _4671_/X vssd1 vssd1 vccd1 vccd1 _4672_/X sky130_fd_sc_hd__a21o_1
X_8588__235 vssd1 vssd1 vccd1 vccd1 _8588__235/HI manufacturerID[7] sky130_fd_sc_hd__conb_1
X_6411_ _6411_/A vssd1 vssd1 vccd1 vccd1 _6437_/A sky130_fd_sc_hd__buf_2
XFILLER_115_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6342_ _7742_/C _6398_/B vssd1 vssd1 vccd1 vccd1 _6397_/A sky130_fd_sc_hd__or2_1
XFILLER_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6273_ _6272_/X _6273_/B vssd1 vssd1 vccd1 vccd1 _6274_/A sky130_fd_sc_hd__and2b_1
XFILLER_103_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8012_ _8531_/CLK _8012_/D vssd1 vssd1 vccd1 vccd1 _8012_/Q sky130_fd_sc_hd__dfxtp_4
X_5224_ _8128_/Q _5040_/X _5349_/A _5223_/X _5107_/X vssd1 vssd1 vccd1 vccd1 _5224_/X
+ sky130_fd_sc_hd__a221o_1
X_6746__343 _6746__343/A vssd1 vssd1 vccd1 vccd1 _8053_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3022_ _6164_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3022_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5155_ _8130_/Q _5040_/X _5348_/A _5154_/X _5107_/X vssd1 vssd1 vccd1 vccd1 _5155_/X
+ sky130_fd_sc_hd__a221o_1
X_4106_ _4023_/X _8406_/Q _4106_/S vssd1 vssd1 vccd1 vccd1 _4107_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5086_ _5250_/A vssd1 vssd1 vccd1 vccd1 _5169_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4037_ _4037_/A vssd1 vssd1 vccd1 vccd1 _8435_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3270_ clkbuf_0__3270_/X vssd1 vssd1 vccd1 vccd1 _6635__298/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7074__513 _7076__515/A vssd1 vssd1 vccd1 vccd1 _8240_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5988_ _6010_/A vssd1 vssd1 vccd1 vccd1 _5997_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7727_ _7728_/C _7727_/B vssd1 vssd1 vccd1 vccd1 _7729_/B sky130_fd_sc_hd__and2b_1
X_4939_ _5014_/C _4943_/A vssd1 vssd1 vccd1 vccd1 _4939_/X sky130_fd_sc_hd__or2_1
X_7658_ _7664_/A vssd1 vssd1 vccd1 vccd1 _7658_/X sky130_fd_sc_hd__buf_1
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6609_ _8180_/Q _8167_/D vssd1 vssd1 vccd1 vccd1 _6610_/A sky130_fd_sc_hd__and2_1
XFILLER_4_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7589_ _7587_/Y _7588_/X _7575_/X _6800_/B vssd1 vssd1 vccd1 vccd1 _7590_/B sky130_fd_sc_hd__o22a_1
Xclkbuf_opt_1_0_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _7120_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_106_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput180 _6091_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[12] sky130_fd_sc_hd__buf_2
Xoutput191 _6130_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[22] sky130_fd_sc_hd__buf_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3468_ clkbuf_0__3468_/X vssd1 vssd1 vccd1 vccd1 _7145__70/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6320__219 _6321__220/A vssd1 vssd1 vccd1 vccd1 _7849_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5911_ _5911_/A vssd1 vssd1 vccd1 vccd1 _5911_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5842_ _5857_/S vssd1 vssd1 vccd1 vccd1 _5851_/S sky130_fd_sc_hd__buf_2
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5773_ _5559_/X _7852_/Q _5779_/S vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3640_ _7402_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3640_/X sky130_fd_sc_hd__clkbuf_16
X_4724_ _4664_/X _4723_/X _4951_/B vssd1 vssd1 vccd1 vccd1 _4724_/X sky130_fd_sc_hd__a21o_1
X_7512_ _7565_/A _7565_/B _7510_/A vssd1 vssd1 vccd1 vccd1 _7513_/D sky130_fd_sc_hd__a21oi_1
X_8492_ _8527_/CLK _8492_/D vssd1 vssd1 vccd1 vccd1 _8492_/Q sky130_fd_sc_hd__dfxtp_2
X_4655_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4655_/X sky130_fd_sc_hd__clkbuf_4
X_4586_ _5661_/A _4959_/A vssd1 vssd1 vccd1 vccd1 _4602_/S sky130_fd_sc_hd__or2_2
Xinput82 wbs_data_i[20] vssd1 vssd1 vccd1 vccd1 _5946_/A sky130_fd_sc_hd__clkbuf_2
Xinput60 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 _3867_/B sky130_fd_sc_hd__clkbuf_1
Xinput71 wbs_data_i[10] vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__clkbuf_2
X_7374_ _8127_/Q _7679_/B _7366_/X _7373_/X _7371_/X vssd1 vssd1 vccd1 vccd1 _8364_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_1_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput93 wbs_data_i[30] vssd1 vssd1 vccd1 vccd1 _5967_/A sky130_fd_sc_hd__buf_4
XFILLER_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6256_ _7637_/A _7814_/Q _6258_/S vssd1 vssd1 vccd1 vccd1 _6257_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5207_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__buf_2
X_6187_ _7726_/A vssd1 vssd1 vccd1 vccd1 _6367_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5138_ _8440_/Q _8432_/Q _7835_/Q _8448_/Q _5066_/X _5080_/X vssd1 vssd1 vccd1 vccd1
+ _5138_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5069_ _8519_/Q _8072_/Q _8045_/Q _8503_/Q _5066_/X _5068_/X vssd1 vssd1 vccd1 vccd1
+ _5069_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3253_ clkbuf_0__3253_/X vssd1 vssd1 vccd1 vccd1 _6576__265/A sky130_fd_sc_hd__clkbuf_4
X_7039__485 _7039__485/A vssd1 vssd1 vccd1 vccd1 _8212_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6985__444 _6986__445/A vssd1 vssd1 vccd1 vccd1 _8169_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4440_ _4440_/A vssd1 vssd1 vccd1 vccd1 _8263_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4371_ _4371_/A vssd1 vssd1 vccd1 vccd1 _8286_/D sky130_fd_sc_hd__clkbuf_1
X_6110_ _6095_/X _6107_/X _6109_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6110_/X sky130_fd_sc_hd__o211a_1
X_7090_ _7114_/A vssd1 vssd1 vccd1 vccd1 _7090_/X sky130_fd_sc_hd__buf_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6041_ _6138_/A vssd1 vssd1 vccd1 vccd1 _7633_/A sky130_fd_sc_hd__clkbuf_8
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7992_ _7992_/CLK _7992_/D vssd1 vssd1 vccd1 vccd1 _7992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6943_ _6955_/A vssd1 vssd1 vccd1 vccd1 _6943_/X sky130_fd_sc_hd__buf_1
XFILLER_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5825_ _7829_/Q _5554_/A _5833_/S vssd1 vssd1 vccd1 vccd1 _5826_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5756_ _5756_/A vssd1 vssd1 vccd1 vccd1 _7908_/D sky130_fd_sc_hd__clkbuf_1
X_8544_ _8550_/CLK _8544_/D vssd1 vssd1 vccd1 vccd1 _8544_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5687_ _7938_/Q _5650_/X _5689_/S vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__mux2_1
X_4707_ _4654_/X _4704_/X _4706_/X vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__a21o_1
X_8475_ _8479_/CLK _8475_/D vssd1 vssd1 vccd1 vccd1 _8475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7426_ _7426_/A vssd1 vssd1 vccd1 vccd1 _7426_/X sky130_fd_sc_hd__buf_1
X_4638_ _4638_/A vssd1 vssd1 vccd1 vccd1 _4638_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4569_ _3954_/X _8212_/Q _4577_/S vssd1 vssd1 vccd1 vccd1 _4570_/A sky130_fd_sc_hd__mux2_1
X_7357_ _7359_/A _7359_/B _7360_/D _7361_/A vssd1 vssd1 vccd1 vccd1 _7357_/X sky130_fd_sc_hd__a31o_1
X_7288_ _7389_/A vssd1 vssd1 vccd1 vccd1 _7288_/X sky130_fd_sc_hd__buf_1
XFILLER_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6239_ _6239_/A vssd1 vssd1 vccd1 vccd1 _6239_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _3893_/X _8502_/Q _3946_/S vssd1 vssd1 vccd1 vccd1 _3941_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3440_ clkbuf_0__3440_/X vssd1 vssd1 vccd1 vccd1 _7002__457/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3871_ _3871_/A _3871_/B _3871_/C _3871_/D vssd1 vssd1 vccd1 vccd1 _6082_/A sky130_fd_sc_hd__nor4_4
X_5610_ _5610_/A vssd1 vssd1 vccd1 vccd1 _7979_/D sky130_fd_sc_hd__clkbuf_1
X_6590_ _6632_/A vssd1 vssd1 vccd1 vccd1 _6590_/X sky130_fd_sc_hd__buf_1
X_5541_ _5541_/A vssd1 vssd1 vccd1 vccd1 _8028_/D sky130_fd_sc_hd__clkbuf_1
X_8260_ _8260_/CLK _8260_/D vssd1 vssd1 vccd1 vccd1 _8260_/Q sky130_fd_sc_hd__dfxtp_1
X_7424__144 _7425__145/A vssd1 vssd1 vccd1 vccd1 _8401_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5472_ _3969_/X _8058_/Q _5474_/S vssd1 vssd1 vccd1 vccd1 _5473_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7211_ _8348_/Q vssd1 vssd1 vccd1 vccd1 _7227_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3270_ _6632_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3270_/X sky130_fd_sc_hd__clkbuf_16
X_8191_ _8191_/CLK _8191_/D vssd1 vssd1 vccd1 vccd1 _8191_/Q sky130_fd_sc_hd__dfxtp_1
X_4423_ _4423_/A vssd1 vssd1 vccd1 vccd1 _8268_/D sky130_fd_sc_hd__clkbuf_1
X_4354_ _4298_/X _8293_/Q _4354_/S vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _4285_/A vssd1 vssd1 vccd1 vccd1 _8322_/D sky130_fd_sc_hd__clkbuf_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _8014_/Q _6030_/B vssd1 vssd1 vccd1 vccd1 _6025_/A sky130_fd_sc_hd__and2_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7975_ _7975_/CLK _7975_/D vssd1 vssd1 vccd1 vccd1 _7975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6926_ _6932_/A vssd1 vssd1 vccd1 vccd1 _6926_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_0_0__3021_ clkbuf_0__3021_/X vssd1 vssd1 vccd1 vccd1 _7494_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3638_ clkbuf_0__3638_/X vssd1 vssd1 vccd1 vccd1 _7400__125/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6857_ _6857_/A _8475_/Q _8474_/Q _6857_/D vssd1 vssd1 vccd1 vccd1 _6857_/X sky130_fd_sc_hd__and4_1
XFILLER_22_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5808_ _5808_/A vssd1 vssd1 vccd1 vccd1 _7837_/D sky130_fd_sc_hd__clkbuf_1
X_6788_ _8472_/Q _8471_/Q _8470_/Q _8469_/Q vssd1 vssd1 vccd1 vccd1 _6796_/A sky130_fd_sc_hd__and4_1
X_7465__1 _7466__2/A vssd1 vssd1 vccd1 vccd1 _8433_/CLK sky130_fd_sc_hd__inv_2
X_8527_ _8527_/CLK _8527_/D vssd1 vssd1 vccd1 vccd1 _8527_/Q sky130_fd_sc_hd__dfxtp_1
X_5739_ _7915_/Q _5647_/X _5743_/S vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8458_ _8458_/CLK _8458_/D vssd1 vssd1 vccd1 vccd1 _8458_/Q sky130_fd_sc_hd__dfxtp_1
X_8389_ _8389_/CLK _8389_/D vssd1 vssd1 vccd1 vccd1 _8389_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3468_ _7140_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3468_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_40 _6129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_51 _6143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_73 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_95 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_84 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_62 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _4027_/X _8421_/Q _4074_/S vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6998__454 _6998__454/A vssd1 vssd1 vccd1 vccd1 _8179_/CLK sky130_fd_sc_hd__inv_2
X_6740__338 _6740__338/A vssd1 vssd1 vccd1 vccd1 _8048_/CLK sky130_fd_sc_hd__inv_2
X_6289__194 _6290__195/A vssd1 vssd1 vccd1 vccd1 _7824_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4972_ _4972_/A vssd1 vssd1 vccd1 vccd1 _8161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7760_ _7631_/A _7702_/X _7744_/X _7729_/A vssd1 vssd1 vccd1 vccd1 _7760_/X sky130_fd_sc_hd__a31o_1
X_3923_ _3896_/X _8509_/Q _3927_/S vssd1 vssd1 vccd1 vccd1 _3924_/A sky130_fd_sc_hd__mux2_1
X_7691_ _7691_/A vssd1 vssd1 vccd1 vccd1 _8528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3423_ clkbuf_0__3423_/X vssd1 vssd1 vccd1 vccd1 _6930__404/A sky130_fd_sc_hd__clkbuf_4
X_3854_ _4076_/A _8116_/Q vssd1 vssd1 vccd1 vccd1 _5034_/A sky130_fd_sc_hd__xnor2_1
XFILLER_32_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8312_ _8312_/CLK _8312_/D vssd1 vssd1 vccd1 vccd1 _8312_/Q sky130_fd_sc_hd__dfxtp_1
X_5524_ _5396_/X _8035_/Q _5528_/S vssd1 vssd1 vccd1 vccd1 _5525_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5455_ _5455_/A vssd1 vssd1 vccd1 vccd1 _8069_/D sky130_fd_sc_hd__clkbuf_1
X_7144__69 _7145__70/A vssd1 vssd1 vccd1 vccd1 _8296_/CLK sky130_fd_sc_hd__inv_2
X_8243_ _8243_/CLK _8243_/D vssd1 vssd1 vccd1 vccd1 _8243_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3253_ _6571_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3253_/X sky130_fd_sc_hd__clkbuf_16
X_4406_ _4382_/X _8274_/Q _4410_/S vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__mux2_1
X_8174_ _8174_/CLK _8174_/D vssd1 vssd1 vccd1 vccd1 _8174_/Q sky130_fd_sc_hd__dfxtp_1
X_5386_ _8106_/Q vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ _4337_/A vssd1 vssd1 vccd1 vccd1 _8301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4268_ _4268_/A vssd1 vssd1 vccd1 vccd1 _8328_/D sky130_fd_sc_hd__clkbuf_1
X_6007_ _6007_/A vssd1 vssd1 vccd1 vccd1 _6007_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4199_ _5500_/B _4199_/B vssd1 vssd1 vccd1 vccd1 _4215_/S sky130_fd_sc_hd__nor2_2
XFILLER_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ _7958_/CLK _7958_/D vssd1 vssd1 vccd1 vccd1 _7958_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _8485_/Q _6911_/B vssd1 vssd1 vccd1 vccd1 _6910_/A sky130_fd_sc_hd__and2_1
X_7889_ _8520_/CLK _7889_/D vssd1 vssd1 vccd1 vccd1 _7889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5240_ _8319_/Q _8056_/Q _5252_/S vssd1 vssd1 vccd1 vccd1 _5240_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5171_ _5092_/X _5170_/X _5131_/X vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__a21o_1
X_4122_ _6329_/A _6398_/A _6461_/B _6461_/C vssd1 vssd1 vccd1 vccd1 _4122_/Y sky130_fd_sc_hd__nor4_4
XFILLER_96_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4053_ _4031_/X _8428_/Q _4055_/S vssd1 vssd1 vccd1 vccd1 _4054_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 caravel_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7812_ _8355_/CLK _7812_/D vssd1 vssd1 vccd1 vccd1 _7812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7743_ _7754_/B vssd1 vssd1 vccd1 vccd1 _7743_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4955_ _4955_/A _4955_/B vssd1 vssd1 vccd1 vccd1 _4955_/Y sky130_fd_sc_hd__nand2_1
X_3906_ _3905_/X _8514_/Q _3912_/S vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__mux2_1
X_4886_ _4886_/A _4886_/B _4886_/C vssd1 vssd1 vccd1 vccd1 _4886_/X sky130_fd_sc_hd__or3_1
Xclkbuf_1_1_0__3406_ clkbuf_0__3406_/X vssd1 vssd1 vccd1 vccd1 _6873__372/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3837_ _4301_/A vssd1 vssd1 vccd1 vccd1 _4256_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5507_ _5507_/A vssd1 vssd1 vccd1 vccd1 _8043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8226_ _8226_/CLK _8226_/D vssd1 vssd1 vccd1 vccd1 _8226_/Q sky130_fd_sc_hd__dfxtp_1
X_6487_ _5995_/A _7886_/Q _6487_/S vssd1 vssd1 vccd1 vccd1 _6488_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5438_ _3972_/X _8076_/Q _5438_/S vssd1 vssd1 vccd1 vccd1 _5439_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5369_ _5369_/A vssd1 vssd1 vccd1 vccd1 _8104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8157_ _8157_/CLK _8157_/D vssd1 vssd1 vccd1 vccd1 _8157_/Q sky130_fd_sc_hd__dfxtp_1
X_7108_ _7108_/A vssd1 vssd1 vccd1 vccd1 _7108_/X sky130_fd_sc_hd__buf_1
XFILLER_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8088_ _8088_/CLK _8088_/D vssd1 vssd1 vccd1 vccd1 _8088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7437__154 _7438__155/A vssd1 vssd1 vccd1 vccd1 _8411_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4740_/A vssd1 vssd1 vccd1 vccd1 _4740_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4671_ _4714_/A _4668_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _4671_/X sky130_fd_sc_hd__a21o_1
X_6410_ _6854_/A _6444_/C _6410_/C vssd1 vssd1 vccd1 vccd1 _6410_/X sky130_fd_sc_hd__and3_1
X_6341_ _6341_/A _7742_/D vssd1 vssd1 vccd1 vccd1 _6398_/B sky130_fd_sc_hd__or2_1
X_6272_ _6272_/A _6272_/B _6272_/C vssd1 vssd1 vccd1 vccd1 _6272_/X sky130_fd_sc_hd__and3_1
XFILLER_88_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5223_ _5350_/B _5202_/X _5206_/X _5222_/X vssd1 vssd1 vccd1 vccd1 _5223_/X sky130_fd_sc_hd__a31o_1
X_8011_ _8531_/CLK _8011_/D vssd1 vssd1 vccd1 vccd1 _8011_/Q sky130_fd_sc_hd__dfxtp_4
X_5154_ _5047_/X _5140_/X _5144_/X _5153_/X vssd1 vssd1 vccd1 vccd1 _5154_/X sky130_fd_sc_hd__a31o_2
Xclkbuf_0__3021_ _6163_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3021_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4105_ _4105_/A vssd1 vssd1 vccd1 vccd1 _8407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5085_ _5055_/X _5078_/X _5084_/X vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4036_ _4035_/X _8435_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5987_ _5987_/A vssd1 vssd1 vccd1 vccd1 _5987_/X sky130_fd_sc_hd__clkbuf_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7726_ _7726_/A vssd1 vssd1 vccd1 vccd1 _7729_/A sky130_fd_sc_hd__buf_2
X_4938_ _4938_/A vssd1 vssd1 vccd1 vccd1 _8176_/D sky130_fd_sc_hd__clkbuf_1
X_4869_ _4811_/A _7951_/Q _7764_/Q _4797_/X _4663_/A vssd1 vssd1 vccd1 vccd1 _4869_/X
+ sky130_fd_sc_hd__o221a_1
X_6608_ _6608_/A vssd1 vssd1 vccd1 vccd1 _7966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7588_ _7588_/A vssd1 vssd1 vccd1 vccd1 _7588_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput170 _5889_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[0] sky130_fd_sc_hd__buf_2
XFILLER_79_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8209_ _8209_/CLK _8209_/D vssd1 vssd1 vccd1 vccd1 _8209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput192 _6132_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput181 _6094_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[13] sky130_fd_sc_hd__buf_2
XFILLER_48_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3467_ clkbuf_0__3467_/X vssd1 vssd1 vccd1 vccd1 _7139__65/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6550__244 _6551__245/A vssd1 vssd1 vccd1 vccd1 _7922_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5910_ _7640_/A _5910_/B vssd1 vssd1 vccd1 vccd1 _5911_/A sky130_fd_sc_hd__or2_1
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6890_ _6890_/A vssd1 vssd1 vccd1 vccd1 _6890_/X sky130_fd_sc_hd__buf_1
XFILLER_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5841_ _5841_/A _5859_/B vssd1 vssd1 vccd1 vccd1 _5857_/S sky130_fd_sc_hd__or2_2
XFILLER_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5772_ _5772_/A vssd1 vssd1 vccd1 vccd1 _7853_/D sky130_fd_sc_hd__clkbuf_1
X_4723_ _8140_/Q _8027_/Q _7923_/Q _7907_/Q _4655_/X _4656_/X vssd1 vssd1 vccd1 vccd1
+ _4723_/X sky130_fd_sc_hd__mux4_1
X_7511_ _7571_/A _7571_/B _8544_/Q vssd1 vssd1 vccd1 vccd1 _7513_/C sky130_fd_sc_hd__a21boi_1
X_8491_ _8530_/CLK _8491_/D vssd1 vssd1 vccd1 vccd1 _8491_/Q sky130_fd_sc_hd__dfxtp_2
X_4654_ _4654_/A vssd1 vssd1 vccd1 vccd1 _4654_/X sky130_fd_sc_hd__buf_2
XFILLER_116_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4585_ _5841_/A vssd1 vssd1 vccd1 vccd1 _5661_/A sky130_fd_sc_hd__buf_4
X_7489__21 _7490__22/A vssd1 vssd1 vccd1 vccd1 _8453_/CLK sky130_fd_sc_hd__inv_2
Xinput61 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 _3867_/A sky130_fd_sc_hd__clkbuf_1
Xinput50 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _3866_/C sky130_fd_sc_hd__clkbuf_1
Xinput72 wbs_data_i[11] vssd1 vssd1 vccd1 vccd1 _5926_/A sky130_fd_sc_hd__clkbuf_2
X_7373_ _8364_/Q _7377_/B vssd1 vssd1 vccd1 vccd1 _7373_/X sky130_fd_sc_hd__or2_1
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput83 wbs_data_i[21] vssd1 vssd1 vccd1 vccd1 _5948_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput94 wbs_data_i[31] vssd1 vssd1 vccd1 vccd1 _5969_/A sky130_fd_sc_hd__buf_4
X_6255_ _6255_/A vssd1 vssd1 vccd1 vccd1 _7813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5206_ _5206_/A _5206_/B vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__or2_1
XFILLER_69_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6186_ _6247_/A vssd1 vssd1 vccd1 vccd1 _7726_/A sky130_fd_sc_hd__clkbuf_4
X_5137_ _8408_/Q _8392_/Q _8384_/Q _8416_/Q _5284_/S _5061_/X vssd1 vssd1 vccd1 vccd1
+ _5137_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5068_ _5080_/A vssd1 vssd1 vccd1 vccd1 _5068_/X sky130_fd_sc_hd__buf_2
X_4019_ _4286_/A vssd1 vssd1 vccd1 vccd1 _4019_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3252_ clkbuf_0__3252_/X vssd1 vssd1 vccd1 vccd1 _6568__258/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7709_ _8533_/Q _7701_/X _7708_/X _7704_/X vssd1 vssd1 vccd1 vccd1 _8533_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _4295_/X _8286_/Q _4372_/S vssd1 vssd1 vccd1 vccd1 _4371_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6040_ _6108_/A vssd1 vssd1 vccd1 vccd1 _6138_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7991_ _7991_/CLK _7991_/D vssd1 vssd1 vccd1 vccd1 _7991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6942_ _6942_/A vssd1 vssd1 vccd1 vccd1 _8134_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3654_ clkbuf_0__3654_/X vssd1 vssd1 vccd1 vccd1 _7479__13/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_16_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8537_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5824_ _5839_/S vssd1 vssd1 vccd1 vccd1 _5833_/S sky130_fd_sc_hd__buf_2
X_5755_ _7908_/Q _5559_/A _5761_/S vssd1 vssd1 vccd1 vccd1 _5756_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8543_ _8543_/CLK _8543_/D vssd1 vssd1 vccd1 vccd1 _8543_/Q sky130_fd_sc_hd__dfxtp_1
X_5686_ _5686_/A vssd1 vssd1 vccd1 vccd1 _7939_/D sky130_fd_sc_hd__clkbuf_1
X_4706_ _4677_/S _4705_/X _4694_/A vssd1 vssd1 vccd1 vccd1 _4706_/X sky130_fd_sc_hd__a21o_1
X_8474_ _8479_/CLK _8474_/D vssd1 vssd1 vccd1 vccd1 _8474_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4637_ _8172_/Q _4683_/B vssd1 vssd1 vccd1 vccd1 _4638_/A sky130_fd_sc_hd__xor2_4
XFILLER_118_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4568_ _4583_/S vssd1 vssd1 vccd1 vccd1 _4577_/S sky130_fd_sc_hd__buf_2
X_7356_ _8360_/Q _7356_/B vssd1 vssd1 vccd1 vccd1 _7360_/D sky130_fd_sc_hd__nand2_1
XFILLER_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4499_ _4499_/A vssd1 vssd1 vccd1 vccd1 _8241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7287_ _7271_/Y _7269_/C _7285_/X _7286_/X vssd1 vssd1 vccd1 vccd1 _8334_/D sky130_fd_sc_hd__o211a_1
X_7045__490 _7045__490/A vssd1 vssd1 vccd1 vccd1 _8217_/CLK sky130_fd_sc_hd__inv_2
X_6238_ _6367_/A vssd1 vssd1 vccd1 vccd1 _6238_/X sky130_fd_sc_hd__clkbuf_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7087__524 _7087__524/A vssd1 vssd1 vccd1 vccd1 _8251_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7483__16 _7485__18/A vssd1 vssd1 vccd1 vccd1 _8448_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3870_ _3870_/A _3870_/B _3870_/C vssd1 vssd1 vccd1 vccd1 _3871_/D sky130_fd_sc_hd__or3_4
X_5540_ _5367_/X _8028_/Q _5546_/S vssd1 vssd1 vccd1 vccd1 _5541_/A sky130_fd_sc_hd__mux2_1
X_5471_ _5471_/A vssd1 vssd1 vccd1 vccd1 _8059_/D sky130_fd_sc_hd__clkbuf_1
X_7156__78 _7156__78/A vssd1 vssd1 vccd1 vccd1 _8305_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4422_ _4418_/X _8268_/Q _4436_/S vssd1 vssd1 vccd1 vccd1 _4423_/A sky130_fd_sc_hd__mux2_1
X_7210_ _7210_/A _7210_/B vssd1 vssd1 vccd1 vccd1 _7272_/B sky130_fd_sc_hd__nand2_1
X_8190_ _8190_/CLK _8190_/D vssd1 vssd1 vccd1 vccd1 _8190_/Q sky130_fd_sc_hd__dfxtp_1
X_4353_ _4353_/A vssd1 vssd1 vccd1 vccd1 _8294_/D sky130_fd_sc_hd__clkbuf_1
X_4284_ _4283_/X _8322_/Q _4290_/S vssd1 vssd1 vccd1 vccd1 _4285_/A sky130_fd_sc_hd__mux2_1
X_6023_ _6023_/A vssd1 vssd1 vccd1 vccd1 _6023_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6563__254 _6563__254/A vssd1 vssd1 vccd1 vccd1 _7932_/CLK sky130_fd_sc_hd__inv_2
X_7974_ _7974_/CLK _7974_/D vssd1 vssd1 vccd1 vccd1 _7974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6925_ _6925_/A vssd1 vssd1 vccd1 vccd1 _6925_/X sky130_fd_sc_hd__buf_1
XFILLER_42_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3637_ clkbuf_0__3637_/X vssd1 vssd1 vccd1 vccd1 _7394__120/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6856_ _8476_/Q vssd1 vssd1 vccd1 vccd1 _6857_/A sky130_fd_sc_hd__inv_2
X_5807_ _3954_/X _7837_/Q _5815_/S vssd1 vssd1 vccd1 vccd1 _5808_/A sky130_fd_sc_hd__mux2_1
X_3999_ _3999_/A vssd1 vssd1 vccd1 vccd1 _8445_/D sky130_fd_sc_hd__clkbuf_1
X_6787_ _7497_/A vssd1 vssd1 vccd1 vccd1 _7505_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8526_ _8526_/CLK _8526_/D vssd1 vssd1 vccd1 vccd1 _8526_/Q sky130_fd_sc_hd__dfxtp_1
X_5738_ _5738_/A vssd1 vssd1 vccd1 vccd1 _7916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5669_ _5611_/X _7946_/Q _5671_/S vssd1 vssd1 vccd1 vccd1 _5670_/A sky130_fd_sc_hd__mux2_1
X_8457_ _8457_/CLK _8457_/D vssd1 vssd1 vccd1 vccd1 _8457_/Q sky130_fd_sc_hd__dfxtp_1
X_7408_ _7420_/A vssd1 vssd1 vccd1 vccd1 _7408_/X sky130_fd_sc_hd__buf_1
X_8388_ _8388_/CLK _8388_/D vssd1 vssd1 vccd1 vccd1 _8388_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3467_ _7134_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3467_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7339_ _7348_/A _7339_/B vssd1 vssd1 vccd1 vccd1 _8354_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_52 _6143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_30 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_41 _6131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_74 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_63 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_85 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_96 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6876__375 _6876__375/A vssd1 vssd1 vccd1 vccd1 _8089_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6917__394 _6918__395/A vssd1 vssd1 vccd1 vccd1 _8116_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4971_ _8161_/Q _4481_/X _4975_/S vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3922_ _3922_/A vssd1 vssd1 vccd1 vccd1 _8510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7690_ _7719_/A _8522_/Q vssd1 vssd1 vccd1 vccd1 _7691_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3422_ clkbuf_0__3422_/X vssd1 vssd1 vccd1 vccd1 _6955_/A sky130_fd_sc_hd__clkbuf_4
X_3853_ _3853_/A _5035_/B vssd1 vssd1 vccd1 vccd1 _3853_/Y sky130_fd_sc_hd__nor2_1
X_8311_ _8311_/CLK _8311_/D vssd1 vssd1 vccd1 vccd1 _8311_/Q sky130_fd_sc_hd__dfxtp_1
X_7129__56 _7130__57/A vssd1 vssd1 vccd1 vccd1 _8283_/CLK sky130_fd_sc_hd__inv_2
X_5523_ _5523_/A vssd1 vssd1 vccd1 vccd1 _8036_/D sky130_fd_sc_hd__clkbuf_1
X_5454_ _8069_/Q _4184_/X _5456_/S vssd1 vssd1 vccd1 vccd1 _5455_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3321_ _6780_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3321_/X sky130_fd_sc_hd__clkbuf_16
X_8242_ _8242_/CLK _8242_/D vssd1 vssd1 vccd1 vccd1 _8242_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3252_ _6565_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3252_/X sky130_fd_sc_hd__clkbuf_16
X_5385_ _5385_/A vssd1 vssd1 vccd1 vccd1 _8099_/D sky130_fd_sc_hd__clkbuf_1
X_4405_ _4405_/A vssd1 vssd1 vccd1 vccd1 _8275_/D sky130_fd_sc_hd__clkbuf_1
X_8173_ _8173_/CLK _8173_/D vssd1 vssd1 vccd1 vccd1 _8173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4336_ _4298_/X _8301_/Q _4336_/S vssd1 vssd1 vccd1 vccd1 _4337_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4267_ _8328_/Q _4187_/X _4267_/S vssd1 vssd1 vccd1 vccd1 _4268_/A sky130_fd_sc_hd__mux2_1
X_6006_ _8006_/Q _6008_/B vssd1 vssd1 vccd1 vccd1 _6007_/A sky130_fd_sc_hd__and2_1
X_4198_ _4198_/A vssd1 vssd1 vccd1 vccd1 _8387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6309__210 _6309__210/A vssd1 vssd1 vccd1 vccd1 _7840_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7957_ _7957_/CLK _7957_/D vssd1 vssd1 vccd1 vccd1 _7957_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7888_ _8063_/CLK _7888_/D vssd1 vssd1 vccd1 vccd1 _7888_/Q sky130_fd_sc_hd__dfxtp_1
X_6908_ _6908_/A vssd1 vssd1 vccd1 vccd1 _8110_/D sky130_fd_sc_hd__clkbuf_1
X_6839_ _7556_/A _7556_/B _6838_/A vssd1 vssd1 vccd1 vccd1 _6839_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8509_ _8509_/CLK _8509_/D vssd1 vssd1 vccd1 vccd1 _8509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5170_ _8209_/Q _8193_/Q _8455_/Q _8225_/Q _5231_/S _5129_/X vssd1 vssd1 vccd1 vccd1
+ _5170_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4121_ _6417_/A _6517_/A vssd1 vssd1 vccd1 vccd1 _6329_/A sky130_fd_sc_hd__or2b_1
X_4052_ _4052_/A vssd1 vssd1 vccd1 vccd1 _8429_/D sky130_fd_sc_hd__clkbuf_1
Xinput4 caravel_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7811_ _8355_/CLK _7811_/D vssd1 vssd1 vccd1 vccd1 _7811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7742_ _7742_/A _7742_/B _7742_/C _7742_/D vssd1 vssd1 vccd1 vccd1 _7754_/B sky130_fd_sc_hd__nor4_2
X_4954_ _4811_/X _4947_/X _4953_/Y _4924_/X vssd1 vssd1 vccd1 vccd1 _8170_/D sky130_fd_sc_hd__o211a_1
X_3905_ _8490_/Q vssd1 vssd1 vccd1 vccd1 _3905_/X sky130_fd_sc_hd__buf_4
X_4885_ _4809_/A _4883_/X _4884_/X vssd1 vssd1 vccd1 vccd1 _4886_/C sky130_fd_sc_hd__o21a_1
XFILLER_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3836_ _8123_/Q vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5506_ _8043_/Q _4283_/A _5510_/S vssd1 vssd1 vccd1 vccd1 _5507_/A sky130_fd_sc_hd__mux2_1
X_8225_ _8225_/CLK _8225_/D vssd1 vssd1 vccd1 vccd1 _8225_/Q sky130_fd_sc_hd__dfxtp_1
X_6486_ _6486_/A vssd1 vssd1 vccd1 vccd1 _7885_/D sky130_fd_sc_hd__clkbuf_1
X_5437_ _5437_/A vssd1 vssd1 vccd1 vccd1 _8077_/D sky130_fd_sc_hd__clkbuf_1
X_5368_ _5367_/X _8104_/Q _5376_/S vssd1 vssd1 vccd1 vccd1 _5369_/A sky130_fd_sc_hd__mux2_1
X_8156_ _8156_/CLK _8156_/D vssd1 vssd1 vccd1 vccd1 _8156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4319_ _4319_/A vssd1 vssd1 vccd1 vccd1 _8309_/D sky130_fd_sc_hd__clkbuf_1
X_5299_ _5306_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _5299_/X sky130_fd_sc_hd__or2_1
X_8087_ _8087_/CLK _8087_/D vssd1 vssd1 vccd1 vccd1 _8087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8572__219 vssd1 vssd1 vccd1 vccd1 _8572__219/HI core0Index[6] sky130_fd_sc_hd__conb_1
XFILLER_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4670_ _4740_/A vssd1 vssd1 vccd1 vccd1 _4670_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__3275_ clkbuf_0__3275_/X vssd1 vssd1 vccd1 vccd1 _6711__315/A sky130_fd_sc_hd__clkbuf_16
X_6340_ _7878_/Q _6348_/B _6348_/C vssd1 vssd1 vccd1 vccd1 _7742_/D sky130_fd_sc_hd__or3_1
X_6889__385 _6889__385/A vssd1 vssd1 vccd1 vccd1 _8099_/CLK sky130_fd_sc_hd__inv_2
X_6271_ _6271_/A vssd1 vssd1 vccd1 vccd1 _7819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5222_ _5293_/A _5210_/X _5213_/X _5221_/X _5047_/X vssd1 vssd1 vccd1 vccd1 _5222_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8010_ _8531_/CLK _8010_/D vssd1 vssd1 vccd1 vccd1 _8010_/Q sky130_fd_sc_hd__dfxtp_4
X_5153_ _5293_/A _5148_/X _5150_/X _5152_/X _5177_/A vssd1 vssd1 vccd1 vccd1 _5153_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4104_ _4019_/X _8407_/Q _4106_/S vssd1 vssd1 vccd1 vccd1 _4105_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5084_ _5079_/X _5081_/X _5083_/X vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4035_ _4298_/A vssd1 vssd1 vccd1 vccd1 _4035_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5986_ _5986_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _5987_/A sky130_fd_sc_hd__and2_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7725_ _7528_/A _7717_/X _7724_/X _7719_/X vssd1 vssd1 vccd1 vccd1 _8538_/D sky130_fd_sc_hd__o211a_1
X_4937_ _7008_/C _4937_/B _4937_/C vssd1 vssd1 vccd1 vccd1 _4938_/A sky130_fd_sc_hd__and3_1
X_4868_ _7847_/Q _7772_/Q _4868_/S vssd1 vssd1 vccd1 vccd1 _4868_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6753__349 _6753__349/A vssd1 vssd1 vccd1 vccd1 _8059_/CLK sky130_fd_sc_hd__inv_2
X_6607_ _8179_/Q _8167_/D vssd1 vssd1 vccd1 vccd1 _6608_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3319_ clkbuf_0__3319_/X vssd1 vssd1 vccd1 vccd1 _6772__359/A sky130_fd_sc_hd__clkbuf_4
X_4799_ _4794_/X _4795_/X _4798_/X vssd1 vssd1 vccd1 vccd1 _4799_/X sky130_fd_sc_hd__o21a_1
X_7587_ _8472_/Q vssd1 vssd1 vccd1 vccd1 _7587_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7081__519 _7082__520/A vssd1 vssd1 vccd1 vccd1 _8246_/CLK sky130_fd_sc_hd__inv_2
X_6469_ _6469_/A vssd1 vssd1 vccd1 vccd1 _7877_/D sky130_fd_sc_hd__clkbuf_1
Xoutput160 _5907_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[2] sky130_fd_sc_hd__buf_2
X_8208_ _8208_/CLK _8208_/D vssd1 vssd1 vccd1 vccd1 _8208_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput171 _5891_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[1] sky130_fd_sc_hd__buf_2
XFILLER_99_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8139_ _8139_/CLK _8139_/D vssd1 vssd1 vccd1 vccd1 _8139_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput193 _6134_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput182 _6099_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[14] sky130_fd_sc_hd__buf_2
XFILLER_102_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3466_ clkbuf_0__3466_/X vssd1 vssd1 vccd1 vccd1 _7133__60/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6769__356 _6773__360/A vssd1 vssd1 vccd1 vccd1 _8069_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8594__241 vssd1 vssd1 vccd1 vccd1 _8594__241/HI partID[5] sky130_fd_sc_hd__conb_1
X_5840_ _5840_/A vssd1 vssd1 vccd1 vccd1 _7822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5771_ _5554_/X _7853_/Q _5779_/S vssd1 vssd1 vccd1 vccd1 _5772_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7510_ _7510_/A _7565_/A _7565_/B vssd1 vssd1 vccd1 vccd1 _7513_/B sky130_fd_sc_hd__and3_1
X_4722_ _8095_/Q _8087_/Q _7915_/Q _8156_/Q _4646_/X _4716_/X vssd1 vssd1 vccd1 vccd1
+ _4722_/X sky130_fd_sc_hd__mux4_1
X_8490_ _8527_/CLK _8490_/D vssd1 vssd1 vccd1 vccd1 _8490_/Q sky130_fd_sc_hd__dfxtp_2
X_4653_ _4663_/A vssd1 vssd1 vccd1 vccd1 _4654_/A sky130_fd_sc_hd__clkbuf_2
Xinput40 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 _5997_/A sky130_fd_sc_hd__buf_4
X_4584_ _4584_/A vssd1 vssd1 vccd1 vccd1 _8205_/D sky130_fd_sc_hd__clkbuf_1
Xinput51 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 _3869_/B sky130_fd_sc_hd__clkbuf_1
Xinput62 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _5978_/A sky130_fd_sc_hd__buf_4
Xinput73 wbs_data_i[12] vssd1 vssd1 vccd1 vccd1 _7728_/A sky130_fd_sc_hd__clkbuf_2
X_7372_ _8126_/Q _7679_/B _7366_/X _7370_/X _7371_/X vssd1 vssd1 vccd1 vccd1 _8363_/D
+ sky130_fd_sc_hd__o311a_1
Xinput84 wbs_data_i[22] vssd1 vssd1 vccd1 vccd1 _5950_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput95 wbs_data_i[3] vssd1 vssd1 vccd1 vccd1 _7637_/A sky130_fd_sc_hd__buf_6
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6254_ _7635_/A _7813_/Q _6258_/S vssd1 vssd1 vccd1 vccd1 _6255_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5205_ _5203_/X _5204_/X _5205_/S vssd1 vssd1 vccd1 vccd1 _5206_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5136_ _3893_/X _5038_/X _5135_/X _5111_/X vssd1 vssd1 vccd1 vccd1 _8131_/D sky130_fd_sc_hd__o211a_1
XFILLER_96_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3320_ clkbuf_0__3320_/X vssd1 vssd1 vccd1 vccd1 _6777__363/A sky130_fd_sc_hd__clkbuf_4
X_5067_ _5181_/A vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__buf_4
Xclkbuf_1_0_0__3251_ clkbuf_0__3251_/X vssd1 vssd1 vccd1 vccd1 _6564__255/A sky130_fd_sc_hd__clkbuf_4
X_4018_ _8492_/Q vssd1 vssd1 vccd1 vccd1 _4286_/A sky130_fd_sc_hd__buf_4
XFILLER_44_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5969_ _5969_/A _5969_/B vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__or2_1
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7708_ _5941_/A _7702_/X _7701_/A vssd1 vssd1 vccd1 vccd1 _7708_/X sky130_fd_sc_hd__a21bo_1
X_7639_ _7702_/A vssd1 vssd1 vccd1 vccd1 _7646_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8578__225 vssd1 vssd1 vccd1 vccd1 _8578__225/HI core1Index[5] sky130_fd_sc_hd__conb_1
XFILLER_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3449_ clkbuf_0__3449_/X vssd1 vssd1 vccd1 vccd1 _7051__495/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7990_ _7990_/CLK _7990_/D vssd1 vssd1 vccd1 vccd1 _7990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6941_ _8370_/Q _6941_/B _6941_/C _7008_/A vssd1 vssd1 vccd1 vccd1 _6942_/A sky130_fd_sc_hd__and4b_1
XFILLER_35_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3653_ clkbuf_0__3653_/X vssd1 vssd1 vccd1 vccd1 _7474__9/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5823_ _5823_/A _5823_/B vssd1 vssd1 vccd1 vccd1 _5839_/S sky130_fd_sc_hd__nor2_2
X_6303__205 _6303__205/A vssd1 vssd1 vccd1 vccd1 _7835_/CLK sky130_fd_sc_hd__inv_2
X_8542_ _8543_/CLK _8542_/D vssd1 vssd1 vccd1 vccd1 _8542_/Q sky130_fd_sc_hd__dfxtp_4
X_5754_ _5754_/A vssd1 vssd1 vccd1 vccd1 _7909_/D sky130_fd_sc_hd__clkbuf_1
X_4705_ _7828_/Q _7948_/Q _7964_/Q _7932_/Q _4876_/A _4649_/A vssd1 vssd1 vccd1 vccd1
+ _4705_/X sky130_fd_sc_hd__mux4_2
X_5685_ _7939_/Q _5647_/X _5689_/S vssd1 vssd1 vccd1 vccd1 _5686_/A sky130_fd_sc_hd__mux2_1
X_8473_ _8473_/CLK _8473_/D vssd1 vssd1 vccd1 vccd1 _8473_/Q sky130_fd_sc_hd__dfxtp_1
X_4636_ _4636_/A vssd1 vssd1 vccd1 vccd1 _4683_/B sky130_fd_sc_hd__buf_2
X_7355_ _7355_/A vssd1 vssd1 vccd1 vccd1 _7359_/B sky130_fd_sc_hd__inv_2
X_4567_ _4567_/A _4604_/A vssd1 vssd1 vccd1 vccd1 _4583_/S sky130_fd_sc_hd__or2_2
XFILLER_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4498_ _4385_/X _8241_/Q _4500_/S vssd1 vssd1 vccd1 vccd1 _4499_/A sky130_fd_sc_hd__mux2_1
X_7286_ _7286_/A vssd1 vssd1 vccd1 vccd1 _7286_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6237_ _8014_/Q _7680_/A _6236_/X _6229_/X _7803_/Q vssd1 vssd1 vccd1 vccd1 _7803_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_103_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _8518_/Q _8071_/Q _8044_/Q _8502_/Q _5290_/S _5080_/X vssd1 vssd1 vccd1 vccd1
+ _5119_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6099_ _6095_/X _6097_/X _6098_/X _6083_/X vssd1 vssd1 vccd1 vccd1 _6099_/X sky130_fd_sc_hd__o211a_1
XFILLER_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7289__106 _7290__107/A vssd1 vssd1 vccd1 vccd1 _8335_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7094__529 _7095__530/A vssd1 vssd1 vccd1 vccd1 _8256_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5470_ _3966_/X _8059_/Q _5474_/S vssd1 vssd1 vccd1 vccd1 _5471_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4421_ _4445_/S vssd1 vssd1 vccd1 vccd1 _4436_/S sky130_fd_sc_hd__clkbuf_2
X_6968__430 _6968__430/A vssd1 vssd1 vccd1 vccd1 _8154_/CLK sky130_fd_sc_hd__inv_2
X_6929__403 _6931__405/A vssd1 vssd1 vccd1 vccd1 _8125_/CLK sky130_fd_sc_hd__inv_2
X_6710__314 _6711__315/A vssd1 vssd1 vccd1 vccd1 _8024_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4352_ _4295_/X _8294_/Q _4354_/S vssd1 vssd1 vccd1 vccd1 _4353_/A sky130_fd_sc_hd__mux2_1
X_7140_ _7146_/A vssd1 vssd1 vccd1 vccd1 _7140_/X sky130_fd_sc_hd__buf_1
XFILLER_86_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4283_ _4283_/A vssd1 vssd1 vccd1 vccd1 _4283_/X sky130_fd_sc_hd__clkbuf_2
X_7071_ _7077_/A vssd1 vssd1 vccd1 vccd1 _7071_/X sky130_fd_sc_hd__buf_1
XFILLER_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _8013_/Q _6030_/B vssd1 vssd1 vccd1 vccd1 _6023_/A sky130_fd_sc_hd__and2_2
XFILLER_100_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7973_ _8520_/CLK _7973_/D vssd1 vssd1 vccd1 vccd1 _7973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6855_ _6855_/A _6855_/B _6855_/C _6855_/D vssd1 vssd1 vccd1 vccd1 _6860_/C sky130_fd_sc_hd__and4_1
X_5806_ _5821_/S vssd1 vssd1 vccd1 vccd1 _5815_/S sky130_fd_sc_hd__buf_2
X_3998_ _3905_/X _8445_/Q _4002_/S vssd1 vssd1 vccd1 vccd1 _3999_/A sky130_fd_sc_hd__mux2_1
X_6786_ _8460_/Q vssd1 vssd1 vccd1 vccd1 _7497_/A sky130_fd_sc_hd__inv_2
XFILLER_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5737_ _7916_/Q _5559_/A _5743_/S vssd1 vssd1 vccd1 vccd1 _5738_/A sky130_fd_sc_hd__mux2_1
X_8525_ _8526_/CLK _8525_/D vssd1 vssd1 vccd1 vccd1 _8525_/Q sky130_fd_sc_hd__dfxtp_1
X_8456_ _8456_/CLK _8456_/D vssd1 vssd1 vccd1 vccd1 _8456_/Q sky130_fd_sc_hd__dfxtp_1
X_5668_ _5668_/A vssd1 vssd1 vccd1 vccd1 _7947_/D sky130_fd_sc_hd__clkbuf_1
X_8387_ _8387_/CLK _8387_/D vssd1 vssd1 vccd1 vccd1 _8387_/Q sky130_fd_sc_hd__dfxtp_1
X_4619_ _4619_/A vssd1 vssd1 vccd1 vccd1 _8190_/D sky130_fd_sc_hd__clkbuf_1
X_5599_ _8106_/Q vssd1 vssd1 vccd1 vccd1 _5599_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3466_ _7128_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3466_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7338_ _8354_/Q _7334_/X _7326_/X _7254_/B vssd1 vssd1 vccd1 vccd1 _7339_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_2_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7269_ _7286_/A _7269_/B _7269_/C vssd1 vssd1 vccd1 vccd1 _7270_/A sky130_fd_sc_hd__and3_1
XFILLER_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_20 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_42 _6131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_31 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_75 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_64 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_86 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_53 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_97 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _8345_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7161__82 _7163__84/A vssd1 vssd1 vccd1 vccd1 _8309_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4970_ _4970_/A vssd1 vssd1 vccd1 vccd1 _8162_/D sky130_fd_sc_hd__clkbuf_1
X_3921_ _3893_/X _8510_/Q _3927_/S vssd1 vssd1 vccd1 vccd1 _3922_/A sky130_fd_sc_hd__mux2_1
X_6640_ _6652_/A vssd1 vssd1 vccd1 vccd1 _6640_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3421_ clkbuf_0__3421_/X vssd1 vssd1 vccd1 vccd1 _6923__399/A sky130_fd_sc_hd__clkbuf_4
X_3852_ _5070_/A _8122_/Q vssd1 vssd1 vccd1 vccd1 _5035_/B sky130_fd_sc_hd__and2b_1
X_6571_ _6571_/A vssd1 vssd1 vccd1 vccd1 _6571_/X sky130_fd_sc_hd__buf_1
XFILLER_118_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5522_ _5367_/X _8036_/Q _5528_/S vssd1 vssd1 vccd1 vccd1 _5523_/A sky130_fd_sc_hd__mux2_1
X_8310_ _8310_/CLK _8310_/D vssd1 vssd1 vccd1 vccd1 _8310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5453_ _5453_/A vssd1 vssd1 vccd1 vccd1 _8070_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3320_ _6774_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3320_/X sky130_fd_sc_hd__clkbuf_16
X_8241_ _8241_/CLK _8241_/D vssd1 vssd1 vccd1 vccd1 _8241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3251_ _6559_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3251_/X sky130_fd_sc_hd__clkbuf_16
X_5384_ _5383_/X _8099_/Q _5388_/S vssd1 vssd1 vccd1 vccd1 _5385_/A sky130_fd_sc_hd__mux2_1
X_4404_ _4379_/X _8275_/Q _4410_/S vssd1 vssd1 vccd1 vccd1 _4405_/A sky130_fd_sc_hd__mux2_1
X_8172_ _8172_/CLK _8172_/D vssd1 vssd1 vccd1 vccd1 _8172_/Q sky130_fd_sc_hd__dfxtp_4
X_4335_ _4335_/A vssd1 vssd1 vccd1 vccd1 _8302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4266_ _4266_/A vssd1 vssd1 vccd1 vccd1 _8329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6005_ _6005_/A vssd1 vssd1 vccd1 vccd1 _6005_/X sky130_fd_sc_hd__clkbuf_1
X_4197_ _8387_/Q _4196_/X _4197_/S vssd1 vssd1 vccd1 vccd1 _4198_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7956_ _7956_/CLK _7956_/D vssd1 vssd1 vccd1 vccd1 _7956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6907_ _8484_/Q _6911_/B vssd1 vssd1 vccd1 vccd1 _6908_/A sky130_fd_sc_hd__and2_1
X_7887_ _8063_/CLK _7887_/D vssd1 vssd1 vccd1 vccd1 _7887_/Q sky130_fd_sc_hd__dfxtp_1
X_6838_ _6838_/A _7556_/A _7556_/B vssd1 vssd1 vccd1 vccd1 _6838_/X sky130_fd_sc_hd__and3_1
XFILLER_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8508_ _8508_/CLK _8508_/D vssd1 vssd1 vccd1 vccd1 _8508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7407__130 _7407__130/A vssd1 vssd1 vccd1 vccd1 _8387_/CLK sky130_fd_sc_hd__inv_2
X_8439_ _8439_/CLK _8439_/D vssd1 vssd1 vccd1 vccd1 _8439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3449_ _7046_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3449_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6169__178 _6170__179/A vssd1 vssd1 vccd1 vccd1 _7765_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4120_ _8173_/Q vssd1 vssd1 vccd1 vccd1 _4944_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4051_ _4027_/X _8429_/Q _4055_/S vssd1 vssd1 vccd1 vccd1 _4052_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput5 caravel_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
X_7810_ _8479_/CLK _7810_/D vssd1 vssd1 vccd1 vccd1 _7810_/Q sky130_fd_sc_hd__dfxtp_1
X_8558__256 vssd1 vssd1 vccd1 vccd1 partID[10] _8558__256/LO sky130_fd_sc_hd__conb_1
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7741_ _7741_/A vssd1 vssd1 vccd1 vccd1 _7742_/A sky130_fd_sc_hd__inv_2
X_4953_ _4955_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _4953_/Y sky130_fd_sc_hd__nand2_1
X_3904_ _3904_/A vssd1 vssd1 vccd1 vccd1 _8515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4884_ _4805_/A _7903_/Q _4806_/A _8136_/Q _4663_/A vssd1 vssd1 vccd1 vccd1 _4884_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3835_ _4057_/B vssd1 vssd1 vccd1 vccd1 _5334_/A sky130_fd_sc_hd__buf_2
XFILLER_20_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5505_ _5505_/A vssd1 vssd1 vccd1 vccd1 _8044_/D sky130_fd_sc_hd__clkbuf_1
X_6485_ _5993_/A _7885_/Q _6487_/S vssd1 vssd1 vccd1 vccd1 _6486_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5436_ _3969_/X _8077_/Q _5438_/S vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__mux2_1
X_8224_ _8224_/CLK _8224_/D vssd1 vssd1 vccd1 vccd1 _8224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5367_ _5559_/A vssd1 vssd1 vccd1 vccd1 _5367_/X sky130_fd_sc_hd__clkbuf_4
X_8155_ _8155_/CLK _8155_/D vssd1 vssd1 vccd1 vccd1 _8155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5298_ _8451_/Q _8189_/Q _5308_/S vssd1 vssd1 vccd1 vccd1 _5299_/B sky130_fd_sc_hd__mux2_1
X_4318_ _4298_/X _8309_/Q _4318_/S vssd1 vssd1 vccd1 vccd1 _4319_/A sky130_fd_sc_hd__mux2_1
X_8086_ _8086_/CLK _8086_/D vssd1 vssd1 vccd1 vccd1 _8086_/Q sky130_fd_sc_hd__dfxtp_1
X_4249_ _4249_/A vssd1 vssd1 vccd1 vccd1 _8338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _7939_/CLK _7939_/D vssd1 vssd1 vccd1 vccd1 _7939_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6576__265 _6576__265/A vssd1 vssd1 vccd1 vccd1 _7943_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6270_ _6273_/B _6270_/B _6272_/C vssd1 vssd1 vccd1 vccd1 _6271_/A sky130_fd_sc_hd__and3_1
X_5221_ _5221_/A _5221_/B _5221_/C vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__or3_1
XFILLER_111_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5152_ _5092_/X _5151_/X _5131_/X vssd1 vssd1 vccd1 vccd1 _5152_/X sky130_fd_sc_hd__a21o_1
X_4103_ _4103_/A vssd1 vssd1 vccd1 vccd1 _8408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5083_ _5258_/A vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4034_ _8488_/Q vssd1 vssd1 vccd1 vccd1 _4298_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5985_ _5985_/A vssd1 vssd1 vccd1 vccd1 _5985_/X sky130_fd_sc_hd__clkbuf_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7115__546 _7118__549/A vssd1 vssd1 vccd1 vccd1 _8273_/CLK sky130_fd_sc_hd__inv_2
X_7724_ _5930_/A _7710_/X _7723_/X vssd1 vssd1 vccd1 vccd1 _7724_/X sky130_fd_sc_hd__a21bo_1
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4936_ _5014_/C _4943_/A _5014_/B vssd1 vssd1 vccd1 vccd1 _4937_/C sky130_fd_sc_hd__a21o_1
X_4867_ _7823_/Q _4791_/X _4809_/A _4866_/X vssd1 vssd1 vccd1 vccd1 _4867_/X sky130_fd_sc_hd__o22a_1
X_7586_ _7586_/A vssd1 vssd1 vccd1 vccd1 _7600_/A sky130_fd_sc_hd__clkbuf_2
X_6606_ _6621_/B vssd1 vssd1 vccd1 vccd1 _8167_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4798_ _4811_/A _7953_/Q _7766_/Q _4797_/X _4733_/A vssd1 vssd1 vccd1 vccd1 _4798_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3249_ clkbuf_0__3249_/X vssd1 vssd1 vccd1 vccd1 _6557__250/A sky130_fd_sc_hd__clkbuf_4
X_6468_ _5975_/A _7877_/Q _6476_/S vssd1 vssd1 vccd1 vccd1 _6469_/A sky130_fd_sc_hd__mux2_1
Xoutput150 _5947_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[20] sky130_fd_sc_hd__buf_2
Xoutput161 _5968_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[30] sky130_fd_sc_hd__buf_2
X_8207_ _8207_/CLK _8207_/D vssd1 vssd1 vccd1 vccd1 _8207_/Q sky130_fd_sc_hd__dfxtp_1
X_6399_ _6396_/X _6397_/X _6398_/Y _8545_/Q vssd1 vssd1 vccd1 vccd1 _6399_/X sky130_fd_sc_hd__a22o_1
X_5419_ _5419_/A vssd1 vssd1 vccd1 vccd1 _8086_/D sky130_fd_sc_hd__clkbuf_1
Xoutput172 _5895_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[2] sky130_fd_sc_hd__buf_2
XFILLER_114_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8138_ _8138_/CLK _8138_/D vssd1 vssd1 vccd1 vccd1 _8138_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput194 _6137_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput183 _6103_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_87_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8069_ _8069_/CLK _8069_/D vssd1 vssd1 vccd1 vccd1 _8069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3465_ clkbuf_0__3465_/X vssd1 vssd1 vccd1 vccd1 _7127__55/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7016__466 _7020__470/A vssd1 vssd1 vccd1 vccd1 _8193_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5770_ _5785_/S vssd1 vssd1 vccd1 vccd1 _5779_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6895__390 _6895__390/A vssd1 vssd1 vccd1 vccd1 _8104_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4721_ _4953_/B _4717_/X _4720_/X vssd1 vssd1 vccd1 vccd1 _4721_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4652_ _4732_/A vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__clkbuf_2
Xinput30 caravel_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4583_ _3981_/X _8205_/Q _4583_/S vssd1 vssd1 vccd1 vccd1 _4584_/A sky130_fd_sc_hd__mux2_1
Xinput52 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _3869_/A sky130_fd_sc_hd__clkbuf_1
Xinput41 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 _6000_/A sky130_fd_sc_hd__buf_4
Xinput63 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _5980_/A sky130_fd_sc_hd__buf_4
X_7371_ _7385_/S vssd1 vssd1 vccd1 vccd1 _7371_/X sky130_fd_sc_hd__clkbuf_2
X_6322_ _6322_/A vssd1 vssd1 vccd1 vccd1 _6322_/X sky130_fd_sc_hd__buf_1
Xinput96 wbs_data_i[4] vssd1 vssd1 vccd1 vccd1 _7640_/A sky130_fd_sc_hd__clkbuf_8
Xinput74 wbs_data_i[13] vssd1 vssd1 vccd1 vccd1 _5930_/A sky130_fd_sc_hd__clkbuf_2
Xinput85 wbs_data_i[23] vssd1 vssd1 vccd1 vccd1 _5952_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6253_ _6253_/A vssd1 vssd1 vccd1 vccd1 _7812_/D sky130_fd_sc_hd__clkbuf_1
X_5204_ _8304_/Q _8296_/Q _8288_/Q _8312_/Q _5095_/X _5088_/X vssd1 vssd1 vccd1 vccd1
+ _5204_/X sky130_fd_sc_hd__mux4_1
X_6184_ _6184_/A vssd1 vssd1 vccd1 vccd1 _6184_/X sky130_fd_sc_hd__buf_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5135_ _8131_/Q _5040_/X _5348_/A _5134_/X _5107_/X vssd1 vssd1 vccd1 vccd1 _5135_/X
+ sky130_fd_sc_hd__a221o_1
X_5066_ _5252_/S vssd1 vssd1 vccd1 vccd1 _5066_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4017_ _4017_/A vssd1 vssd1 vccd1 vccd1 _8440_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3250_ clkbuf_0__3250_/X vssd1 vssd1 vccd1 vccd1 _6583_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5968_ _5968_/A vssd1 vssd1 vccd1 vccd1 _5968_/X sky130_fd_sc_hd__clkbuf_1
X_4919_ _4949_/B _4908_/Y _4911_/Y _4918_/X vssd1 vssd1 vccd1 vccd1 _4920_/B sky130_fd_sc_hd__a31o_1
X_7707_ _8532_/Q _7701_/X _7706_/X _7704_/X vssd1 vssd1 vccd1 vccd1 _8532_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5899_ _5956_/A vssd1 vssd1 vccd1 vccd1 _5969_/B sky130_fd_sc_hd__buf_8
X_7638_ _7638_/A vssd1 vssd1 vccd1 vccd1 _8491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7569_ _8467_/Q vssd1 vssd1 vccd1 vccd1 _7569_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7057__500 _7057__500/A vssd1 vssd1 vccd1 vccd1 _8227_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3448_ clkbuf_0__3448_/X vssd1 vssd1 vccd1 vccd1 _7045__490/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3463_ clkbuf_0__3463_/X vssd1 vssd1 vccd1 vccd1 _7432_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6775__361 _6777__363/A vssd1 vssd1 vccd1 vccd1 _8074_/CLK sky130_fd_sc_hd__inv_2
X_7168__88 _7169__89/A vssd1 vssd1 vccd1 vccd1 _8315_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6940_ _6462_/A _7680_/B _6336_/X _7640_/C _7747_/A vssd1 vssd1 vccd1 vccd1 _8133_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_93_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3652_ clkbuf_0__3652_/X vssd1 vssd1 vccd1 vccd1 _7466__2/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6871_ _6871_/A vssd1 vssd1 vccd1 vccd1 _6871_/X sky130_fd_sc_hd__buf_1
X_5822_ _5822_/A vssd1 vssd1 vccd1 vccd1 _7830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8541_ _8543_/CLK _8541_/D vssd1 vssd1 vccd1 vccd1 _8541_/Q sky130_fd_sc_hd__dfxtp_1
X_5753_ _7909_/Q _5554_/A _5761_/S vssd1 vssd1 vccd1 vccd1 _5754_/A sky130_fd_sc_hd__mux2_1
X_4704_ _7769_/Q _7777_/Q _7852_/Q _7956_/Q _4666_/X _4667_/X vssd1 vssd1 vccd1 vccd1
+ _4704_/X sky130_fd_sc_hd__mux4_2
X_5684_ _5684_/A vssd1 vssd1 vccd1 vccd1 _7940_/D sky130_fd_sc_hd__clkbuf_1
X_8472_ _8473_/CLK _8472_/D vssd1 vssd1 vccd1 vccd1 _8472_/Q sky130_fd_sc_hd__dfxtp_1
X_4635_ _8171_/Q _4651_/A vssd1 vssd1 vccd1 vccd1 _4636_/A sky130_fd_sc_hd__and2_1
XFILLER_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4566_ _4566_/A vssd1 vssd1 vccd1 vccd1 _8213_/D sky130_fd_sc_hd__clkbuf_1
X_6533__230 _6533__230/A vssd1 vssd1 vccd1 vccd1 _7908_/CLK sky130_fd_sc_hd__inv_2
X_7354_ _7354_/A _7361_/A vssd1 vssd1 vccd1 vccd1 _7354_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4497_ _4497_/A vssd1 vssd1 vccd1 vccd1 _8242_/D sky130_fd_sc_hd__clkbuf_1
X_7285_ _7359_/A _7285_/B vssd1 vssd1 vccd1 vccd1 _7285_/X sky130_fd_sc_hd__or2_1
X_6236_ _6272_/A vssd1 vssd1 vccd1 vccd1 _6236_/X sky130_fd_sc_hd__clkbuf_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5252_/S vssd1 vssd1 vccd1 vccd1 _5290_/S sky130_fd_sc_hd__buf_2
XFILLER_85_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _7793_/Q _6105_/B vssd1 vssd1 vccd1 vccd1 _6098_/X sky130_fd_sc_hd__or2_1
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5049_ _8114_/Q vssd1 vssd1 vccd1 vccd1 _5182_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7456__170 _7456__170/A vssd1 vssd1 vccd1 vccd1 _8427_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4420_ _5602_/A _5841_/A vssd1 vssd1 vccd1 vccd1 _4445_/S sky130_fd_sc_hd__or2_2
XFILLER_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4351_ _4351_/A vssd1 vssd1 vccd1 vccd1 _8295_/D sky130_fd_sc_hd__clkbuf_1
X_7029__476 _7030__477/A vssd1 vssd1 vccd1 vccd1 _8203_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4282_ _4282_/A vssd1 vssd1 vccd1 vccd1 _8323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _6021_/A vssd1 vssd1 vccd1 vccd1 _6030_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7972_ _8520_/CLK _7972_/D vssd1 vssd1 vccd1 vccd1 _7972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6854_ _6854_/A _7514_/B vssd1 vssd1 vccd1 vccd1 _6855_/D sky130_fd_sc_hd__xor2_1
XFILLER_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3997_ _3997_/A vssd1 vssd1 vccd1 vccd1 _8446_/D sky130_fd_sc_hd__clkbuf_1
X_5805_ _5805_/A _5805_/B vssd1 vssd1 vccd1 vccd1 _5821_/S sky130_fd_sc_hd__or2_2
XFILLER_50_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6785_ _7586_/A vssd1 vssd1 vccd1 vccd1 _7568_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8524_ _8530_/CLK _8524_/D vssd1 vssd1 vccd1 vccd1 _8524_/Q sky130_fd_sc_hd__dfxtp_1
X_5736_ _5736_/A vssd1 vssd1 vccd1 vccd1 _7917_/D sky130_fd_sc_hd__clkbuf_1
X_5667_ _5608_/X _7947_/Q _5671_/S vssd1 vssd1 vccd1 vccd1 _5668_/A sky130_fd_sc_hd__mux2_1
X_8455_ _8455_/CLK _8455_/D vssd1 vssd1 vccd1 vccd1 _8455_/Q sky130_fd_sc_hd__dfxtp_1
X_4618_ _8190_/Q _4193_/X _4620_/S vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__mux2_1
X_8386_ _8386_/CLK _8386_/D vssd1 vssd1 vccd1 vccd1 _8386_/Q sky130_fd_sc_hd__dfxtp_1
X_5598_ _5598_/A vssd1 vssd1 vccd1 vccd1 _7983_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3465_ _7122_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3465_/X sky130_fd_sc_hd__clkbuf_16
X_7399__124 _7399__124/A vssd1 vssd1 vccd1 vccd1 _8381_/CLK sky130_fd_sc_hd__inv_2
X_4549_ _5823_/A _4959_/A vssd1 vssd1 vccd1 vccd1 _4565_/S sky130_fd_sc_hd__or2_2
X_7337_ _7360_/B vssd1 vssd1 vccd1 vccd1 _7348_/A sky130_fd_sc_hd__buf_2
X_7268_ _7355_/A _7303_/A vssd1 vssd1 vccd1 vccd1 _7269_/C sky130_fd_sc_hd__nand2_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7295__111 _7388__115/A vssd1 vssd1 vccd1 vccd1 _8340_/CLK sky130_fd_sc_hd__inv_2
X_6219_ _6272_/A vssd1 vssd1 vccd1 vccd1 _6219_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_10 _6272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7199_ _7199_/A vssd1 vssd1 vccd1 vccd1 _7344_/A sky130_fd_sc_hd__dlymetal6s2s_1
XINSDIODE2_43 _6131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_32 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_21 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_54 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_76 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_65 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_87 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_98 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3920_ _3920_/A vssd1 vssd1 vccd1 vccd1 _8511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3851_ _4057_/B _5070_/A vssd1 vssd1 vccd1 vccd1 _3853_/A sky130_fd_sc_hd__and2b_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5521_ _5521_/A vssd1 vssd1 vccd1 vccd1 _8037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8240_ _8240_/CLK _8240_/D vssd1 vssd1 vccd1 vccd1 _8240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5452_ _8070_/Q _4181_/X _5456_/S vssd1 vssd1 vccd1 vccd1 _5453_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3250_ _6558_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3250_/X sky130_fd_sc_hd__clkbuf_16
X_5383_ _5572_/A vssd1 vssd1 vccd1 vccd1 _5383_/X sky130_fd_sc_hd__buf_2
X_4403_ _4403_/A vssd1 vssd1 vccd1 vccd1 _8276_/D sky130_fd_sc_hd__clkbuf_1
X_8171_ _8171_/CLK _8171_/D vssd1 vssd1 vccd1 vccd1 _8171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4334_ _4295_/X _8302_/Q _4336_/S vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__mux2_1
X_7122_ _7122_/A vssd1 vssd1 vccd1 vccd1 _7122_/X sky130_fd_sc_hd__buf_1
XFILLER_113_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6004_ _8005_/Q _6008_/B vssd1 vssd1 vccd1 vccd1 _6005_/A sky130_fd_sc_hd__and2_1
X_4265_ _8329_/Q _4184_/X _4267_/S vssd1 vssd1 vccd1 vccd1 _4266_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4196_ _8488_/Q vssd1 vssd1 vccd1 vccd1 _4196_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7955_ _7955_/CLK _7955_/D vssd1 vssd1 vccd1 vccd1 _7955_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7886_ _8551_/CLK _7886_/D vssd1 vssd1 vccd1 vccd1 _7886_/Q sky130_fd_sc_hd__dfxtp_1
X_6906_ _6906_/A vssd1 vssd1 vccd1 vccd1 _8109_/D sky130_fd_sc_hd__clkbuf_1
X_6837_ _7550_/A _8461_/Q _8463_/Q vssd1 vssd1 vccd1 vccd1 _7556_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6768_ _6780_/A vssd1 vssd1 vccd1 vccd1 _6768_/X sky130_fd_sc_hd__buf_1
X_8507_ _8507_/CLK _8507_/D vssd1 vssd1 vccd1 vccd1 _8507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5719_ _7924_/Q _5583_/X _5725_/S vssd1 vssd1 vccd1 vccd1 _5720_/A sky130_fd_sc_hd__mux2_1
X_6699_ _6699_/A vssd1 vssd1 vccd1 vccd1 _8017_/D sky130_fd_sc_hd__clkbuf_1
X_8438_ _8438_/CLK _8438_/D vssd1 vssd1 vccd1 vccd1 _8438_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3448_ _7040_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3448_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8369_ _8370_/CLK _8369_/D vssd1 vssd1 vccd1 vccd1 _8369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _4050_/A vssd1 vssd1 vccd1 vccd1 _8430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 caravel_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7740_ _6854_/A _7717_/A _7739_/X _7737_/X vssd1 vssd1 vccd1 vccd1 _8543_/D sky130_fd_sc_hd__o211a_1
X_4952_ _8171_/Q _4947_/X _4951_/Y _4924_/X vssd1 vssd1 vccd1 vccd1 _8171_/D sky130_fd_sc_hd__o211a_1
XFILLER_45_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3903_ _3902_/X _8515_/Q _3903_/S vssd1 vssd1 vccd1 vccd1 _3904_/A sky130_fd_sc_hd__mux2_1
X_4883_ _7919_/Q _8023_/Q _4883_/S vssd1 vssd1 vccd1 vccd1 _4883_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6622_ _6622_/A vssd1 vssd1 vccd1 vccd1 _7973_/D sky130_fd_sc_hd__clkbuf_1
X_3834_ _8122_/Q vssd1 vssd1 vccd1 vccd1 _4057_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5504_ _8044_/Q _4280_/A _5510_/S vssd1 vssd1 vccd1 vccd1 _5505_/A sky130_fd_sc_hd__mux2_1
X_6484_ _6484_/A vssd1 vssd1 vccd1 vccd1 _7884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5435_ _5435_/A vssd1 vssd1 vccd1 vccd1 _8078_/D sky130_fd_sc_hd__clkbuf_1
X_8223_ _8223_/CLK _8223_/D vssd1 vssd1 vccd1 vccd1 _8223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5366_ _8112_/Q vssd1 vssd1 vccd1 vccd1 _5559_/A sky130_fd_sc_hd__clkbuf_4
X_8154_ _8154_/CLK _8154_/D vssd1 vssd1 vccd1 vccd1 _8154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4317_ _4317_/A vssd1 vssd1 vccd1 vccd1 _8310_/D sky130_fd_sc_hd__clkbuf_1
X_8085_ _8085_/CLK _8085_/D vssd1 vssd1 vccd1 vccd1 _8085_/Q sky130_fd_sc_hd__dfxtp_1
X_5297_ _3908_/X _5038_/A _5296_/X _5262_/X vssd1 vssd1 vccd1 vccd1 _8126_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4248_ _8338_/Q _4160_/X _4248_/S vssd1 vssd1 vccd1 vccd1 _4249_/A sky130_fd_sc_hd__mux2_1
X_6723__325 _6723__325/A vssd1 vssd1 vccd1 vccd1 _8035_/CLK sky130_fd_sc_hd__inv_2
X_4179_ _8393_/Q _4178_/X _4188_/S vssd1 vssd1 vccd1 vccd1 _4180_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7938_ _7938_/CLK _7938_/D vssd1 vssd1 vccd1 vccd1 _7938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7869_ _8537_/CLK _7869_/D vssd1 vssd1 vccd1 vccd1 _7869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6175__183 _6175__183/A vssd1 vssd1 vccd1 vccd1 _7770_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6624__289 _6625__290/A vssd1 vssd1 vccd1 vccd1 _7975_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3411_ clkbuf_0__3411_/X vssd1 vssd1 vccd1 vccd1 _6918__395/A sky130_fd_sc_hd__clkbuf_16
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220_ _5244_/A _5218_/X _5219_/X vssd1 vssd1 vccd1 vccd1 _5221_/C sky130_fd_sc_hd__o21a_1
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5151_ _8210_/Q _8194_/Q _8456_/Q _8226_/Q _5231_/S _5129_/X vssd1 vssd1 vccd1 vccd1
+ _5151_/X sky130_fd_sc_hd__mux4_2
X_4102_ _4015_/X _8408_/Q _4106_/S vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__mux2_1
X_5082_ _5103_/B _5082_/B vssd1 vssd1 vccd1 vccd1 _5258_/A sky130_fd_sc_hd__nor2_1
X_4033_ _4033_/A vssd1 vssd1 vccd1 vccd1 _8436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5984_ _5984_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _5985_/A sky130_fd_sc_hd__and2_1
X_7723_ _7728_/C vssd1 vssd1 vccd1 vccd1 _7723_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4935_ _5014_/A _4924_/X _4937_/B _4934_/Y vssd1 vssd1 vccd1 vccd1 _8177_/D sky130_fd_sc_hd__a31o_1
X_4866_ _7959_/Q _7943_/Q _4866_/S vssd1 vssd1 vccd1 vccd1 _4866_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4797_ _4797_/A vssd1 vssd1 vccd1 vccd1 _4797_/X sky130_fd_sc_hd__clkbuf_2
X_7585_ _7585_/A _7585_/B vssd1 vssd1 vccd1 vccd1 _8471_/D sky130_fd_sc_hd__nor2_1
X_6605_ _7726_/A _6605_/B vssd1 vssd1 vccd1 vccd1 _6621_/B sky130_fd_sc_hd__nor2_1
XFILLER_118_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3248_ clkbuf_0__3248_/X vssd1 vssd1 vccd1 vccd1 _6549__243/A sky130_fd_sc_hd__clkbuf_4
X_6467_ _6511_/A vssd1 vssd1 vccd1 vccd1 _6476_/S sky130_fd_sc_hd__clkbuf_2
Xoutput151 _5949_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[21] sky130_fd_sc_hd__buf_2
Xoutput140 _5927_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[11] sky130_fd_sc_hd__buf_2
X_8206_ _8206_/CLK _8206_/D vssd1 vssd1 vccd1 vccd1 _8206_/Q sky130_fd_sc_hd__dfxtp_1
X_6398_ _6398_/A _6398_/B vssd1 vssd1 vccd1 vccd1 _6398_/Y sky130_fd_sc_hd__nor2_1
X_5418_ _5399_/X _8086_/Q _5420_/S vssd1 vssd1 vccd1 vccd1 _5419_/A sky130_fd_sc_hd__mux2_1
Xoutput173 _5897_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[3] sky130_fd_sc_hd__buf_2
Xoutput162 _5970_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[31] sky130_fd_sc_hd__buf_2
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8137_ _8137_/CLK _8137_/D vssd1 vssd1 vccd1 vccd1 _8137_/Q sky130_fd_sc_hd__dfxtp_1
X_5349_ _5349_/A vssd1 vssd1 vccd1 vccd1 _5356_/A sky130_fd_sc_hd__clkbuf_2
Xoutput195 _6141_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[26] sky130_fd_sc_hd__buf_2
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput184 _6106_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_114_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8068_ _8068_/CLK _8068_/D vssd1 vssd1 vccd1 vccd1 _8068_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3464_ clkbuf_0__3464_/X vssd1 vssd1 vccd1 vccd1 _7146_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6582__270 _6582__270/A vssd1 vssd1 vccd1 vccd1 _7948_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7450__165 _7450__165/A vssd1 vssd1 vccd1 vccd1 _8422_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4664_/X _4719_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__a21o_1
X_4651_ _4651_/A _4783_/A vssd1 vssd1 vccd1 vccd1 _4732_/A sky130_fd_sc_hd__nor2_1
Xinput20 caravel_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 _6135_/A sky130_fd_sc_hd__clkbuf_4
Xinput31 caravel_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
X_4582_ _4582_/A vssd1 vssd1 vccd1 vccd1 _8206_/D sky130_fd_sc_hd__clkbuf_1
Xinput53 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _3869_/D sky130_fd_sc_hd__clkbuf_1
Xinput64 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _5982_/A sky130_fd_sc_hd__buf_4
Xinput42 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 _6002_/A sky130_fd_sc_hd__buf_4
X_7370_ _8363_/Q _7377_/B vssd1 vssd1 vccd1 vccd1 _7370_/X sky130_fd_sc_hd__or2_1
Xinput86 wbs_data_i[24] vssd1 vssd1 vccd1 vccd1 _5954_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput97 wbs_data_i[5] vssd1 vssd1 vccd1 vccd1 _7642_/A sky130_fd_sc_hd__buf_4
Xinput75 wbs_data_i[14] vssd1 vssd1 vccd1 vccd1 _5932_/A sky130_fd_sc_hd__clkbuf_2
X_6252_ _7633_/B _7812_/Q _6258_/S vssd1 vssd1 vccd1 vccd1 _6253_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5203_ _8422_/Q _8320_/Q _8057_/Q _8272_/Q _5080_/A _5308_/S vssd1 vssd1 vccd1 vccd1
+ _5203_/X sky130_fd_sc_hd__mux4_1
X_8562__209 vssd1 vssd1 vccd1 vccd1 _8562__209/HI caravel_irq[0] sky130_fd_sc_hd__conb_1
X_7393__119 _7394__120/A vssd1 vssd1 vccd1 vccd1 _8376_/CLK sky130_fd_sc_hd__inv_2
X_5134_ _5047_/X _5116_/X _5121_/X _5133_/X vssd1 vssd1 vccd1 vccd1 _5134_/X sky130_fd_sc_hd__a31o_2
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5065_ _5250_/A vssd1 vssd1 vccd1 vccd1 _5354_/B sky130_fd_sc_hd__clkbuf_4
X_4016_ _4015_/X _8440_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4017_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7468__4 _7469__5/A vssd1 vssd1 vccd1 vccd1 _8436_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5967_ _5967_/A _5969_/B vssd1 vssd1 vccd1 vccd1 _5968_/A sky130_fd_sc_hd__or2_1
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4918_ _4638_/A _4914_/Y _4917_/Y _4951_/B vssd1 vssd1 vccd1 vccd1 _4918_/X sky130_fd_sc_hd__a31o_1
X_7706_ _5943_/A _7702_/X _7701_/A vssd1 vssd1 vccd1 vccd1 _7706_/X sky130_fd_sc_hd__a21bo_1
XFILLER_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5898_ _5898_/A vssd1 vssd1 vccd1 vccd1 _5956_/A sky130_fd_sc_hd__buf_6
X_7637_ _7637_/A _7637_/B _7640_/C vssd1 vssd1 vccd1 vccd1 _7638_/A sky130_fd_sc_hd__and3_1
X_4849_ _4803_/A _4847_/X _4848_/X vssd1 vssd1 vccd1 vccd1 _4853_/B sky130_fd_sc_hd__o21a_1
XFILLER_107_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7568_ _7568_/A vssd1 vssd1 vccd1 vccd1 _7585_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7499_ _7502_/A input1/X vssd1 vssd1 vccd1 vccd1 _7499_/X sky130_fd_sc_hd__or2_1
X_6519_ _7689_/A _6519_/B vssd1 vssd1 vccd1 vccd1 _6522_/B sky130_fd_sc_hd__and2_1
XFILLER_88_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7022__471 _7023__472/A vssd1 vssd1 vccd1 vccd1 _8198_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3447_ clkbuf_0__3447_/X vssd1 vssd1 vccd1 vccd1 _7039__485/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6736__335 _6736__335/A vssd1 vssd1 vccd1 vccd1 _8045_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7064__505 _7064__505/A vssd1 vssd1 vccd1 vccd1 _8232_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3651_ clkbuf_0__3651_/X vssd1 vssd1 vccd1 vccd1 _7488_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5821_ _3981_/X _7830_/Q _5821_/S vssd1 vssd1 vccd1 vccd1 _5822_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5752_ _5767_/S vssd1 vssd1 vccd1 vccd1 _5761_/S sky130_fd_sc_hd__clkbuf_2
X_8540_ _8540_/CLK _8540_/D vssd1 vssd1 vccd1 vccd1 _8540_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4703_ _4701_/X _4702_/X _4760_/S vssd1 vssd1 vccd1 vccd1 _4703_/X sky130_fd_sc_hd__mux2_1
X_5683_ _7940_/Q _5583_/X _5689_/S vssd1 vssd1 vccd1 vccd1 _5684_/A sky130_fd_sc_hd__mux2_1
X_8471_ _8473_/CLK _8471_/D vssd1 vssd1 vccd1 vccd1 _8471_/Q sky130_fd_sc_hd__dfxtp_1
X_4634_ _8170_/Q _4767_/A _8168_/Q vssd1 vssd1 vccd1 vccd1 _4651_/A sky130_fd_sc_hd__and3_1
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4565_ _4444_/X _8213_/Q _4565_/S vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__mux2_1
X_7353_ _7354_/A _7361_/A _7352_/X _7286_/X vssd1 vssd1 vccd1 vccd1 _8359_/D sky130_fd_sc_hd__o211a_1
X_6304_ _6310_/A vssd1 vssd1 vccd1 vccd1 _6304_/X sky130_fd_sc_hd__buf_1
XFILLER_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4496_ _4382_/X _8242_/Q _4500_/S vssd1 vssd1 vccd1 vccd1 _4497_/A sky130_fd_sc_hd__mux2_1
X_7284_ _8333_/Q _7284_/B _7284_/C _7284_/D vssd1 vssd1 vccd1 vccd1 _7285_/B sky130_fd_sc_hd__and4_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6235_ _6235_/A vssd1 vssd1 vccd1 vccd1 _7680_/A sky130_fd_sc_hd__buf_6
X_6166_ _6291_/A vssd1 vssd1 vccd1 vccd1 _6166_/X sky130_fd_sc_hd__buf_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5117_ _7844_/Q _8052_/Q _8331_/Q _8079_/Q _5273_/S _5068_/X vssd1 vssd1 vccd1 vccd1
+ _5117_/X sky130_fd_sc_hd__mux4_2
XFILLER_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _7868_/Q input8/X _6111_/S vssd1 vssd1 vccd1 vccd1 _6097_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5048_ _8115_/Q vssd1 vssd1 vccd1 vccd1 _5181_/A sky130_fd_sc_hd__buf_2
XFILLER_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7173__92 _7173__92/A vssd1 vssd1 vccd1 vccd1 _8319_/CLK sky130_fd_sc_hd__inv_2
X_8584__231 vssd1 vssd1 vccd1 vccd1 _8584__231/HI manufacturerID[3] sky130_fd_sc_hd__conb_1
XFILLER_4_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6595__280 _6595__280/A vssd1 vssd1 vccd1 vccd1 _7958_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4350_ _4292_/X _8295_/Q _4354_/S vssd1 vssd1 vccd1 vccd1 _4351_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4281_ _4280_/X _8323_/Q _4290_/S vssd1 vssd1 vccd1 vccd1 _4282_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6020_ _6020_/A vssd1 vssd1 vccd1 vccd1 _6020_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7971_ _8520_/CLK _7971_/D vssd1 vssd1 vccd1 vccd1 _7971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6853_ _6853_/A _6853_/B vssd1 vssd1 vccd1 vccd1 _7514_/B sky130_fd_sc_hd__xnor2_2
X_6936__409 _6936__409/A vssd1 vssd1 vccd1 vccd1 _8131_/CLK sky130_fd_sc_hd__inv_2
X_6604__287 _6604__287/A vssd1 vssd1 vccd1 vccd1 _7965_/CLK sky130_fd_sc_hd__inv_2
X_5804_ _5804_/A vssd1 vssd1 vccd1 vccd1 _7838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3996_ _3902_/X _8446_/Q _3996_/S vssd1 vssd1 vccd1 vccd1 _3997_/A sky130_fd_sc_hd__mux2_1
X_6784_ _7552_/A vssd1 vssd1 vccd1 vccd1 _7586_/A sky130_fd_sc_hd__inv_2
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8523_ _8530_/CLK _8523_/D vssd1 vssd1 vccd1 vccd1 _8523_/Q sky130_fd_sc_hd__dfxtp_1
X_5735_ _7917_/Q _5554_/A _5743_/S vssd1 vssd1 vccd1 vccd1 _5736_/A sky130_fd_sc_hd__mux2_1
X_5666_ _5666_/A vssd1 vssd1 vccd1 vccd1 _7948_/D sky130_fd_sc_hd__clkbuf_1
X_8454_ _8454_/CLK _8454_/D vssd1 vssd1 vccd1 vccd1 _8454_/Q sky130_fd_sc_hd__dfxtp_1
X_4617_ _4617_/A vssd1 vssd1 vccd1 vccd1 _8191_/D sky130_fd_sc_hd__clkbuf_1
X_8568__215 vssd1 vssd1 vccd1 vccd1 _8568__215/HI core0Index[2] sky130_fd_sc_hd__conb_1
X_8385_ _8385_/CLK _8385_/D vssd1 vssd1 vccd1 vccd1 _8385_/Q sky130_fd_sc_hd__dfxtp_1
X_5597_ _7983_/Q _5596_/X _5600_/S vssd1 vssd1 vccd1 vccd1 _5598_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3464_ _7121_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3464_/X sky130_fd_sc_hd__clkbuf_16
X_4548_ _4548_/A vssd1 vssd1 vccd1 vccd1 _8221_/D sky130_fd_sc_hd__clkbuf_1
X_7336_ _7336_/A _7336_/B vssd1 vssd1 vccd1 vccd1 _8353_/D sky130_fd_sc_hd__nor2_1
XFILLER_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4479_ _8248_/Q _4478_/X _4479_/S vssd1 vssd1 vccd1 vccd1 _4480_/A sky130_fd_sc_hd__mux2_1
X_7267_ _7350_/B _7303_/A _7383_/B _7355_/A vssd1 vssd1 vccd1 vccd1 _7269_/B sky130_fd_sc_hd__a211o_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6218_ _6217_/X _8003_/Q _6211_/X _6213_/X _7792_/Q vssd1 vssd1 vccd1 vccd1 _7792_/D
+ sky130_fd_sc_hd__o32a_1
X_7198_ _8357_/Q _8356_/Q _7257_/A vssd1 vssd1 vccd1 vccd1 _7199_/A sky130_fd_sc_hd__nand3_1
XINSDIODE2_22 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_11 _7552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_33 _6123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6149_ _6149_/A _6151_/B vssd1 vssd1 vccd1 vccd1 _6149_/X sky130_fd_sc_hd__and2_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_44 _6131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_77 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_66 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_55 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_88 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_99 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3850_ _8117_/Q vssd1 vssd1 vccd1 vccd1 _5070_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7035__481 _7039__485/A vssd1 vssd1 vccd1 vccd1 _8208_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5520_ _5361_/X _8037_/Q _5528_/S vssd1 vssd1 vccd1 vccd1 _5521_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5451_ _5451_/A vssd1 vssd1 vccd1 vccd1 _8071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5382_ _8107_/Q vssd1 vssd1 vccd1 vccd1 _5572_/A sky130_fd_sc_hd__clkbuf_2
X_4402_ _4374_/X _8276_/Q _4410_/S vssd1 vssd1 vccd1 vccd1 _4403_/A sky130_fd_sc_hd__mux2_1
X_8170_ _8170_/CLK _8170_/D vssd1 vssd1 vccd1 vccd1 _8170_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4333_ _4333_/A vssd1 vssd1 vccd1 vccd1 _8303_/D sky130_fd_sc_hd__clkbuf_1
X_7121_ _7152_/A vssd1 vssd1 vccd1 vccd1 _7121_/X sky130_fd_sc_hd__buf_1
XFILLER_115_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4264_ _4264_/A vssd1 vssd1 vccd1 vccd1 _8330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7052_ _7052_/A vssd1 vssd1 vccd1 vccd1 _7052_/X sky130_fd_sc_hd__buf_1
X_6003_ _6003_/A vssd1 vssd1 vccd1 vccd1 _6003_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4195_ _4195_/A vssd1 vssd1 vccd1 vccd1 _8388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7003__458 _7005__460/A vssd1 vssd1 vccd1 vccd1 _8183_/CLK sky130_fd_sc_hd__inv_2
X_7954_ _7954_/CLK _7954_/D vssd1 vssd1 vccd1 vccd1 _7954_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ _8483_/Q _6911_/B vssd1 vssd1 vccd1 vccd1 _6906_/A sky130_fd_sc_hd__and2_1
X_7885_ _8551_/CLK _7885_/D vssd1 vssd1 vccd1 vccd1 _7885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6836_ _7518_/B vssd1 vssd1 vccd1 vccd1 _7556_/A sky130_fd_sc_hd__clkbuf_2
X_3979_ _8452_/Q _3978_/X _3982_/S vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__mux2_1
X_8506_ _8506_/CLK _8506_/D vssd1 vssd1 vccd1 vccd1 _8506_/Q sky130_fd_sc_hd__dfxtp_1
X_5718_ _5718_/A vssd1 vssd1 vccd1 vccd1 _7925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6698_ _8017_/Q _5961_/A _6700_/S vssd1 vssd1 vccd1 vccd1 _6699_/A sky130_fd_sc_hd__mux2_1
X_5649_ _5649_/A vssd1 vssd1 vccd1 vccd1 _7955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8437_ _8437_/CLK _8437_/D vssd1 vssd1 vccd1 vccd1 _8437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3447_ _7034_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3447_/X sky130_fd_sc_hd__clkbuf_16
X_8368_ _8368_/CLK _8368_/D vssd1 vssd1 vccd1 vccd1 _8368_/Q sky130_fd_sc_hd__dfxtp_1
X_7319_ _7319_/A _7319_/B vssd1 vssd1 vccd1 vccd1 _7319_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8299_ _8299_/CLK _8299_/D vssd1 vssd1 vccd1 vccd1 _8299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 caravel_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ _4955_/A _4951_/B vssd1 vssd1 vccd1 vccd1 _4951_/Y sky130_fd_sc_hd__nand2_1
X_7670_ _7670_/A vssd1 vssd1 vccd1 vccd1 _7670_/X sky130_fd_sc_hd__buf_1
X_4882_ _8091_/Q _4781_/A _4726_/A _4881_/X vssd1 vssd1 vccd1 vccd1 _4886_/B sky130_fd_sc_hd__o211a_1
X_3902_ _8491_/Q vssd1 vssd1 vccd1 vccd1 _3902_/X sky130_fd_sc_hd__buf_4
X_3833_ _4076_/A vssd1 vssd1 vccd1 vccd1 _4256_/C sky130_fd_sc_hd__buf_2
X_6621_ _8186_/Q _6621_/B vssd1 vssd1 vccd1 vccd1 _6622_/A sky130_fd_sc_hd__and2_1
XFILLER_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6552_ _6552_/A vssd1 vssd1 vccd1 vccd1 _6552_/X sky130_fd_sc_hd__buf_1
XFILLER_118_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5503_ _5503_/A vssd1 vssd1 vccd1 vccd1 _8045_/D sky130_fd_sc_hd__clkbuf_1
X_6483_ _5991_/A _7884_/Q _6487_/S vssd1 vssd1 vccd1 vccd1 _6484_/A sky130_fd_sc_hd__mux2_1
X_5434_ _3966_/X _8078_/Q _5438_/S vssd1 vssd1 vccd1 vccd1 _5435_/A sky130_fd_sc_hd__mux2_1
X_8222_ _8222_/CLK _8222_/D vssd1 vssd1 vccd1 vccd1 _8222_/Q sky130_fd_sc_hd__dfxtp_1
X_8153_ _8153_/CLK _8153_/D vssd1 vssd1 vccd1 vccd1 _8153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5365_ _5365_/A vssd1 vssd1 vccd1 vccd1 _8105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4316_ _4295_/X _8310_/Q _4318_/S vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__mux2_1
X_8084_ _8084_/CLK _8084_/D vssd1 vssd1 vccd1 vccd1 _8084_/Q sky130_fd_sc_hd__dfxtp_1
X_5296_ _8126_/Q _5041_/A _5349_/A _5295_/Y _5107_/A vssd1 vssd1 vccd1 vccd1 _5296_/X
+ sky130_fd_sc_hd__a221o_1
X_4247_ _4247_/A vssd1 vssd1 vccd1 vccd1 _8339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4178_ _8494_/Q vssd1 vssd1 vccd1 vccd1 _4178_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7937_ _7937_/CLK _7937_/D vssd1 vssd1 vccd1 vccd1 _7937_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ _8537_/CLK _7868_/D vssd1 vssd1 vccd1 vccd1 _7868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6819_ _8466_/Q _8465_/Q vssd1 vssd1 vccd1 vccd1 _6830_/B sky130_fd_sc_hd__and2_1
XFILLER_51_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7799_ _8531_/CLK _7799_/D vssd1 vssd1 vccd1 vccd1 _7799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6988__446 _6989__447/A vssd1 vssd1 vccd1 vccd1 _8171_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5150_ _5169_/A _5150_/B vssd1 vssd1 vccd1 vccd1 _5150_/X sky130_fd_sc_hd__and2_1
X_4101_ _4101_/A vssd1 vssd1 vccd1 vccd1 _8409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5081_ _8442_/Q _8434_/Q _7837_/Q _8450_/Q _5066_/X _5080_/X vssd1 vssd1 vccd1 vccd1
+ _5081_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4032_ _4031_/X _8436_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4033_/A sky130_fd_sc_hd__mux2_1
X_6642__302 _6643__303/A vssd1 vssd1 vccd1 vccd1 _7988_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5983_ _5983_/A vssd1 vssd1 vccd1 vccd1 _5983_/X sky130_fd_sc_hd__clkbuf_1
X_4934_ _5733_/A _5859_/B vssd1 vssd1 vccd1 vccd1 _4934_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7722_ _6440_/A _7717_/X _7721_/X _7719_/X vssd1 vssd1 vccd1 vccd1 _8537_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_19_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _8550_/CLK sky130_fd_sc_hd__clkbuf_16
X_4865_ _7927_/Q _4658_/B _4784_/X vssd1 vssd1 vccd1 vccd1 _4865_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4796_ _8170_/Q vssd1 vssd1 vccd1 vccd1 _4811_/A sky130_fd_sc_hd__clkbuf_2
X_7584_ _6816_/A _7570_/X _7575_/X _7525_/B vssd1 vssd1 vccd1 vccd1 _7585_/B sky130_fd_sc_hd__o22a_1
Xclkbuf_1_1_0__3247_ clkbuf_0__3247_/X vssd1 vssd1 vccd1 vccd1 _6545__240/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8205_ _8205_/CLK _8205_/D vssd1 vssd1 vccd1 vccd1 _8205_/Q sky130_fd_sc_hd__dfxtp_1
X_6466_ _6466_/A _6466_/B _6466_/C _6284_/X vssd1 vssd1 vccd1 vccd1 _6511_/A sky130_fd_sc_hd__or4b_4
Xoutput141 _5929_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[12] sky130_fd_sc_hd__buf_2
Xoutput130 _5979_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[3] sky130_fd_sc_hd__buf_2
Xoutput152 _5951_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[22] sky130_fd_sc_hd__buf_2
X_6397_ _6397_/A _6397_/B vssd1 vssd1 vccd1 vccd1 _6397_/X sky130_fd_sc_hd__and2_1
X_5417_ _5417_/A vssd1 vssd1 vccd1 vccd1 _8087_/D sky130_fd_sc_hd__clkbuf_1
Xoutput174 _5885_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_stb_o sky130_fd_sc_hd__buf_2
Xoutput163 _5909_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_114_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8136_ _8136_/CLK _8136_/D vssd1 vssd1 vccd1 vccd1 _8136_/Q sky130_fd_sc_hd__dfxtp_1
X_5348_ _5348_/A vssd1 vssd1 vccd1 vccd1 _5348_/X sky130_fd_sc_hd__clkbuf_2
Xoutput185 _6110_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8067_ _8067_/CLK _8067_/D vssd1 vssd1 vccd1 vccd1 _8067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput196 _6144_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[27] sky130_fd_sc_hd__buf_2
X_5279_ _5235_/A _5275_/Y _5278_/Y _5047_/A vssd1 vssd1 vccd1 vccd1 _5279_/X sky130_fd_sc_hd__a31o_1
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7188__104 _7189__105/A vssd1 vssd1 vccd1 vccd1 _8331_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6630__294 _6631__295/A vssd1 vssd1 vccd1 vccd1 _7980_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7655__33 _7656__34/A vssd1 vssd1 vccd1 vccd1 _8502_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _8097_/Q _8089_/Q _7917_/Q _8158_/Q _4646_/X _4649_/X vssd1 vssd1 vccd1 vccd1
+ _4650_/X sky130_fd_sc_hd__mux4_1
Xinput21 caravel_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 _6140_/A sky130_fd_sc_hd__clkbuf_4
Xinput10 caravel_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_4
X_7427__146 _7429__148/A vssd1 vssd1 vccd1 vccd1 _8403_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput32 caravel_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_4
X_4581_ _3978_/X _8206_/Q _4583_/S vssd1 vssd1 vccd1 vccd1 _4582_/A sky130_fd_sc_hd__mux2_1
Xinput54 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _3869_/C sky130_fd_sc_hd__clkbuf_1
Xinput43 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _6108_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput65 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _5984_/A sky130_fd_sc_hd__buf_4
Xinput76 wbs_data_i[15] vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__buf_4
Xinput87 wbs_data_i[25] vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__buf_4
Xinput98 wbs_data_i[6] vssd1 vssd1 vccd1 vccd1 _7644_/A sky130_fd_sc_hd__buf_4
X_6251_ _6251_/A vssd1 vssd1 vccd1 vccd1 _7811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5202_ _5354_/B _5191_/X _5200_/X _5352_/B vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__a211o_1
X_5133_ _5206_/A _5126_/X _5128_/X _5132_/X _5177_/A vssd1 vssd1 vccd1 vccd1 _5133_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5064_ _5100_/A vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4015_ _4283_/A vssd1 vssd1 vccd1 vccd1 _4015_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _5966_/A vssd1 vssd1 vccd1 vccd1 _5966_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5897_ _5897_/A vssd1 vssd1 vccd1 vccd1 _5897_/X sky130_fd_sc_hd__clkbuf_1
X_4917_ _4794_/X _4915_/X _4916_/X vssd1 vssd1 vccd1 vccd1 _4917_/Y sky130_fd_sc_hd__o21ai_1
X_7705_ _8531_/Q _7701_/X _7703_/X _7704_/X vssd1 vssd1 vccd1 vccd1 _8531_/D sky130_fd_sc_hd__o211a_1
X_4848_ _4805_/A _7904_/Q _4797_/A _8137_/Q _4732_/A vssd1 vssd1 vccd1 vccd1 _4848_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7636_ _7636_/A vssd1 vssd1 vccd1 vccd1 _8490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _4770_/X _4773_/X _4778_/X vssd1 vssd1 vccd1 vccd1 _4779_/X sky130_fd_sc_hd__o21a_1
X_7567_ _7567_/A _7567_/B vssd1 vssd1 vccd1 vccd1 _8466_/D sky130_fd_sc_hd__nor2_1
X_7498_ _8479_/Q _8478_/Q _8477_/Q vssd1 vssd1 vccd1 vccd1 _7609_/B sky130_fd_sc_hd__and3_1
X_6518_ _6465_/A _6284_/X _6161_/C _6382_/A vssd1 vssd1 vccd1 vccd1 _6519_/B sky130_fd_sc_hd__a31o_1
X_6449_ _8534_/Q vssd1 vssd1 vccd1 vccd1 _7008_/A sky130_fd_sc_hd__buf_4
X_6649__308 _6649__308/A vssd1 vssd1 vccd1 vccd1 _7994_/CLK sky130_fd_sc_hd__inv_2
X_8119_ _8119_/CLK _8119_/D vssd1 vssd1 vccd1 vccd1 _8119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3446_ clkbuf_0__3446_/X vssd1 vssd1 vccd1 vccd1 _7030__477/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6879__376 _6881__378/A vssd1 vssd1 vccd1 vccd1 _8090_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6782__367 _6782__367/A vssd1 vssd1 vccd1 vccd1 _8080_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3650_ clkbuf_0__3650_/X vssd1 vssd1 vccd1 vccd1 _7462__175/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5820_ _5820_/A vssd1 vssd1 vccd1 vccd1 _7831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5751_ _5751_/A _5751_/B vssd1 vssd1 vccd1 vccd1 _5767_/S sky130_fd_sc_hd__nor2_2
X_4702_ _8149_/Q _8104_/Q _7996_/Q _8341_/Q _4646_/A _4649_/A vssd1 vssd1 vccd1 vccd1
+ _4702_/X sky130_fd_sc_hd__mux4_1
X_8470_ _8473_/CLK _8470_/D vssd1 vssd1 vccd1 vccd1 _8470_/Q sky130_fd_sc_hd__dfxtp_1
X_5682_ _5682_/A vssd1 vssd1 vccd1 vccd1 _7941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4633_ _8169_/Q vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4564_ _4564_/A vssd1 vssd1 vccd1 vccd1 _8214_/D sky130_fd_sc_hd__clkbuf_1
X_7352_ _7359_/A _7303_/A _7350_/Y _7356_/B vssd1 vssd1 vccd1 vccd1 _7352_/X sky130_fd_sc_hd__a31o_1
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7283_ _7278_/X _7279_/Y _7280_/X _7281_/X _7282_/X vssd1 vssd1 vccd1 vccd1 _7284_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_104_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4495_ _4495_/A vssd1 vssd1 vccd1 vccd1 _8243_/D sky130_fd_sc_hd__clkbuf_1
X_6234_ _6233_/X _8013_/Q _6227_/X _6229_/X _7802_/Q vssd1 vssd1 vccd1 vccd1 _7802_/D
+ sky130_fd_sc_hd__o32a_1
X_6165_ _6297_/A vssd1 vssd1 vccd1 vccd1 _6165_/X sky130_fd_sc_hd__buf_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _5055_/X _5113_/X _5115_/X vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6114_/A vssd1 vssd1 vccd1 vccd1 _6111_/S sky130_fd_sc_hd__clkbuf_2
X_5047_ _5047_/A vssd1 vssd1 vccd1 vccd1 _5047_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5949_ _5949_/A vssd1 vssd1 vccd1 vccd1 _5949_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7619_ _8482_/Q _7614_/X vssd1 vssd1 vccd1 vccd1 _7619_/X sky130_fd_sc_hd__or2b_1
XFILLER_119_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6742__340 _6742__340/A vssd1 vssd1 vccd1 vccd1 _8050_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3429_ clkbuf_0__3429_/X vssd1 vssd1 vccd1 vccd1 _6952__418/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7070__510 _7070__510/A vssd1 vssd1 vccd1 vccd1 _8237_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4280_ _4280_/A vssd1 vssd1 vccd1 vccd1 _4280_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7970_ _8526_/CLK _7970_/D vssd1 vssd1 vccd1 vccd1 _7970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6852_ _8469_/Q vssd1 vssd1 vccd1 vccd1 _6853_/A sky130_fd_sc_hd__inv_2
XFILLER_35_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5803_ _7838_/Q _4298_/A _5803_/S vssd1 vssd1 vccd1 vccd1 _5804_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3995_ _3995_/A vssd1 vssd1 vccd1 vccd1 _8447_/D sky130_fd_sc_hd__clkbuf_1
X_6783_ _7631_/A _6465_/B _4122_/Y _6466_/A vssd1 vssd1 vccd1 vccd1 _7552_/A sky130_fd_sc_hd__a31oi_4
X_8522_ _8530_/CLK _8522_/D vssd1 vssd1 vccd1 vccd1 _8522_/Q sky130_fd_sc_hd__dfxtp_1
X_5734_ _5749_/S vssd1 vssd1 vccd1 vccd1 _5743_/S sky130_fd_sc_hd__buf_2
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5665_ _5559_/X _7948_/Q _5671_/S vssd1 vssd1 vccd1 vccd1 _5666_/A sky130_fd_sc_hd__mux2_1
X_8453_ _8453_/CLK _8453_/D vssd1 vssd1 vccd1 vccd1 _8453_/Q sky130_fd_sc_hd__dfxtp_1
X_8384_ _8384_/CLK _8384_/D vssd1 vssd1 vccd1 vccd1 _8384_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3463_ _7120_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3463_/X sky130_fd_sc_hd__clkbuf_16
X_4616_ _8191_/Q _4190_/X _4620_/S vssd1 vssd1 vccd1 vccd1 _4617_/A sky130_fd_sc_hd__mux2_1
X_5596_ _8107_/Q vssd1 vssd1 vccd1 vccd1 _5596_/X sky130_fd_sc_hd__clkbuf_2
X_7335_ _8353_/Q _7334_/X _7326_/X _7221_/B vssd1 vssd1 vccd1 vccd1 _7336_/B sky130_fd_sc_hd__o2bb2a_1
X_4547_ _4397_/X _8221_/Q _4547_/S vssd1 vssd1 vccd1 vccd1 _4548_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4478_ _8109_/Q vssd1 vssd1 vccd1 vccd1 _4478_/X sky130_fd_sc_hd__clkbuf_4
X_7266_ _7363_/A _7365_/A vssd1 vssd1 vccd1 vccd1 _7383_/B sky130_fd_sc_hd__nor2_2
X_6217_ _6235_/A vssd1 vssd1 vccd1 vccd1 _6217_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7197_ _8355_/Q _7236_/B _7232_/C _7197_/D vssd1 vssd1 vccd1 vccd1 _7257_/A sky130_fd_sc_hd__and4_2
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6148_ _7808_/Q _6138_/X _6139_/X _6147_/X _6136_/X vssd1 vssd1 vccd1 vccd1 _6148_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_12 _8539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_23 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_34 _6123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_67 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_56 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6079_ _6075_/X _6077_/X _6078_/X _6063_/X vssd1 vssd1 vccd1 vccd1 _6079_/X sky130_fd_sc_hd__o211a_1
XINSDIODE2_45 _6135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_89 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_78 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5450_ _8071_/Q _4178_/X _5456_/S vssd1 vssd1 vccd1 vccd1 _5451_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4401_ _4416_/S vssd1 vssd1 vccd1 vccd1 _4410_/S sky130_fd_sc_hd__clkbuf_2
X_5381_ _5381_/A vssd1 vssd1 vccd1 vccd1 _8100_/D sky130_fd_sc_hd__clkbuf_1
X_4332_ _4292_/X _8303_/Q _4336_/S vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__mux2_1
X_7120_ _7120_/A vssd1 vssd1 vccd1 vccd1 _7120_/X sky130_fd_sc_hd__buf_1
X_4263_ _8330_/Q _4181_/X _4267_/S vssd1 vssd1 vccd1 vccd1 _4264_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6002_ _6002_/A _6008_/B vssd1 vssd1 vccd1 vccd1 _6003_/A sky130_fd_sc_hd__and2_1
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4194_ _8388_/Q _4193_/X _4197_/S vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7953_ _7953_/CLK _7953_/D vssd1 vssd1 vccd1 vccd1 _7953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6904_ _6904_/A vssd1 vssd1 vccd1 vccd1 _8108_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7884_ _8551_/CLK _7884_/D vssd1 vssd1 vccd1 vccd1 _7884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6835_ _8463_/Q _7550_/A _8461_/Q vssd1 vssd1 vccd1 vccd1 _7518_/B sky130_fd_sc_hd__nand3_1
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3978_ _8489_/Q vssd1 vssd1 vccd1 vccd1 _3978_/X sky130_fd_sc_hd__buf_2
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8505_ _8505_/CLK _8505_/D vssd1 vssd1 vccd1 vccd1 _8505_/Q sky130_fd_sc_hd__dfxtp_1
X_5717_ _7925_/Q _5578_/X _5725_/S vssd1 vssd1 vccd1 vccd1 _5718_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6697_ _6697_/A vssd1 vssd1 vccd1 vccd1 _8016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5648_ _7955_/Q _5647_/X _5653_/S vssd1 vssd1 vccd1 vccd1 _5649_/A sky130_fd_sc_hd__mux2_1
X_8436_ _8436_/CLK _8436_/D vssd1 vssd1 vccd1 vccd1 _8436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5579_ _5679_/B _5733_/A vssd1 vssd1 vccd1 vccd1 _5600_/S sky130_fd_sc_hd__nor2_2
Xclkbuf_0__3446_ _7028_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3446_/X sky130_fd_sc_hd__clkbuf_16
X_8367_ _8368_/CLK _8367_/D vssd1 vssd1 vccd1 vccd1 _8367_/Q sky130_fd_sc_hd__dfxtp_1
X_8298_ _8298_/CLK _8298_/D vssd1 vssd1 vccd1 vccd1 _8298_/Q sky130_fd_sc_hd__dfxtp_1
X_7318_ _7334_/A vssd1 vssd1 vccd1 vccd1 _7318_/X sky130_fd_sc_hd__clkbuf_1
X_7249_ _7242_/X _7243_/Y _7246_/Y _7247_/Y _7248_/X vssd1 vssd1 vccd1 vccd1 _7281_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_77_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6553__246 _6554__247/A vssd1 vssd1 vccd1 vccd1 _7924_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 caravel_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4950_ _8172_/Q _4947_/X _4949_/Y _4857_/X vssd1 vssd1 vccd1 vccd1 _8172_/D sky130_fd_sc_hd__o211a_1
X_3901_ _3901_/A vssd1 vssd1 vccd1 vccd1 _8516_/D sky130_fd_sc_hd__clkbuf_1
X_4881_ _8152_/Q _4784_/A _4880_/X _4786_/A vssd1 vssd1 vccd1 vccd1 _4881_/X sky130_fd_sc_hd__o22a_1
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6620_ _6620_/A vssd1 vssd1 vccd1 vccd1 _7972_/D sky130_fd_sc_hd__clkbuf_1
X_3832_ _8121_/Q vssd1 vssd1 vccd1 vccd1 _4076_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5502_ _8045_/Q _4275_/A _5510_/S vssd1 vssd1 vccd1 vccd1 _5503_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6482_ _6482_/A vssd1 vssd1 vccd1 vccd1 _7883_/D sky130_fd_sc_hd__clkbuf_1
X_5433_ _5433_/A vssd1 vssd1 vccd1 vccd1 _8079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8221_ _8221_/CLK _8221_/D vssd1 vssd1 vccd1 vccd1 _8221_/Q sky130_fd_sc_hd__dfxtp_1
X_5364_ _5361_/X _8105_/Q _5376_/S vssd1 vssd1 vccd1 vccd1 _5365_/A sky130_fd_sc_hd__mux2_1
X_8152_ _8152_/CLK _8152_/D vssd1 vssd1 vccd1 vccd1 _8152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4315_ _4315_/A vssd1 vssd1 vccd1 vccd1 _8311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5295_ _5295_/A _5295_/B vssd1 vssd1 vccd1 vccd1 _5295_/Y sky130_fd_sc_hd__nand2_2
X_8083_ _8083_/CLK _8083_/D vssd1 vssd1 vccd1 vccd1 _8083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4246_ _8339_/Q _4157_/X _4248_/S vssd1 vssd1 vccd1 vccd1 _4247_/A sky130_fd_sc_hd__mux2_1
X_7034_ _7052_/A vssd1 vssd1 vccd1 vccd1 _7034_/X sky130_fd_sc_hd__buf_1
X_4177_ _4177_/A vssd1 vssd1 vccd1 vccd1 _8394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7936_ _7936_/CLK _7936_/D vssd1 vssd1 vccd1 vccd1 _7936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7867_ _8537_/CLK _7867_/D vssd1 vssd1 vccd1 vccd1 _7867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6818_ _6818_/A vssd1 vssd1 vccd1 vccd1 _6849_/B sky130_fd_sc_hd__buf_2
X_7798_ _8548_/CLK _7798_/D vssd1 vssd1 vccd1 vccd1 _7798_/Q sky130_fd_sc_hd__dfxtp_1
X_6749_ _6749_/A vssd1 vssd1 vccd1 vccd1 _6749_/X sky130_fd_sc_hd__buf_1
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8419_ _8419_/CLK _8419_/D vssd1 vssd1 vccd1 vccd1 _8419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3429_ _6949_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3429_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_104_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6182__189 _6183__190/A vssd1 vssd1 vccd1 vccd1 _7776_/CLK sky130_fd_sc_hd__inv_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4100_ _4011_/X _8409_/Q _4106_/S vssd1 vssd1 vccd1 vccd1 _4101_/A sky130_fd_sc_hd__mux2_1
X_5080_ _5080_/A vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__buf_2
X_4031_ _4295_/A vssd1 vssd1 vccd1 vccd1 _4031_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5982_ _5982_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _5983_/A sky130_fd_sc_hd__and2_1
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4933_ _5014_/A _5014_/B _4933_/C vssd1 vssd1 vccd1 vccd1 _5859_/B sky130_fd_sc_hd__nand3b_4
X_7721_ _5932_/A _7710_/X _7717_/A vssd1 vssd1 vccd1 vccd1 _7721_/X sky130_fd_sc_hd__a21bo_1
X_4864_ _8246_/Q _4781_/X _4755_/A _4863_/X vssd1 vssd1 vccd1 vccd1 _4864_/X sky130_fd_sc_hd__o211a_1
X_7652_ _7664_/A vssd1 vssd1 vccd1 vccd1 _7652_/X sky130_fd_sc_hd__buf_1
XFILLER_32_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4795_ _7849_/Q _7774_/Q _4868_/S vssd1 vssd1 vccd1 vccd1 _4795_/X sky130_fd_sc_hd__mux2_1
X_6872__371 _6873__372/A vssd1 vssd1 vccd1 vccd1 _8085_/CLK sky130_fd_sc_hd__inv_2
X_7583_ _7585_/A _7583_/B vssd1 vssd1 vccd1 vccd1 _8470_/D sky130_fd_sc_hd__nor2_1
XFILLER_118_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3315_ clkbuf_0__3315_/X vssd1 vssd1 vccd1 vccd1 _6767__355/A sky130_fd_sc_hd__clkbuf_4
X_6534_ _6540_/A vssd1 vssd1 vccd1 vccd1 _6534_/X sky130_fd_sc_hd__buf_1
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3246_ clkbuf_0__3246_/X vssd1 vssd1 vccd1 vccd1 _6538__234/A sky130_fd_sc_hd__clkbuf_4
X_6465_ _6465_/A _6465_/B _7696_/A vssd1 vssd1 vccd1 vccd1 _6466_/C sky130_fd_sc_hd__nand3_1
X_5416_ _5396_/X _8087_/Q _5420_/S vssd1 vssd1 vccd1 vccd1 _5417_/A sky130_fd_sc_hd__mux2_1
X_8204_ _8204_/CLK _8204_/D vssd1 vssd1 vccd1 vccd1 _8204_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput142 _5931_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput120 _5974_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[1] sky130_fd_sc_hd__buf_2
Xoutput131 _5981_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[4] sky130_fd_sc_hd__buf_2
X_7048__492 _7049__493/A vssd1 vssd1 vccd1 vccd1 _8219_/CLK sky130_fd_sc_hd__inv_2
X_6396_ _6362_/A _7972_/Q _6410_/C _7010_/B vssd1 vssd1 vccd1 vccd1 _6396_/X sky130_fd_sc_hd__a31o_1
Xoutput175 _5887_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_we_o sky130_fd_sc_hd__buf_2
Xoutput153 _5953_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput164 _5911_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8135_ _8135_/CLK _8135_/D vssd1 vssd1 vccd1 vccd1 _8135_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput186 _6113_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[18] sky130_fd_sc_hd__buf_2
X_5347_ _5347_/A vssd1 vssd1 vccd1 vccd1 _8119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8066_ _8066_/CLK _8066_/D vssd1 vssd1 vccd1 vccd1 _8066_/Q sky130_fd_sc_hd__dfxtp_1
X_5278_ _5193_/X _5276_/X _5277_/X vssd1 vssd1 vccd1 vccd1 _5278_/Y sky130_fd_sc_hd__o21ai_1
Xoutput197 _6146_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[28] sky130_fd_sc_hd__buf_2
X_4229_ _8374_/Q _4160_/X _4229_/S vssd1 vssd1 vccd1 vccd1 _4230_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3462_ clkbuf_0__3462_/X vssd1 vssd1 vccd1 vccd1 _7118__549/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7919_ _7919_/CLK _7919_/D vssd1 vssd1 vccd1 vccd1 _7919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 caravel_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 _6143_/A sky130_fd_sc_hd__clkbuf_4
Xinput11 caravel_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_4
X_4580_ _4580_/A vssd1 vssd1 vccd1 vccd1 _8207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput33 caravel_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
Xinput55 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _3868_/B sky130_fd_sc_hd__clkbuf_1
Xinput44 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 _3871_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_115_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput66 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _5986_/A sky130_fd_sc_hd__buf_4
Xinput77 wbs_data_i[16] vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__buf_4
Xinput88 wbs_data_i[26] vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__buf_4
X_6250_ _7631_/A _7811_/Q _6258_/S vssd1 vssd1 vccd1 vccd1 _6251_/A sky130_fd_sc_hd__mux2_1
Xinput99 wbs_data_i[7] vssd1 vssd1 vccd1 vccd1 _7646_/A sky130_fd_sc_hd__buf_4
X_5201_ _5221_/A vssd1 vssd1 vccd1 vccd1 _5352_/B sky130_fd_sc_hd__buf_2
XFILLER_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5132_ _5092_/X _5130_/X _5131_/X vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5063_ _5070_/B _5063_/B vssd1 vssd1 vccd1 vccd1 _5100_/A sky130_fd_sc_hd__or2_2
XFILLER_84_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6566__256 _6568__258/A vssd1 vssd1 vccd1 vccd1 _7934_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4014_ _8493_/Q vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__buf_4
XFILLER_53_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5965_ _5965_/A _5965_/B vssd1 vssd1 vccd1 vccd1 _5966_/A sky130_fd_sc_hd__or2_1
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5896_ _6690_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5897_/A sky130_fd_sc_hd__and2_1
X_4916_ _4811_/A _7902_/Q _4797_/X _8135_/Q _4733_/A vssd1 vssd1 vccd1 vccd1 _4916_/X
+ sky130_fd_sc_hd__o221a_1
X_7704_ _7719_/A vssd1 vssd1 vccd1 vccd1 _7704_/X sky130_fd_sc_hd__clkbuf_2
X_4847_ _7920_/Q _8024_/Q _4883_/S vssd1 vssd1 vccd1 vccd1 _4847_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7635_ _7635_/A _7637_/B _7640_/C vssd1 vssd1 vccd1 vccd1 _7636_/A sky130_fd_sc_hd__and3_1
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4778_ _8338_/Q _4775_/X _8146_/Q _4777_/X _4654_/A vssd1 vssd1 vccd1 vccd1 _4778_/X
+ sky130_fd_sc_hd__o221a_1
X_7566_ _7564_/Y _7542_/X _7555_/X _7565_/Y vssd1 vssd1 vccd1 vccd1 _7567_/B sky130_fd_sc_hd__o22a_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7497_ _7497_/A _8459_/Q vssd1 vssd1 vccd1 vccd1 _7609_/A sky130_fd_sc_hd__or2_1
X_6517_ _6517_/A _6521_/C vssd1 vssd1 vccd1 vccd1 _6517_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6448_ _7870_/Q _6442_/X _6437_/X _6447_/X _6435_/X vssd1 vssd1 vccd1 vccd1 _7870_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6379_ _8528_/Q _6356_/X _6378_/X _6350_/X _6358_/X vssd1 vssd1 vccd1 vccd1 _6379_/X
+ sky130_fd_sc_hd__a221o_1
X_8118_ _8118_/CLK _8118_/D vssd1 vssd1 vccd1 vccd1 _8118_/Q sky130_fd_sc_hd__dfxtp_2
X_8049_ _8049_/CLK _8049_/D vssd1 vssd1 vccd1 vccd1 _8049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3445_ clkbuf_0__3445_/X vssd1 vssd1 vccd1 vccd1 _7052_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _8368_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5750_ _5750_/A vssd1 vssd1 vccd1 vccd1 _7910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4701_ _8251_/Q _8036_/Q _7988_/Q _7940_/Q _4646_/A _4674_/X vssd1 vssd1 vccd1 vccd1
+ _4701_/X sky130_fd_sc_hd__mux4_1
X_5681_ _7941_/Q _5578_/X _5689_/S vssd1 vssd1 vccd1 vccd1 _5682_/A sky130_fd_sc_hd__mux2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7420_ _7420_/A vssd1 vssd1 vccd1 vccd1 _7420_/X sky130_fd_sc_hd__buf_1
X_4632_ _4823_/A vssd1 vssd1 vccd1 vccd1 _4947_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4563_ _4441_/X _8214_/Q _4565_/S vssd1 vssd1 vccd1 vccd1 _4564_/A sky130_fd_sc_hd__mux2_1
X_7351_ _7008_/A _7299_/B _7303_/A _7271_/Y _7350_/Y vssd1 vssd1 vccd1 vccd1 _7361_/A
+ sky130_fd_sc_hd__o221ai_4
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4494_ _4379_/X _8243_/Q _4500_/S vssd1 vssd1 vccd1 vccd1 _4495_/A sky130_fd_sc_hd__mux2_1
X_7282_ _7514_/A _7261_/B _7221_/B _7529_/A vssd1 vssd1 vccd1 vccd1 _7282_/X sky130_fd_sc_hd__o2bb2a_1
X_6945__412 _6948__415/A vssd1 vssd1 vccd1 vccd1 _8136_/CLK sky130_fd_sc_hd__inv_2
X_6233_ _6367_/A vssd1 vssd1 vccd1 vccd1 _6233_/X sky130_fd_sc_hd__buf_2
X_6164_ _6961_/A vssd1 vssd1 vccd1 vccd1 _6164_/X sky130_fd_sc_hd__buf_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5354_/B _5114_/X _5083_/X vssd1 vssd1 vccd1 vccd1 _5115_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6095_/A vssd1 vssd1 vccd1 vccd1 _6095_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5046_ _8118_/Q _5103_/B vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__xor2_2
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3092_ clkbuf_0__3092_/X vssd1 vssd1 vccd1 vccd1 _6526__225/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5948_ _5948_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _5949_/A sky130_fd_sc_hd__or2_4
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5879_ _8014_/Q _8015_/Q _8016_/Q _8017_/Q vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__and4_2
X_7158__80 _7158__80/A vssd1 vssd1 vccd1 vccd1 _8307_/CLK sky130_fd_sc_hd__inv_2
X_7618_ _8482_/Q _7613_/X _7617_/X _7552_/X vssd1 vssd1 vccd1 vccd1 _8481_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7549_ _7567_/A _7549_/B vssd1 vssd1 vccd1 vccd1 _8461_/D sky130_fd_sc_hd__nor2_1
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6885__381 _6887__383/A vssd1 vssd1 vccd1 vccd1 _8095_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3428_ clkbuf_0__3428_/X vssd1 vssd1 vccd1 vccd1 _6946__413/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__3022_ clkbuf_0__3022_/X vssd1 vssd1 vccd1 vccd1 _6297_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6851_ _6832_/Y _6833_/X _6845_/X _6848_/X _6850_/X vssd1 vssd1 vccd1 vccd1 _6855_/C
+ sky130_fd_sc_hd__o2111a_1
X_5802_ _5802_/A vssd1 vssd1 vccd1 vccd1 _7839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3994_ _3899_/X _8447_/Q _3996_/S vssd1 vssd1 vccd1 vccd1 _3995_/A sky130_fd_sc_hd__mux2_1
X_6719__321 _6720__322/A vssd1 vssd1 vccd1 vccd1 _8031_/CLK sky130_fd_sc_hd__inv_2
X_8521_ _8527_/CLK _8521_/D vssd1 vssd1 vccd1 vccd1 _8521_/Q sky130_fd_sc_hd__dfxtp_1
X_5733_ _5733_/A _5733_/B vssd1 vssd1 vccd1 vccd1 _5749_/S sky130_fd_sc_hd__nor2_2
X_5664_ _5664_/A vssd1 vssd1 vccd1 vccd1 _7949_/D sky130_fd_sc_hd__clkbuf_1
X_8452_ _8452_/CLK _8452_/D vssd1 vssd1 vccd1 vccd1 _8452_/Q sky130_fd_sc_hd__dfxtp_1
X_8383_ _8383_/CLK _8383_/D vssd1 vssd1 vccd1 vccd1 _8383_/Q sky130_fd_sc_hd__dfxtp_1
X_4615_ _4615_/A vssd1 vssd1 vccd1 vccd1 _8192_/D sky130_fd_sc_hd__clkbuf_1
X_5595_ _5595_/A vssd1 vssd1 vccd1 vccd1 _7984_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3462_ _7114_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3462_/X sky130_fd_sc_hd__clkbuf_16
X_4546_ _4546_/A vssd1 vssd1 vccd1 vccd1 _8222_/D sky130_fd_sc_hd__clkbuf_1
X_7334_ _7334_/A vssd1 vssd1 vccd1 vccd1 _7334_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4477_ _4477_/A vssd1 vssd1 vccd1 vccd1 _8249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7265_ _8534_/Q _7308_/A vssd1 vssd1 vccd1 vccd1 _7365_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7196_ _8354_/Q _8353_/Q _8352_/Q _8351_/Q vssd1 vssd1 vccd1 vccd1 _7197_/D sky130_fd_sc_hd__and4_1
X_6216_ _6208_/X _8002_/Q _6211_/X _6213_/X _7791_/Q vssd1 vssd1 vccd1 vccd1 _7791_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6147_ _6147_/A _6151_/B vssd1 vssd1 vccd1 vccd1 _6147_/X sky130_fd_sc_hd__and2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_24 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_13 _8392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_35 _6123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_68 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6078_ _7788_/Q _6086_/B vssd1 vssd1 vccd1 vccd1 _6078_/X sky130_fd_sc_hd__or2_1
XINSDIODE2_46 _6135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_57 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_79 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5029_ _4441_/X _8136_/Q _5031_/S vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ _4531_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _4416_/S sky130_fd_sc_hd__or2_2
X_5380_ _5379_/X _8100_/Q _5388_/S vssd1 vssd1 vccd1 vccd1 _5381_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4331_ _4331_/A vssd1 vssd1 vccd1 vccd1 _8304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4262_ _4262_/A vssd1 vssd1 vccd1 vccd1 _8331_/D sky130_fd_sc_hd__clkbuf_1
X_6001_ _6001_/A vssd1 vssd1 vccd1 vccd1 _6001_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4193_ _8489_/Q vssd1 vssd1 vccd1 vccd1 _4193_/X sky130_fd_sc_hd__clkbuf_2
X_7042__487 _7043__488/A vssd1 vssd1 vccd1 vccd1 _8214_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7952_ _7952_/CLK _7952_/D vssd1 vssd1 vccd1 vccd1 _7952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6903_ _8482_/Q _6911_/B vssd1 vssd1 vccd1 vccd1 _6904_/A sky130_fd_sc_hd__and2_1
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7883_ _8551_/CLK _7883_/D vssd1 vssd1 vccd1 vccd1 _7883_/Q sky130_fd_sc_hd__dfxtp_1
X_8574__221 vssd1 vssd1 vccd1 vccd1 _8574__221/HI core1Index[1] sky130_fd_sc_hd__conb_1
XFILLER_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6834_ _8462_/Q vssd1 vssd1 vccd1 vccd1 _7550_/A sky130_fd_sc_hd__buf_2
X_3977_ _3977_/A vssd1 vssd1 vccd1 vccd1 _8453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3477_ clkbuf_0__3477_/X vssd1 vssd1 vccd1 vccd1 _7189__105/A sky130_fd_sc_hd__clkbuf_4
X_8504_ _8504_/CLK _8504_/D vssd1 vssd1 vccd1 vccd1 _8504_/Q sky130_fd_sc_hd__dfxtp_1
X_5716_ _5731_/S vssd1 vssd1 vccd1 vccd1 _5725_/S sky130_fd_sc_hd__clkbuf_2
X_7446__161 _7447__162/A vssd1 vssd1 vccd1 vccd1 _8418_/CLK sky130_fd_sc_hd__inv_2
X_8435_ _8435_/CLK _8435_/D vssd1 vssd1 vccd1 vccd1 _8435_/Q sky130_fd_sc_hd__dfxtp_1
X_6696_ _8016_/Q _5959_/A _6700_/S vssd1 vssd1 vccd1 vccd1 _6697_/A sky130_fd_sc_hd__mux2_1
X_5647_ _8111_/Q vssd1 vssd1 vccd1 vccd1 _5647_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3445_ _7027_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3445_/X sky130_fd_sc_hd__clkbuf_16
X_5578_ _8113_/Q vssd1 vssd1 vccd1 vccd1 _5578_/X sky130_fd_sc_hd__buf_4
X_8366_ _8368_/CLK _8366_/D vssd1 vssd1 vccd1 vccd1 _8366_/Q sky130_fd_sc_hd__dfxtp_1
X_4529_ _8229_/Q _4487_/X _4529_/S vssd1 vssd1 vccd1 vccd1 _4530_/A sky130_fd_sc_hd__mux2_1
X_8297_ _8297_/CLK _8297_/D vssd1 vssd1 vccd1 vccd1 _8297_/Q sky130_fd_sc_hd__dfxtp_1
X_7317_ _7321_/A _7317_/B vssd1 vssd1 vccd1 vccd1 _8347_/D sky130_fd_sc_hd__nor2_1
XFILLER_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7248_ _8551_/Q _7302_/A vssd1 vssd1 vccd1 vccd1 _7248_/X sky130_fd_sc_hd__or2_1
XFILLER_58_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 caravel_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3900_ _3899_/X _8516_/Q _3903_/S vssd1 vssd1 vccd1 vccd1 _3901_/A sky130_fd_sc_hd__mux2_1
X_4880_ _7911_/Q _8083_/Q _4880_/S vssd1 vssd1 vccd1 vccd1 _4880_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3831_ _8495_/Q vssd1 vssd1 vccd1 vccd1 _3831_/X sky130_fd_sc_hd__buf_4
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5501_ _5516_/S vssd1 vssd1 vccd1 vccd1 _5510_/S sky130_fd_sc_hd__buf_2
XFILLER_118_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6481_ _5989_/A _7883_/Q _6487_/S vssd1 vssd1 vccd1 vccd1 _6482_/A sky130_fd_sc_hd__mux2_1
X_5432_ _3963_/X _8079_/Q _5438_/S vssd1 vssd1 vccd1 vccd1 _5433_/A sky130_fd_sc_hd__mux2_1
X_8220_ _8220_/CLK _8220_/D vssd1 vssd1 vccd1 vccd1 _8220_/Q sky130_fd_sc_hd__dfxtp_1
X_5363_ _5388_/S vssd1 vssd1 vccd1 vccd1 _5376_/S sky130_fd_sc_hd__buf_2
X_8151_ _8151_/CLK _8151_/D vssd1 vssd1 vccd1 vccd1 _8151_/Q sky130_fd_sc_hd__dfxtp_1
X_7125__53 _7127__55/A vssd1 vssd1 vccd1 vccd1 _8280_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4314_ _4292_/X _8311_/Q _4318_/S vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__mux2_1
X_7102_ _7108_/A vssd1 vssd1 vccd1 vccd1 _7102_/X sky130_fd_sc_hd__buf_1
XFILLER_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5294_ _5352_/B _5283_/Y _5286_/Y _5293_/X _5350_/B vssd1 vssd1 vccd1 vccd1 _5295_/B
+ sky130_fd_sc_hd__a311o_1
X_8082_ _8082_/CLK _8082_/D vssd1 vssd1 vccd1 vccd1 _8082_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3092_ _6322_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3092_/X sky130_fd_sc_hd__clkbuf_16
X_4245_ _4245_/A vssd1 vssd1 vccd1 vccd1 _8340_/D sky130_fd_sc_hd__clkbuf_1
X_4176_ _8394_/Q _4172_/X _4188_/S vssd1 vssd1 vccd1 vccd1 _4177_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7935_ _7935_/CLK _7935_/D vssd1 vssd1 vccd1 vccd1 _7935_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7866_ _8550_/CLK _7866_/D vssd1 vssd1 vccd1 vccd1 _7866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6817_ _7529_/A _7525_/B vssd1 vssd1 vccd1 vccd1 _6855_/A sky130_fd_sc_hd__xor2_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7797_ _8537_/CLK _7797_/D vssd1 vssd1 vccd1 vccd1 _7797_/Q sky130_fd_sc_hd__dfxtp_1
X_6679_ _6679_/A vssd1 vssd1 vccd1 vccd1 _8008_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8418_ _8418_/CLK _8418_/D vssd1 vssd1 vccd1 vccd1 _8418_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3428_ _6943_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3428_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8349_ _8358_/CLK _8349_/D vssd1 vssd1 vccd1 vccd1 _8349_/Q sky130_fd_sc_hd__dfxtp_1
X_7667__43 _7669__45/A vssd1 vssd1 vccd1 vccd1 _8512_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4030_ _8489_/Q vssd1 vssd1 vccd1 vccd1 _4295_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5981_ _5981_/A vssd1 vssd1 vccd1 vccd1 _5981_/X sky130_fd_sc_hd__clkbuf_1
X_6306__207 _6306__207/A vssd1 vssd1 vccd1 vccd1 _7837_/CLK sky130_fd_sc_hd__inv_2
X_4932_ _5769_/A vssd1 vssd1 vccd1 vccd1 _5733_/A sky130_fd_sc_hd__clkbuf_4
X_7720_ _7201_/A _7717_/X _7718_/X _7719_/X vssd1 vssd1 vccd1 vccd1 _8536_/D sky130_fd_sc_hd__o211a_1
XFILLER_45_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6602_ _6626_/A vssd1 vssd1 vccd1 vccd1 _6602_/X sky130_fd_sc_hd__buf_1
X_4863_ _7935_/Q _4784_/A _4862_/X _4787_/X vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__o22a_1
X_4794_ _4803_/A vssd1 vssd1 vccd1 vccd1 _4794_/X sky130_fd_sc_hd__buf_2
X_7582_ _7581_/Y _7570_/X _7575_/X _7529_/B vssd1 vssd1 vccd1 vccd1 _7583_/B sky130_fd_sc_hd__o22a_1
XFILLER_20_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3245_ clkbuf_0__3245_/X vssd1 vssd1 vccd1 vccd1 _6530__227/A sky130_fd_sc_hd__clkbuf_4
X_6464_ _6388_/X _6521_/B _6522_/A _7876_/Q _7687_/A vssd1 vssd1 vccd1 vccd1 _7876_/D
+ sky130_fd_sc_hd__o221a_1
Xoutput110 _5994_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[10] sky130_fd_sc_hd__buf_2
XFILLER_118_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5415_ _5415_/A vssd1 vssd1 vccd1 vccd1 _8088_/D sky130_fd_sc_hd__clkbuf_1
X_8203_ _8203_/CLK _8203_/D vssd1 vssd1 vccd1 vccd1 _8203_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput121 _6016_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput132 _5983_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[5] sky130_fd_sc_hd__buf_2
Xoutput143 _5933_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[14] sky130_fd_sc_hd__buf_2
X_6395_ _6395_/A vssd1 vssd1 vccd1 vccd1 _7010_/B sky130_fd_sc_hd__clkbuf_2
Xoutput154 _5955_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput165 _5914_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_114_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput176 _6157_/X vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
X_8134_ _8530_/CLK _8134_/D vssd1 vssd1 vccd1 vccd1 _8134_/Q sky130_fd_sc_hd__dfxtp_1
X_5346_ _5346_/A _6941_/B _5346_/C vssd1 vssd1 vccd1 vccd1 _5347_/A sky130_fd_sc_hd__and3_1
XFILLER_102_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8065_ _8065_/CLK _8065_/D vssd1 vssd1 vccd1 vccd1 _8065_/Q sky130_fd_sc_hd__dfxtp_1
X_5277_ _8310_/Q _5196_/X _5239_/X _8302_/Q _5167_/S vssd1 vssd1 vccd1 vccd1 _5277_/X
+ sky130_fd_sc_hd__o221a_1
Xoutput187 _6117_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput198 _6148_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[29] sky130_fd_sc_hd__buf_2
X_4228_ _4228_/A vssd1 vssd1 vccd1 vccd1 _8375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3461_ clkbuf_0__3461_/X vssd1 vssd1 vccd1 vccd1 _7113__545/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4159_ _4159_/A vssd1 vssd1 vccd1 vccd1 _8399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7918_ _7918_/CLK _7918_/D vssd1 vssd1 vccd1 vccd1 _7918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7849_ _7849_/CLK _7849_/D vssd1 vssd1 vccd1 vccd1 _7849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6292__196 _6294__198/A vssd1 vssd1 vccd1 vccd1 _7826_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 caravel_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 caravel_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 _6145_/A sky130_fd_sc_hd__clkbuf_4
Xinput34 caravel_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_4
X_6713__316 _6716__319/A vssd1 vssd1 vccd1 vccd1 _8026_/CLK sky130_fd_sc_hd__inv_2
Xinput45 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _3871_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput67 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _5989_/A sky130_fd_sc_hd__buf_4
Xinput78 wbs_data_i[17] vssd1 vssd1 vccd1 vccd1 _5939_/A sky130_fd_sc_hd__buf_4
Xinput89 wbs_data_i[27] vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__buf_4
Xinput56 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _3868_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5200_ _5193_/X _5195_/X _5199_/X vssd1 vssd1 vccd1 vccd1 _5200_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5131_ _5221_/A vssd1 vssd1 vccd1 vccd1 _5131_/X sky130_fd_sc_hd__buf_2
X_5062_ _7845_/Q _8053_/Q _8332_/Q _8080_/Q _5284_/S _5061_/X vssd1 vssd1 vccd1 vccd1
+ _5062_/X sky130_fd_sc_hd__mux4_1
X_4013_ _4013_/A vssd1 vssd1 vccd1 vccd1 _8441_/D sky130_fd_sc_hd__clkbuf_1
X_7661__38 _7663__40/A vssd1 vssd1 vccd1 vccd1 _8507_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5964_ _5964_/A vssd1 vssd1 vccd1 vccd1 _5964_/X sky130_fd_sc_hd__clkbuf_1
X_7703_ _5946_/A _7702_/X _7701_/A vssd1 vssd1 vccd1 vccd1 _7703_/X sky130_fd_sc_hd__a21bo_1
X_5895_ _5895_/A vssd1 vssd1 vccd1 vccd1 _5895_/X sky130_fd_sc_hd__clkbuf_1
X_4915_ _7918_/Q _8022_/Q _4915_/S vssd1 vssd1 vccd1 vccd1 _4915_/X sky130_fd_sc_hd__mux2_1
X_4846_ _4770_/X _4844_/X _4845_/X vssd1 vssd1 vccd1 vccd1 _4846_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7634_ _7634_/A vssd1 vssd1 vccd1 vccd1 _8489_/D sky130_fd_sc_hd__clkbuf_1
X_7565_ _7565_/A _7565_/B vssd1 vssd1 vccd1 vccd1 _7565_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4777_ _4806_/A vssd1 vssd1 vccd1 vccd1 _4777_/X sky130_fd_sc_hd__clkbuf_2
X_6516_ _6269_/C _6284_/X _6456_/B vssd1 vssd1 vccd1 vccd1 _6521_/C sky130_fd_sc_hd__a21oi_1
XFILLER_119_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6447_ _8535_/Q _6452_/B _6454_/C vssd1 vssd1 vccd1 vccd1 _6447_/X sky130_fd_sc_hd__and3_1
X_6378_ _7741_/A _7969_/Q _6352_/X _6364_/X vssd1 vssd1 vccd1 vccd1 _6378_/X sky130_fd_sc_hd__a31o_1
XFILLER_114_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8117_ _8117_/CLK _8117_/D vssd1 vssd1 vccd1 vccd1 _8117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5329_ _8124_/Q _5106_/A _5345_/B _5262_/X vssd1 vssd1 vccd1 vccd1 _8124_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8048_ _8048_/CLK _8048_/D vssd1 vssd1 vccd1 vccd1 _8048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3444_ clkbuf_0__3444_/X vssd1 vssd1 vccd1 vccd1 _7026__475/A sky130_fd_sc_hd__clkbuf_4
XFILLER_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8554__252 vssd1 vssd1 vccd1 vccd1 partID[2] _8554__252/LO sky130_fd_sc_hd__conb_1
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7486__19 _7487__20/A vssd1 vssd1 vccd1 vccd1 _8451_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7105__538 _7106__539/A vssd1 vssd1 vccd1 vccd1 _8265_/CLK sky130_fd_sc_hd__inv_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5680_ _5695_/S vssd1 vssd1 vccd1 vccd1 _5689_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4664_/X _4697_/X _4699_/X vssd1 vssd1 vccd1 vccd1 _4700_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4631_ _4713_/A _6605_/B vssd1 vssd1 vccd1 vccd1 _4823_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6572__261 _6574__263/A vssd1 vssd1 vccd1 vccd1 _7939_/CLK sky130_fd_sc_hd__inv_2
X_4562_ _4562_/A vssd1 vssd1 vccd1 vccd1 _8215_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7350_ _7355_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7350_/Y sky130_fd_sc_hd__nor2_1
X_4493_ _4493_/A vssd1 vssd1 vccd1 vccd1 _8244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7281_ _7281_/A _7281_/B _7281_/C _7281_/D vssd1 vssd1 vccd1 vccd1 _7281_/X sky130_fd_sc_hd__and4_1
XFILLER_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7440__156 _7441__157/A vssd1 vssd1 vccd1 vccd1 _8413_/CLK sky130_fd_sc_hd__inv_2
X_6232_ _6225_/X _8012_/Q _6227_/X _6229_/X _7801_/Q vssd1 vssd1 vccd1 vccd1 _7801_/D
+ sky130_fd_sc_hd__o32a_1
X_6163_ _6163_/A vssd1 vssd1 vccd1 vccd1 _6163_/X sky130_fd_sc_hd__buf_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _8441_/Q _8433_/Q _7836_/Q _8449_/Q _5066_/X _5080_/X vssd1 vssd1 vccd1 vccd1
+ _5114_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6075_/X _6092_/X _6093_/X _6083_/X vssd1 vssd1 vccd1 vccd1 _6094_/X sky130_fd_sc_hd__o211a_1
XFILLER_85_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5045_ _5045_/A vssd1 vssd1 vccd1 vccd1 _5103_/B sky130_fd_sc_hd__clkbuf_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5947_ _5947_/A vssd1 vssd1 vccd1 vccd1 _5947_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__3091_ clkbuf_0__3091_/X vssd1 vssd1 vccd1 vccd1 _6318__217/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5878_ _6035_/A _5878_/B vssd1 vssd1 vccd1 vccd1 _5881_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7617_ _8481_/Q _7614_/X vssd1 vssd1 vccd1 vccd1 _7617_/X sky130_fd_sc_hd__or2b_1
X_4829_ _4770_/X _4827_/X _4828_/X vssd1 vssd1 vccd1 vccd1 _4829_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7548_ _7547_/X _7588_/A _7548_/S vssd1 vssd1 vccd1 vccd1 _7549_/B sky130_fd_sc_hd__mux2_1
XFILLER_111_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8591__238 vssd1 vssd1 vccd1 vccd1 _8591__238/HI manufacturerID[10] sky130_fd_sc_hd__conb_1
XFILLER_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6850_ _8547_/Q _7522_/B vssd1 vssd1 vccd1 vccd1 _6850_/X sky130_fd_sc_hd__xor2_1
XFILLER_23_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5801_ _7839_/Q _4295_/A _5803_/S vssd1 vssd1 vccd1 vccd1 _5802_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3993_ _3993_/A vssd1 vssd1 vccd1 vccd1 _8448_/D sky130_fd_sc_hd__clkbuf_1
X_5732_ _5732_/A vssd1 vssd1 vccd1 vccd1 _7918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8520_ _8520_/CLK _8520_/D vssd1 vssd1 vccd1 vccd1 _8520_/Q sky130_fd_sc_hd__dfxtp_1
X_5663_ _5554_/X _7949_/Q _5671_/S vssd1 vssd1 vccd1 vccd1 _5664_/A sky130_fd_sc_hd__mux2_1
X_8451_ _8451_/CLK _8451_/D vssd1 vssd1 vccd1 vccd1 _8451_/Q sky130_fd_sc_hd__dfxtp_1
X_7402_ _7426_/A vssd1 vssd1 vccd1 vccd1 _7402_/X sky130_fd_sc_hd__buf_1
X_8382_ _8382_/CLK _8382_/D vssd1 vssd1 vccd1 vccd1 _8382_/Q sky130_fd_sc_hd__dfxtp_1
X_5594_ _7984_/Q _5593_/X _5600_/S vssd1 vssd1 vccd1 vccd1 _5595_/A sky130_fd_sc_hd__mux2_1
X_4614_ _8192_/Q _4187_/X _4614_/S vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3461_ _7108_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3461_/X sky130_fd_sc_hd__clkbuf_16
X_4545_ _4394_/X _8222_/Q _4547_/S vssd1 vssd1 vccd1 vccd1 _4546_/A sky130_fd_sc_hd__mux2_1
X_7333_ _7336_/A _7333_/B vssd1 vssd1 vccd1 vccd1 _8352_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4476_ _8249_/Q _4157_/X _4479_/S vssd1 vssd1 vccd1 vccd1 _4477_/A sky130_fd_sc_hd__mux2_1
X_7264_ _7308_/B vssd1 vssd1 vccd1 vccd1 _7303_/A sky130_fd_sc_hd__clkbuf_2
X_6215_ _6208_/X _8001_/Q _6211_/X _6213_/X _7790_/Q vssd1 vssd1 vccd1 vccd1 _7790_/D
+ sky130_fd_sc_hd__o32a_1
X_7195_ _8350_/Q _8349_/Q _8348_/Q _8347_/Q vssd1 vssd1 vccd1 vccd1 _7232_/C sky130_fd_sc_hd__and4_2
XFILLER_112_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6765__353 _6767__355/A vssd1 vssd1 vccd1 vccd1 _8066_/CLK sky130_fd_sc_hd__inv_2
X_6146_ _7807_/Q _6138_/X _6139_/X _6145_/X _6136_/X vssd1 vssd1 vccd1 vccd1 _6146_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_25 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_14 _8394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6726__326 _6727__327/A vssd1 vssd1 vccd1 vccd1 _8036_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_47 _6135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_36 _6123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_58 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6077_ _7863_/Q input34/X _6092_/S vssd1 vssd1 vccd1 vccd1 _6077_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5028_ _5028_/A vssd1 vssd1 vccd1 vccd1 _8137_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_69 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6579__267 _6579__267/A vssd1 vssd1 vccd1 vccd1 _7945_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4289_/X _8304_/Q _4330_/S vssd1 vssd1 vccd1 vccd1 _4331_/A sky130_fd_sc_hd__mux2_1
X_4261_ _8331_/Q _4178_/X _4267_/S vssd1 vssd1 vccd1 vccd1 _4262_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6000_ _6000_/A _6008_/B vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__and2_1
XFILLER_113_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4192_ _4192_/A vssd1 vssd1 vccd1 vccd1 _8389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7951_ _7951_/CLK _7951_/D vssd1 vssd1 vccd1 vccd1 _7951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7882_ _8551_/CLK _7882_/D vssd1 vssd1 vccd1 vccd1 _7882_/Q sky130_fd_sc_hd__dfxtp_1
X_6902_ _6902_/A vssd1 vssd1 vccd1 vccd1 _6911_/B sky130_fd_sc_hd__clkbuf_1
X_6833_ _8546_/Q _7565_/A _7565_/B vssd1 vssd1 vccd1 vccd1 _6833_/X sky130_fd_sc_hd__and3_1
XFILLER_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3976_ _8453_/Q _3975_/X _3982_/S vssd1 vssd1 vccd1 vccd1 _3977_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8503_ _8503_/CLK _8503_/D vssd1 vssd1 vccd1 vccd1 _8503_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3476_ clkbuf_0__3476_/X vssd1 vssd1 vccd1 vccd1 _7389_/A sky130_fd_sc_hd__clkbuf_4
X_5715_ _5733_/A _5751_/B vssd1 vssd1 vccd1 vccd1 _5731_/S sky130_fd_sc_hd__nor2_2
X_6695_ _6695_/A vssd1 vssd1 vccd1 vccd1 _8015_/D sky130_fd_sc_hd__clkbuf_1
X_5646_ _5646_/A vssd1 vssd1 vccd1 vccd1 _7956_/D sky130_fd_sc_hd__clkbuf_1
X_8434_ _8434_/CLK _8434_/D vssd1 vssd1 vccd1 vccd1 _8434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5577_ _5577_/A vssd1 vssd1 vccd1 vccd1 _7990_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3444_ _7021_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3444_/X sky130_fd_sc_hd__clkbuf_16
X_8365_ _8368_/CLK _8365_/D vssd1 vssd1 vccd1 vccd1 _8365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4528_ _4528_/A vssd1 vssd1 vccd1 vccd1 _8230_/D sky130_fd_sc_hd__clkbuf_1
X_8296_ _8296_/CLK _8296_/D vssd1 vssd1 vccd1 vccd1 _8296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7316_ _7236_/A _7301_/X _7310_/X _7237_/B vssd1 vssd1 vccd1 vccd1 _7317_/B sky130_fd_sc_hd__o2bb2a_1
X_4459_ _4391_/X _8255_/Q _4463_/S vssd1 vssd1 vccd1 vccd1 _4460_/A sky130_fd_sc_hd__mux2_1
X_7247_ _7247_/A _7302_/A vssd1 vssd1 vccd1 vccd1 _7247_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6129_ _6129_/A _6140_/B vssd1 vssd1 vccd1 vccd1 _6129_/X sky130_fd_sc_hd__and2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6958__423 _6960__425/A vssd1 vssd1 vccd1 vccd1 _8147_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6965__427 _6968__430/A vssd1 vssd1 vccd1 vccd1 _8151_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8597__244 vssd1 vssd1 vccd1 vccd1 _8597__244/HI partID[12] sky130_fd_sc_hd__conb_1
XFILLER_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5500_ _5500_/A _5500_/B vssd1 vssd1 vccd1 vccd1 _5516_/S sky130_fd_sc_hd__nor2_2
X_6480_ _6480_/A vssd1 vssd1 vccd1 vccd1 _7882_/D sky130_fd_sc_hd__clkbuf_1
X_5431_ _5431_/A vssd1 vssd1 vccd1 vccd1 _8080_/D sky130_fd_sc_hd__clkbuf_1
X_8150_ _8150_/CLK _8150_/D vssd1 vssd1 vccd1 vccd1 _8150_/Q sky130_fd_sc_hd__dfxtp_1
X_5362_ _5555_/A _5841_/A vssd1 vssd1 vccd1 vccd1 _5388_/S sky130_fd_sc_hd__or2_2
X_4313_ _4313_/A vssd1 vssd1 vccd1 vccd1 _8312_/D sky130_fd_sc_hd__clkbuf_1
X_8081_ _8487_/CLK _8081_/D vssd1 vssd1 vccd1 vccd1 _8081_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5293_ _5293_/A _5293_/B _5293_/C vssd1 vssd1 vccd1 vccd1 _5293_/X sky130_fd_sc_hd__and3_1
Xclkbuf_0__3091_ _6316_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3091_/X sky130_fd_sc_hd__clkbuf_16
X_4244_ _8340_/Q _4154_/X _4248_/S vssd1 vssd1 vccd1 vccd1 _4245_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4175_ _4197_/S vssd1 vssd1 vccd1 vccd1 _4188_/S sky130_fd_sc_hd__buf_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7934_ _7934_/CLK _7934_/D vssd1 vssd1 vccd1 vccd1 _7934_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7865_ _8550_/CLK _7865_/D vssd1 vssd1 vccd1 vccd1 _7865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6816_ _6816_/A _6816_/B vssd1 vssd1 vccd1 vccd1 _7525_/B sky130_fd_sc_hd__xnor2_4
X_7796_ _8537_/CLK _7796_/D vssd1 vssd1 vccd1 vccd1 _7796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3959_ _4604_/A _5500_/B vssd1 vssd1 vccd1 vccd1 _3982_/S sky130_fd_sc_hd__nor2_2
XFILLER_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3459_ clkbuf_0__3459_/X vssd1 vssd1 vccd1 vccd1 _7101__535/A sky130_fd_sc_hd__clkbuf_4
X_6678_ _5941_/A _8008_/Q _6682_/S vssd1 vssd1 vccd1 vccd1 _6679_/A sky130_fd_sc_hd__mux2_1
X_8417_ _8417_/CLK _8417_/D vssd1 vssd1 vccd1 vccd1 _8417_/Q sky130_fd_sc_hd__dfxtp_1
X_5629_ _5608_/X _7963_/Q _5633_/S vssd1 vssd1 vccd1 vccd1 _5630_/A sky130_fd_sc_hd__mux2_1
X_8348_ _8370_/CLK _8348_/D vssd1 vssd1 vccd1 vccd1 _8348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8279_ _8279_/CLK _8279_/D vssd1 vssd1 vccd1 vccd1 _8279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _5980_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__and2_1
XFILLER_92_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _4931_/A _4931_/B vssd1 vssd1 vccd1 vccd1 _5769_/A sky130_fd_sc_hd__or2_4
X_4862_ _7983_/Q _8031_/Q _4883_/S vssd1 vssd1 vccd1 vccd1 _4862_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3313_ clkbuf_0__3313_/X vssd1 vssd1 vccd1 vccd1 _6754__350/A sky130_fd_sc_hd__clkbuf_4
X_4793_ _7825_/Q _4791_/X _4787_/X _4792_/X vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__o22a_1
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7581_ _8470_/Q vssd1 vssd1 vccd1 vccd1 _7581_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7473__8 _7474__9/A vssd1 vssd1 vccd1 vccd1 _8440_/CLK sky130_fd_sc_hd__inv_2
X_6536__232 _6538__234/A vssd1 vssd1 vccd1 vccd1 _7910_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3244_ clkbuf_0__3244_/X vssd1 vssd1 vccd1 vccd1 _6552_/A sky130_fd_sc_hd__clkbuf_4
X_6463_ _7689_/A vssd1 vssd1 vccd1 vccd1 _7687_/A sky130_fd_sc_hd__buf_2
X_7404__127 _7405__128/A vssd1 vssd1 vccd1 vccd1 _8384_/CLK sky130_fd_sc_hd__inv_2
X_8202_ _8202_/CLK _8202_/D vssd1 vssd1 vccd1 vccd1 _8202_/Q sky130_fd_sc_hd__dfxtp_1
X_5414_ _5367_/X _8088_/Q _5420_/S vssd1 vssd1 vccd1 vccd1 _5415_/A sky130_fd_sc_hd__mux2_1
Xoutput111 _5996_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[11] sky130_fd_sc_hd__buf_2
Xoutput122 _6018_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput133 _5985_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[6] sky130_fd_sc_hd__buf_2
X_6394_ _7859_/Q _6388_/X _6393_/X vssd1 vssd1 vccd1 vccd1 _7859_/D sky130_fd_sc_hd__a21o_1
X_8133_ _8530_/CLK _8133_/D vssd1 vssd1 vccd1 vccd1 _8133_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput155 _5958_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput166 _5916_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[6] sky130_fd_sc_hd__buf_2
Xoutput144 _5936_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_102_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput177 _6045_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[0] sky130_fd_sc_hd__buf_2
X_5345_ _5345_/A _5345_/B vssd1 vssd1 vccd1 vccd1 _5346_/C sky130_fd_sc_hd__nand2_1
XFILLER_114_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5276_ _8286_/Q _8294_/Q _5315_/S vssd1 vssd1 vccd1 vccd1 _5276_/X sky130_fd_sc_hd__mux2_1
Xoutput188 _6048_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput199 _6052_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[2] sky130_fd_sc_hd__buf_2
X_8064_ _8548_/CLK _8064_/D vssd1 vssd1 vccd1 vccd1 _8064_/Q sky130_fd_sc_hd__dfxtp_1
X_4227_ _8375_/Q _4157_/X _4229_/S vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__3460_ clkbuf_0__3460_/X vssd1 vssd1 vccd1 vccd1 _7107__540/A sky130_fd_sc_hd__clkbuf_4
X_7015_ _7021_/A vssd1 vssd1 vccd1 vccd1 _7015_/X sky130_fd_sc_hd__buf_1
XFILLER_68_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4158_ _8399_/Q _4157_/X _4161_/S vssd1 vssd1 vccd1 vccd1 _4159_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4089_ _4089_/A vssd1 vssd1 vccd1 vccd1 _8414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6920__396 _6923__399/A vssd1 vssd1 vccd1 vccd1 _8118_/CLK sky130_fd_sc_hd__inv_2
X_7917_ _7917_/CLK _7917_/D vssd1 vssd1 vccd1 vccd1 _7917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7848_ _7848_/CLK _7848_/D vssd1 vssd1 vccd1 vccd1 _7848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7055__498 _7057__500/A vssd1 vssd1 vccd1 vccd1 _8225_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7779_ _8355_/CLK _7779_/D vssd1 vssd1 vccd1 vccd1 _7779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7459__172 _7460__173/A vssd1 vssd1 vccd1 vccd1 _8429_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3658_ clkbuf_0__3658_/X vssd1 vssd1 vccd1 vccd1 _7650__29/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3321_ clkbuf_0__3321_/X vssd1 vssd1 vccd1 vccd1 _6782__367/A sky130_fd_sc_hd__clkbuf_16
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 caravel_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_4
Xinput24 caravel_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 _6147_/A sky130_fd_sc_hd__clkbuf_4
Xinput35 caravel_wb_error_i vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_4
Xinput46 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _3866_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_116_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput57 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
Xinput79 wbs_data_i[18] vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__buf_4
Xinput68 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _5991_/A sky130_fd_sc_hd__buf_4
XFILLER_6_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6312__212 _6312__212/A vssd1 vssd1 vccd1 vccd1 _7842_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5130_ _8211_/Q _8195_/Q _8457_/Q _8227_/Q _5231_/S _5129_/X vssd1 vssd1 vccd1 vccd1
+ _5130_/X sky130_fd_sc_hd__mux4_2
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5061_ _5061_/A vssd1 vssd1 vccd1 vccd1 _5061_/X sky130_fd_sc_hd__buf_4
X_4012_ _4011_/X _8441_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4013_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5963_ _5963_/A _5965_/B vssd1 vssd1 vccd1 vccd1 _5964_/A sky130_fd_sc_hd__or2_1
X_4914_ _4794_/X _4912_/X _4913_/X vssd1 vssd1 vccd1 vccd1 _4914_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7702_ _7702_/A vssd1 vssd1 vccd1 vccd1 _7702_/X sky130_fd_sc_hd__buf_2
XFILLER_18_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5894_ _6672_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5895_/A sky130_fd_sc_hd__and2_1
X_4845_ _8231_/Q _4811_/X _4806_/X _8215_/Q _4760_/S vssd1 vssd1 vccd1 vccd1 _4845_/X
+ sky130_fd_sc_hd__o221a_1
X_7633_ _7633_/A _7633_/B _7633_/C _7646_/C vssd1 vssd1 vccd1 vccd1 _7634_/A sky130_fd_sc_hd__and4_1
X_4776_ _4797_/A vssd1 vssd1 vccd1 vccd1 _4806_/A sky130_fd_sc_hd__clkbuf_2
X_7564_ _8466_/Q vssd1 vssd1 vccd1 vccd1 _7564_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6515_ _6515_/A vssd1 vssd1 vccd1 vccd1 _7898_/D sky130_fd_sc_hd__clkbuf_1
X_7495_ _7670_/A vssd1 vssd1 vccd1 vccd1 _7495_/X sky130_fd_sc_hd__buf_1
XFILLER_119_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6446_ _8064_/Q vssd1 vssd1 vccd1 vccd1 _6454_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6377_ _7754_/A _6362_/X _6336_/X _6343_/X vssd1 vssd1 vccd1 vccd1 _6377_/X sky130_fd_sc_hd__a31o_1
XFILLER_114_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3089_ clkbuf_0__3089_/X vssd1 vssd1 vccd1 vccd1 _6309__210/A sky130_fd_sc_hd__clkbuf_4
X_8116_ _8116_/CLK _8116_/D vssd1 vssd1 vccd1 vccd1 _8116_/Q sky130_fd_sc_hd__dfxtp_2
X_5328_ _3911_/X _5038_/A _5327_/X _5262_/X vssd1 vssd1 vccd1 vccd1 _8125_/D sky130_fd_sc_hd__o211a_1
X_8047_ _8047_/CLK _8047_/D vssd1 vssd1 vccd1 vccd1 _8047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5259_ _5352_/B _5247_/X _5251_/X _5258_/X _5047_/A vssd1 vssd1 vccd1 vccd1 _5259_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_102_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3443_ clkbuf_0__3443_/X vssd1 vssd1 vccd1 vccd1 _7020__470/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _8188_/Q vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__inv_2
X_4561_ _4438_/X _8215_/Q _4565_/S vssd1 vssd1 vccd1 vccd1 _4562_/A sky130_fd_sc_hd__mux2_1
X_4492_ _4374_/X _8244_/Q _4500_/S vssd1 vssd1 vccd1 vccd1 _4493_/A sky130_fd_sc_hd__mux2_1
X_7280_ _7280_/A _7280_/B _7280_/C vssd1 vssd1 vccd1 vccd1 _7280_/X sky130_fd_sc_hd__and3_1
X_6231_ _6225_/X _8011_/Q _6227_/X _6229_/X _7800_/Q vssd1 vssd1 vccd1 vccd1 _7800_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6162_/A vssd1 vssd1 vccd1 vccd1 _7762_/D sky130_fd_sc_hd__clkbuf_1
X_5113_ _8409_/Q _8393_/Q _8385_/Q _8417_/Q _5284_/S _5061_/X vssd1 vssd1 vccd1 vccd1
+ _5113_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _7792_/Q _6105_/B vssd1 vssd1 vccd1 vccd1 _6093_/X sky130_fd_sc_hd__or2_1
X_5044_ _5070_/A _5070_/B vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__and2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3776_ clkbuf_0__3776_/X vssd1 vssd1 vccd1 vccd1 _7675__50/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3090_ clkbuf_0__3090_/X vssd1 vssd1 vccd1 vccd1 _6312__212/A sky130_fd_sc_hd__clkbuf_4
X_5946_ _5946_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _5947_/A sky130_fd_sc_hd__or2_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6952__418 _6952__418/A vssd1 vssd1 vccd1 vccd1 _8142_/CLK sky130_fd_sc_hd__inv_2
X_5877_ _8020_/Q _8021_/Q _8018_/Q _8019_/Q vssd1 vssd1 vccd1 vccd1 _5878_/B sky130_fd_sc_hd__and4bb_4
XFILLER_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4828_ _8337_/Q _4775_/X _8145_/Q _4777_/X _4654_/A vssd1 vssd1 vccd1 vccd1 _4828_/X
+ sky130_fd_sc_hd__o221a_1
X_7616_ _8481_/Q _7613_/X _7615_/X _7552_/X vssd1 vssd1 vccd1 vccd1 _8480_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6319__218 _6321__220/A vssd1 vssd1 vccd1 vccd1 _7848_/CLK sky130_fd_sc_hd__inv_2
X_4759_ _8147_/Q _8102_/Q _7994_/Q _8339_/Q _4868_/S _4674_/X vssd1 vssd1 vccd1 vccd1
+ _4759_/X sky130_fd_sc_hd__mux4_1
X_7547_ _7575_/A vssd1 vssd1 vccd1 vccd1 _7547_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6429_ _7865_/Q _6424_/X _6415_/X _6428_/X _6422_/X vssd1 vssd1 vccd1 vccd1 _7865_/D
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_12_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8486_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7491__23 _7493__25/A vssd1 vssd1 vccd1 vccd1 _8455_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6892__387 _6892__387/A vssd1 vssd1 vccd1 vccd1 _8101_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7111__543 _7113__545/A vssd1 vssd1 vccd1 vccd1 _8270_/CLK sky130_fd_sc_hd__inv_2
X_7164__85 _7164__85/A vssd1 vssd1 vccd1 vccd1 _8312_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _3896_/X _8448_/Q _3996_/S vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__mux2_1
X_5800_ _5800_/A vssd1 vssd1 vccd1 vccd1 _7840_/D sky130_fd_sc_hd__clkbuf_1
X_6780_ _6780_/A vssd1 vssd1 vccd1 vccd1 _6780_/X sky130_fd_sc_hd__buf_1
XFILLER_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5731_ _7918_/Q _5599_/X _5731_/S vssd1 vssd1 vccd1 vccd1 _5732_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8450_ _8450_/CLK _8450_/D vssd1 vssd1 vccd1 vccd1 _8450_/Q sky130_fd_sc_hd__dfxtp_1
X_5662_ _5677_/S vssd1 vssd1 vccd1 vccd1 _5671_/S sky130_fd_sc_hd__buf_2
X_7401_ _7432_/A vssd1 vssd1 vccd1 vccd1 _7401_/X sky130_fd_sc_hd__buf_1
X_8381_ _8381_/CLK _8381_/D vssd1 vssd1 vccd1 vccd1 _8381_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3460_ _7102_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3460_/X sky130_fd_sc_hd__clkbuf_16
X_7012__463 _7014__465/A vssd1 vssd1 vccd1 vccd1 _8190_/CLK sky130_fd_sc_hd__inv_2
X_4613_ _4613_/A vssd1 vssd1 vccd1 vccd1 _8193_/D sky130_fd_sc_hd__clkbuf_1
X_5593_ _8108_/Q vssd1 vssd1 vccd1 vccd1 _5593_/X sky130_fd_sc_hd__clkbuf_2
X_4544_ _4544_/A vssd1 vssd1 vccd1 vccd1 _8223_/D sky130_fd_sc_hd__clkbuf_1
X_7332_ _8352_/Q _7318_/X _7326_/X _7261_/B vssd1 vssd1 vccd1 vccd1 _7333_/B sky130_fd_sc_hd__o2bb2a_1
X_7263_ _7284_/B _7263_/B _7263_/C _7263_/D vssd1 vssd1 vccd1 vccd1 _7308_/B sky130_fd_sc_hd__and4_1
XFILLER_104_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4475_ _4475_/A vssd1 vssd1 vccd1 vccd1 _8250_/D sky130_fd_sc_hd__clkbuf_1
X_6214_ _6208_/X _8000_/Q _6211_/X _6213_/X _7789_/Q vssd1 vssd1 vccd1 vccd1 _7789_/D
+ sky130_fd_sc_hd__o32a_1
X_7194_ _7213_/A vssd1 vssd1 vccd1 vccd1 _7236_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6145_ _6145_/A _6151_/B vssd1 vssd1 vccd1 vccd1 _6145_/X sky130_fd_sc_hd__and2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_15 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6076_ _6114_/A vssd1 vssd1 vccd1 vccd1 _6092_/S sky130_fd_sc_hd__clkbuf_2
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_48 _6135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_26 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5027_ _4438_/X _8137_/Q _5031_/S vssd1 vssd1 vccd1 vccd1 _5028_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_37 _6129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_59 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5929_ _5929_/A vssd1 vssd1 vccd1 vccd1 _5929_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3658_ _7495_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3658_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3409_ clkbuf_0__3409_/X vssd1 vssd1 vccd1 vccd1 _6887__383/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7137__63 _7139__65/A vssd1 vssd1 vccd1 vccd1 _8290_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6530__227 _6530__227/A vssd1 vssd1 vccd1 vccd1 _7905_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ _4260_/A vssd1 vssd1 vccd1 vccd1 _8332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4191_ _8389_/Q _4190_/X _4197_/S vssd1 vssd1 vccd1 vccd1 _4192_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7950_ _7950_/CLK _7950_/D vssd1 vssd1 vccd1 vccd1 _7950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7881_ _8345_/CLK _7881_/D vssd1 vssd1 vccd1 vccd1 _7881_/Q sky130_fd_sc_hd__dfxtp_1
X_6901_ _6901_/A vssd1 vssd1 vccd1 vccd1 _8107_/D sky130_fd_sc_hd__clkbuf_1
X_7118__549 _7118__549/A vssd1 vssd1 vccd1 vccd1 _8276_/CLK sky130_fd_sc_hd__inv_2
X_6832_ _7565_/A _7565_/B _7522_/A vssd1 vssd1 vccd1 vccd1 _6832_/Y sky130_fd_sc_hd__a21oi_1
X_3975_ _8490_/Q vssd1 vssd1 vccd1 vccd1 _3975_/X sky130_fd_sc_hd__buf_2
X_6763_ _6763_/A vssd1 vssd1 vccd1 vccd1 _8064_/D sky130_fd_sc_hd__clkbuf_1
X_8502_ _8502_/CLK _8502_/D vssd1 vssd1 vccd1 vccd1 _8502_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3475_ clkbuf_0__3475_/X vssd1 vssd1 vccd1 vccd1 _7181__99/A sky130_fd_sc_hd__clkbuf_4
X_5714_ _5714_/A vssd1 vssd1 vccd1 vccd1 _7926_/D sky130_fd_sc_hd__clkbuf_1
X_6694_ _8015_/Q _5957_/A _6700_/S vssd1 vssd1 vccd1 vccd1 _6695_/A sky130_fd_sc_hd__mux2_1
X_5645_ _7956_/Q _5583_/X _5653_/S vssd1 vssd1 vccd1 vccd1 _5646_/A sky130_fd_sc_hd__mux2_1
X_8433_ _8433_/CLK _8433_/D vssd1 vssd1 vccd1 vccd1 _8433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6732__331 _6733__332/A vssd1 vssd1 vccd1 vccd1 _8041_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3443_ _7015_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3443_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5576_ _5575_/X _7990_/Q _5576_/S vssd1 vssd1 vccd1 vccd1 _5577_/A sky130_fd_sc_hd__mux2_1
X_8364_ _8368_/CLK _8364_/D vssd1 vssd1 vccd1 vccd1 _8364_/Q sky130_fd_sc_hd__dfxtp_1
X_4527_ _8230_/Q _4484_/X _4529_/S vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__mux2_1
X_8295_ _8295_/CLK _8295_/D vssd1 vssd1 vccd1 vccd1 _8295_/Q sky130_fd_sc_hd__dfxtp_1
X_7315_ _7321_/A _7315_/B vssd1 vssd1 vccd1 vccd1 _8346_/D sky130_fd_sc_hd__nor2_1
X_4458_ _4458_/A vssd1 vssd1 vccd1 vccd1 _8256_/D sky130_fd_sc_hd__clkbuf_1
X_7060__501 _7064__505/A vssd1 vssd1 vccd1 vccd1 _8228_/CLK sky130_fd_sc_hd__inv_2
X_7246_ _8550_/Q _7246_/B vssd1 vssd1 vccd1 vccd1 _7246_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_104_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7177_ _7177_/A vssd1 vssd1 vccd1 vccd1 _7177_/X sky130_fd_sc_hd__buf_1
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4389_ _4388_/X _8280_/Q _4389_/S vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__mux2_1
X_6128_ _6153_/B vssd1 vssd1 vccd1 vccd1 _6140_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6585__272 _6588__275/A vssd1 vssd1 vccd1 vccd1 _7950_/CLK sky130_fd_sc_hd__inv_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6059_ _7783_/Q _6066_/B vssd1 vssd1 vccd1 vccd1 _6059_/X sky130_fd_sc_hd__or2_1
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7453__167 _7453__167/A vssd1 vssd1 vccd1 vccd1 _8424_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7019__469 _7019__469/A vssd1 vssd1 vccd1 vccd1 _8196_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5430_ _3954_/X _8080_/Q _5438_/S vssd1 vssd1 vccd1 vccd1 _5431_/A sky130_fd_sc_hd__mux2_1
X_5361_ _5554_/A vssd1 vssd1 vccd1 vccd1 _5361_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8080_ _8080_/CLK _8080_/D vssd1 vssd1 vccd1 vccd1 _8080_/Q sky130_fd_sc_hd__dfxtp_1
X_5292_ _5230_/X _5290_/X _5291_/X vssd1 vssd1 vccd1 vccd1 _5293_/C sky130_fd_sc_hd__o21ai_1
X_4312_ _4289_/X _8312_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4243_ _4243_/A vssd1 vssd1 vccd1 vccd1 _8341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3090_ _6310_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3090_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4174_ _5482_/A _4199_/B vssd1 vssd1 vccd1 vccd1 _4197_/S sky130_fd_sc_hd__nor2_2
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7933_ _7933_/CLK _7933_/D vssd1 vssd1 vccd1 vccd1 _7933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7864_ _8550_/CLK _7864_/D vssd1 vssd1 vccd1 vccd1 _7864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7795_ _8537_/CLK _7795_/D vssd1 vssd1 vccd1 vccd1 _7795_/Q sky130_fd_sc_hd__dfxtp_1
X_6815_ _8471_/Q vssd1 vssd1 vccd1 vccd1 _6816_/A sky130_fd_sc_hd__clkinv_2
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3958_ _5805_/A vssd1 vssd1 vccd1 vccd1 _5500_/B sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3458_ clkbuf_0__3458_/X vssd1 vssd1 vccd1 vccd1 _7093__528/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3889_ _5500_/A _4567_/A vssd1 vssd1 vccd1 vccd1 _3912_/S sky130_fd_sc_hd__or2_2
X_6677_ _6677_/A vssd1 vssd1 vccd1 vccd1 _8007_/D sky130_fd_sc_hd__clkbuf_1
X_8416_ _8416_/CLK _8416_/D vssd1 vssd1 vccd1 vccd1 _8416_/Q sky130_fd_sc_hd__dfxtp_1
X_5628_ _5628_/A vssd1 vssd1 vccd1 vccd1 _7964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5559_ _5559_/A vssd1 vssd1 vccd1 vccd1 _5559_/X sky130_fd_sc_hd__clkbuf_4
X_8347_ _8370_/CLK _8347_/D vssd1 vssd1 vccd1 vccd1 _8347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7131__58 _7133__60/A vssd1 vssd1 vccd1 vccd1 _8285_/CLK sky130_fd_sc_hd__inv_2
X_8278_ _8278_/CLK _8278_/D vssd1 vssd1 vccd1 vccd1 _8278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7229_ _7319_/A _7319_/B _8546_/Q vssd1 vssd1 vccd1 vccd1 _7280_/B sky130_fd_sc_hd__a21bo_1
XFILLER_86_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6778__364 _6779__365/A vssd1 vssd1 vccd1 vccd1 _8077_/CLK sky130_fd_sc_hd__inv_2
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6739__337 _6740__338/A vssd1 vssd1 vccd1 vccd1 _8047_/CLK sky130_fd_sc_hd__inv_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6971__432 _6973__434/A vssd1 vssd1 vccd1 vccd1 _8156_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7067__507 _7070__510/A vssd1 vssd1 vccd1 vccd1 _8234_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8564__211 vssd1 vssd1 vccd1 vccd1 _8564__211/HI caravel_irq[2] sky130_fd_sc_hd__conb_1
X_7673__48 _7675__50/A vssd1 vssd1 vccd1 vccd1 _8517_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4930_ _5014_/B _5014_/C _4943_/A vssd1 vssd1 vccd1 vccd1 _4937_/B sky130_fd_sc_hd__nand3_1
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4861_ _4770_/X _4859_/X _4860_/X vssd1 vssd1 vccd1 vccd1 _4861_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4792_ _7961_/Q _7945_/Q _4866_/S vssd1 vssd1 vccd1 vccd1 _4792_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3312_ clkbuf_0__3312_/X vssd1 vssd1 vccd1 vccd1 _6746__343/A sky130_fd_sc_hd__clkbuf_4
X_7580_ _7585_/A _7580_/B vssd1 vssd1 vccd1 vccd1 _8469_/D sky130_fd_sc_hd__nor2_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6462_ _6462_/A _7502_/A _7680_/B _6938_/B vssd1 vssd1 vccd1 vccd1 _6522_/A sky130_fd_sc_hd__or4b_1
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8201_ _8201_/CLK _8201_/D vssd1 vssd1 vccd1 vccd1 _8201_/Q sky130_fd_sc_hd__dfxtp_1
X_6393_ _6331_/A _6390_/X _6392_/X _6367_/X vssd1 vssd1 vccd1 vccd1 _6393_/X sky130_fd_sc_hd__a31o_1
X_5413_ _5413_/A vssd1 vssd1 vccd1 vccd1 _8089_/D sky130_fd_sc_hd__clkbuf_1
Xoutput123 _6020_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput112 _5998_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[12] sky130_fd_sc_hd__buf_2
Xoutput134 _5987_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[7] sky130_fd_sc_hd__buf_2
X_5344_ _5344_/A vssd1 vssd1 vccd1 vccd1 _8120_/D sky130_fd_sc_hd__clkbuf_1
X_8132_ _8132_/CLK _8132_/D vssd1 vssd1 vccd1 vccd1 _8132_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput156 _5960_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[26] sky130_fd_sc_hd__buf_2
Xoutput145 _5938_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[16] sky130_fd_sc_hd__buf_2
Xoutput167 _5918_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_114_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5275_ _5193_/X _5273_/X _5274_/X vssd1 vssd1 vccd1 vccd1 _5275_/Y sky130_fd_sc_hd__o21ai_1
Xoutput178 _6084_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput189 _6121_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[20] sky130_fd_sc_hd__buf_2
X_8063_ _8063_/CLK _8063_/D vssd1 vssd1 vccd1 vccd1 _8063_/Q sky130_fd_sc_hd__dfxtp_1
X_4226_ _4226_/A vssd1 vssd1 vccd1 vccd1 _8376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4157_ _8110_/Q vssd1 vssd1 vccd1 vccd1 _4157_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4088_ _4023_/X _8414_/Q _4088_/S vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7916_ _7916_/CLK _7916_/D vssd1 vssd1 vccd1 vccd1 _7916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7847_ _7847_/CLK _7847_/D vssd1 vssd1 vccd1 vccd1 _7847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7778_ _7778_/CLK _7778_/D vssd1 vssd1 vccd1 vccd1 _7778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3409_ _6884_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3409_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3657_ clkbuf_0__3657_/X vssd1 vssd1 vccd1 vccd1 _7664_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6598__282 _6600__284/A vssd1 vssd1 vccd1 vccd1 _7960_/CLK sky130_fd_sc_hd__inv_2
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput25 caravel_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_4
Xinput14 caravel_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_4
Xinput36 wb_rst_i vssd1 vssd1 vccd1 vccd1 _6247_/A sky130_fd_sc_hd__buf_4
XFILLER_116_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput58 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_1
Xinput47 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _3866_/A sky130_fd_sc_hd__clkbuf_1
Xinput69 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5060_ _5129_/A vssd1 vssd1 vccd1 vccd1 _5061_/A sky130_fd_sc_hd__buf_2
X_4011_ _4280_/A vssd1 vssd1 vccd1 vccd1 _4011_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6978__438 _6980__440/A vssd1 vssd1 vccd1 vccd1 _8162_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5962_ _5962_/A vssd1 vssd1 vccd1 vccd1 _5962_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4913_ _8151_/Q _4768_/A _4797_/X _8090_/Q _4782_/A vssd1 vssd1 vccd1 vccd1 _4913_/X
+ sky130_fd_sc_hd__o221a_1
X_7701_ _7701_/A vssd1 vssd1 vccd1 vccd1 _7701_/X sky130_fd_sc_hd__clkbuf_2
X_5893_ _6010_/A vssd1 vssd1 vccd1 vccd1 _5975_/B sky130_fd_sc_hd__clkbuf_2
X_7410__132 _7411__133/A vssd1 vssd1 vccd1 vccd1 _8389_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4844_ _8161_/Q _8199_/Q _4873_/S vssd1 vssd1 vccd1 vccd1 _4844_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7632_ _7632_/A vssd1 vssd1 vccd1 vccd1 _8488_/D sky130_fd_sc_hd__clkbuf_1
X_4775_ _4805_/A vssd1 vssd1 vccd1 vccd1 _4775_/X sky130_fd_sc_hd__clkbuf_2
X_7563_ _7567_/A _7563_/B vssd1 vssd1 vccd1 vccd1 _8465_/D sky130_fd_sc_hd__nor2_1
X_6514_ _8013_/Q _7898_/Q _6762_/S vssd1 vssd1 vccd1 vccd1 _6515_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7494_ _7494_/A vssd1 vssd1 vccd1 vccd1 _7494_/X sky130_fd_sc_hd__buf_1
X_6445_ _7869_/Q _6442_/X _6437_/X _6444_/X _6435_/X vssd1 vssd1 vccd1 vccd1 _7869_/D
+ sky130_fd_sc_hd__a221o_1
X_6376_ _8548_/Q vssd1 vssd1 vccd1 vccd1 _7754_/A sky130_fd_sc_hd__buf_4
Xclkbuf_1_1_0__3088_ clkbuf_0__3088_/X vssd1 vssd1 vccd1 vccd1 _6299__201/A sky130_fd_sc_hd__clkbuf_4
X_8115_ _8115_/CLK _8115_/D vssd1 vssd1 vccd1 vccd1 _8115_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5327_ _8125_/Q _5041_/A _5349_/A _5326_/X _5107_/A vssd1 vssd1 vccd1 vccd1 _5327_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8046_ _8046_/CLK _8046_/D vssd1 vssd1 vccd1 vccd1 _8046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5258_ _5258_/A _5258_/B _5258_/C vssd1 vssd1 vccd1 vccd1 _5258_/X sky130_fd_sc_hd__or3_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4209_ _8382_/Q _4187_/X _4209_/S vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__mux2_1
X_5189_ _5214_/A vssd1 vssd1 vccd1 vccd1 _5207_/A sky130_fd_sc_hd__buf_2
XFILLER_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__3655_ clkbuf_0__3655_/X vssd1 vssd1 vccd1 vccd1 _7487__20/A sky130_fd_sc_hd__clkbuf_16
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4560_ _4560_/A vssd1 vssd1 vccd1 vccd1 _8216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4491_ _4506_/S vssd1 vssd1 vccd1 vccd1 _4500_/S sky130_fd_sc_hd__clkbuf_2
X_6230_ _6225_/X _8010_/Q _6227_/X _6229_/X _7799_/Q vssd1 vssd1 vccd1 vccd1 _7799_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _7737_/A _7637_/B _6161_/C vssd1 vssd1 vccd1 vccd1 _6162_/A sky130_fd_sc_hd__and3_1
XFILLER_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _3831_/X _5038_/X _5108_/X _5111_/X vssd1 vssd1 vccd1 vccd1 _8132_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _7867_/Q input7/X _6092_/S vssd1 vssd1 vccd1 vccd1 _6092_/X sky130_fd_sc_hd__mux2_1
X_6171__180 _6171__180/A vssd1 vssd1 vccd1 vccd1 _7767_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5043_ _8116_/Q _8115_/Q _8114_/Q vssd1 vssd1 vccd1 vccd1 _5070_/B sky130_fd_sc_hd__and3_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3775_ clkbuf_0__3775_/X vssd1 vssd1 vccd1 vccd1 _7669__45/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6994_ _7006_/A vssd1 vssd1 vccd1 vccd1 _6994_/X sky130_fd_sc_hd__buf_1
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5945_ _5956_/A vssd1 vssd1 vccd1 vccd1 _5954_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_43_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5876_ _5876_/A vssd1 vssd1 vccd1 vccd1 _7763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4827_ _7992_/Q _8100_/Q _4873_/S vssd1 vssd1 vccd1 vccd1 _4827_/X sky130_fd_sc_hd__mux2_1
X_7615_ _8480_/Q _7614_/X vssd1 vssd1 vccd1 vccd1 _7615_/X sky130_fd_sc_hd__or2b_1
X_4758_ _8249_/Q _8034_/Q _7986_/Q _7938_/Q _4729_/X _4674_/X vssd1 vssd1 vccd1 vccd1
+ _4758_/X sky130_fd_sc_hd__mux4_2
X_7546_ _7568_/A vssd1 vssd1 vccd1 vccd1 _7567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4689_ _6902_/A vssd1 vssd1 vccd1 vccd1 _6900_/B sky130_fd_sc_hd__buf_2
XFILLER_108_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6428_ _8540_/Q _6434_/B _6431_/C vssd1 vssd1 vccd1 vccd1 _6428_/X sky130_fd_sc_hd__and3_1
XFILLER_108_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6359_ _6350_/X _6354_/X _6356_/X _8525_/Q _6358_/X vssd1 vssd1 vccd1 vccd1 _6359_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6549__243 _6549__243/A vssd1 vssd1 vccd1 vccd1 _7921_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8029_ _8029_/CLK _8029_/D vssd1 vssd1 vccd1 vccd1 _8029_/Q sky130_fd_sc_hd__dfxtp_1
X_7417__138 _7419__140/A vssd1 vssd1 vccd1 vccd1 _8395_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7005__460 _7005__460/A vssd1 vssd1 vccd1 vccd1 _8185_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3991_ _3991_/A vssd1 vssd1 vccd1 vccd1 _8449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5730_ _5730_/A vssd1 vssd1 vccd1 vccd1 _7919_/D sky130_fd_sc_hd__clkbuf_1
X_5661_ _5661_/A _5823_/B vssd1 vssd1 vccd1 vccd1 _5677_/S sky130_fd_sc_hd__or2_2
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5592_ _5592_/A vssd1 vssd1 vccd1 vccd1 _7985_/D sky130_fd_sc_hd__clkbuf_1
X_8380_ _8380_/CLK _8380_/D vssd1 vssd1 vccd1 vccd1 _8380_/Q sky130_fd_sc_hd__dfxtp_1
X_4612_ _8193_/Q _4184_/X _4614_/S vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__mux2_1
X_4543_ _4391_/X _8223_/Q _4547_/S vssd1 vssd1 vccd1 vccd1 _4544_/A sky130_fd_sc_hd__mux2_1
X_7331_ _7336_/A _7331_/B vssd1 vssd1 vccd1 vccd1 _8351_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7262_ _7277_/B _7262_/B _7262_/C _7262_/D vssd1 vssd1 vccd1 vccd1 _7263_/D sky130_fd_sc_hd__and4_1
XFILLER_104_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4474_ _8250_/Q _4154_/X _4479_/S vssd1 vssd1 vccd1 vccd1 _4475_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6213_ _6213_/A vssd1 vssd1 vccd1 vccd1 _6213_/X sky130_fd_sc_hd__clkbuf_2
X_7193_ _8346_/Q _8345_/Q _8344_/Q _8343_/Q vssd1 vssd1 vccd1 vccd1 _7213_/A sky130_fd_sc_hd__and4_1
X_6144_ _7806_/Q _6138_/X _6139_/X _6143_/X _6136_/X vssd1 vssd1 vccd1 vccd1 _6144_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6075_ _6075_/A vssd1 vssd1 vccd1 vccd1 _6075_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_16 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5026_ _5026_/A vssd1 vssd1 vccd1 vccd1 _8138_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_27 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_49 _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_38 _6129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6325__223 _6325__223/A vssd1 vssd1 vccd1 vccd1 _7853_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5928_ _7728_/A _5932_/B vssd1 vssd1 vccd1 vccd1 _5929_/A sky130_fd_sc_hd__or2_4
X_6772__359 _6772__359/A vssd1 vssd1 vccd1 vccd1 _8072_/CLK sky130_fd_sc_hd__inv_2
X_5859_ _5859_/A _5859_/B vssd1 vssd1 vccd1 vccd1 _5875_/S sky130_fd_sc_hd__or2_2
Xclkbuf_0__3657_ _7494_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3657_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7529_ _7529_/A _7529_/B vssd1 vssd1 vccd1 vccd1 _7530_/D sky130_fd_sc_hd__xor2_1
XFILLER_119_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3408_ clkbuf_0__3408_/X vssd1 vssd1 vccd1 vccd1 _6883__380/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4190_ _8490_/Q vssd1 vssd1 vccd1 vccd1 _4190_/X sky130_fd_sc_hd__buf_2
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7880_ _8345_/CLK _7880_/D vssd1 vssd1 vccd1 vccd1 _7880_/Q sky130_fd_sc_hd__dfxtp_1
X_6900_ _8481_/Q _6900_/B vssd1 vssd1 vccd1 vccd1 _6901_/A sky130_fd_sc_hd__and2_1
X_6831_ _8465_/Q _6818_/A _8466_/Q vssd1 vssd1 vccd1 vccd1 _7565_/B sky130_fd_sc_hd__a21o_1
XINSDIODE2_120 _7201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8501_ _8501_/CLK _8501_/D vssd1 vssd1 vccd1 vccd1 _8501_/Q sky130_fd_sc_hd__dfxtp_1
X_3974_ _3974_/A vssd1 vssd1 vccd1 vccd1 _8454_/D sky130_fd_sc_hd__clkbuf_1
X_6762_ _6672_/A _6454_/C _6762_/S vssd1 vssd1 vccd1 vccd1 _6763_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3474_ clkbuf_0__3474_/X vssd1 vssd1 vccd1 vccd1 _7173__92/A sky130_fd_sc_hd__clkbuf_4
X_5713_ _7926_/Q _5599_/X _5713_/S vssd1 vssd1 vccd1 vccd1 _5714_/A sky130_fd_sc_hd__mux2_1
X_6693_ _6693_/A vssd1 vssd1 vccd1 vccd1 _8014_/D sky130_fd_sc_hd__clkbuf_1
X_5644_ _5644_/A vssd1 vssd1 vccd1 vccd1 _7957_/D sky130_fd_sc_hd__clkbuf_1
X_8432_ _8432_/CLK _8432_/D vssd1 vssd1 vccd1 vccd1 _8432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8363_ _8368_/CLK _8363_/D vssd1 vssd1 vccd1 vccd1 _8363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5575_ _5575_/A vssd1 vssd1 vccd1 vccd1 _5575_/X sky130_fd_sc_hd__clkbuf_2
X_7314_ _8346_/Q _7301_/X _7310_/X _7240_/B vssd1 vssd1 vccd1 vccd1 _7315_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4526_ _4526_/A vssd1 vssd1 vccd1 vccd1 _8231_/D sky130_fd_sc_hd__clkbuf_1
X_8294_ _8294_/CLK _8294_/D vssd1 vssd1 vccd1 vccd1 _8294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4457_ _4388_/X _8256_/Q _4457_/S vssd1 vssd1 vccd1 vccd1 _4458_/A sky130_fd_sc_hd__mux2_1
X_7245_ _8344_/Q _7302_/A vssd1 vssd1 vccd1 vccd1 _7246_/B sky130_fd_sc_hd__xor2_2
X_8581__228 vssd1 vssd1 vccd1 vccd1 _8581__228/HI manufacturerID[0] sky130_fd_sc_hd__conb_1
XFILLER_104_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4388_ _8491_/Q vssd1 vssd1 vccd1 vccd1 _4388_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6127_ _7800_/Q _6122_/X _6123_/X _6126_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6127_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6058_ _7858_/Q input29/X _6072_/S vssd1 vssd1 vccd1 vccd1 _6058_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ _5009_/A vssd1 vssd1 vccd1 vccd1 _8145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6592__277 _6594__279/A vssd1 vssd1 vccd1 vccd1 _7955_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6633__296 _6635__298/A vssd1 vssd1 vccd1 vccd1 _7982_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5360_ _8113_/Q vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5291_ _5270_/A _8074_/Q _7839_/Q _5214_/X _5092_/A vssd1 vssd1 vccd1 vccd1 _5291_/X
+ sky130_fd_sc_hd__o221a_1
X_4311_ _4311_/A vssd1 vssd1 vccd1 vccd1 _8313_/D sky130_fd_sc_hd__clkbuf_1
X_4242_ _8341_/Q _4151_/X _4248_/S vssd1 vssd1 vccd1 vccd1 _4243_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4173_ _5464_/A vssd1 vssd1 vccd1 vccd1 _5482_/A sky130_fd_sc_hd__buf_4
X_7292__109 _7293__110/A vssd1 vssd1 vccd1 vccd1 _8338_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7932_ _7932_/CLK _7932_/D vssd1 vssd1 vccd1 vccd1 _7932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7863_ _8550_/CLK _7863_/D vssd1 vssd1 vccd1 vccd1 _7863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7794_ _8537_/CLK _7794_/D vssd1 vssd1 vccd1 vccd1 _7794_/Q sky130_fd_sc_hd__dfxtp_1
X_6814_ _8537_/Q _6814_/B vssd1 vssd1 vccd1 vccd1 _6860_/B sky130_fd_sc_hd__xor2_1
XFILLER_23_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3957_ _5109_/A _5330_/A vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_1_1_0__3457_ clkbuf_0__3457_/X vssd1 vssd1 vccd1 vccd1 _7108_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8415_ _8415_/CLK _8415_/D vssd1 vssd1 vccd1 vccd1 _8415_/Q sky130_fd_sc_hd__dfxtp_1
X_6676_ _5939_/A _8007_/Q _6682_/S vssd1 vssd1 vccd1 vccd1 _6677_/A sky130_fd_sc_hd__mux2_1
X_3888_ _3956_/B _5346_/A _5109_/A vssd1 vssd1 vccd1 vccd1 _4567_/A sky130_fd_sc_hd__or3b_4
X_5627_ _5559_/X _7964_/Q _5633_/S vssd1 vssd1 vccd1 vccd1 _5628_/A sky130_fd_sc_hd__mux2_1
X_5558_ _5558_/A vssd1 vssd1 vccd1 vccd1 _7997_/D sky130_fd_sc_hd__clkbuf_1
X_8346_ _8358_/CLK _8346_/D vssd1 vssd1 vccd1 vccd1 _8346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8277_ _8277_/CLK _8277_/D vssd1 vssd1 vccd1 vccd1 _8277_/Q sky130_fd_sc_hd__dfxtp_1
X_4509_ _5622_/A vssd1 vssd1 vccd1 vccd1 _5014_/A sky130_fd_sc_hd__buf_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5489_ _5489_/A vssd1 vssd1 vccd1 vccd1 _8051_/D sky130_fd_sc_hd__clkbuf_1
X_7228_ _8347_/Q _7236_/B _7227_/A vssd1 vssd1 vccd1 vccd1 _7319_/B sky130_fd_sc_hd__a21o_1
XFILLER_59_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7159_ _7177_/A vssd1 vssd1 vccd1 vccd1 _7159_/X sky130_fd_sc_hd__buf_1
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7025__474 _7026__475/A vssd1 vssd1 vccd1 vccd1 _8201_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6600__284 _6600__284/A vssd1 vssd1 vccd1 vccd1 _7962_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8526_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4860_ _8336_/Q _4775_/X _8144_/Q _4777_/X _4654_/A vssd1 vssd1 vccd1 vccd1 _4860_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_1_0__3311_ clkbuf_0__3311_/X vssd1 vssd1 vccd1 vccd1 _6742__340/A sky130_fd_sc_hd__clkbuf_4
X_4791_ _4806_/A vssd1 vssd1 vccd1 vccd1 _4791_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6461_ _7742_/B _6461_/B _6461_/C _6461_/D vssd1 vssd1 vccd1 vccd1 _6938_/B sky130_fd_sc_hd__nor4_1
X_8200_ _8200_/CLK _8200_/D vssd1 vssd1 vccd1 vccd1 _8200_/Q sky130_fd_sc_hd__dfxtp_1
X_6392_ _8530_/Q _6356_/A _6391_/X _6397_/B _6411_/A vssd1 vssd1 vccd1 vccd1 _6392_/X
+ sky130_fd_sc_hd__a221o_1
X_5412_ _5361_/X _8089_/Q _5420_/S vssd1 vssd1 vccd1 vccd1 _5413_/A sky130_fd_sc_hd__mux2_1
Xoutput124 _6023_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput113 _6001_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[13] sky130_fd_sc_hd__buf_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5343_ _5343_/A _5343_/B _5343_/C vssd1 vssd1 vccd1 vccd1 _5344_/A sky130_fd_sc_hd__and3_1
X_8131_ _8131_/CLK _8131_/D vssd1 vssd1 vccd1 vccd1 _8131_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput157 _5962_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput135 _5990_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[8] sky130_fd_sc_hd__buf_2
Xoutput146 _5940_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[17] sky130_fd_sc_hd__buf_2
Xoutput168 _5920_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[8] sky130_fd_sc_hd__buf_2
X_5274_ _8270_/Q _5180_/X _5239_/X _8420_/Q _5250_/A vssd1 vssd1 vccd1 vccd1 _5274_/X
+ sky130_fd_sc_hd__o221a_1
Xoutput179 _6087_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[11] sky130_fd_sc_hd__buf_2
X_8062_ _8530_/CLK _8062_/D vssd1 vssd1 vccd1 vccd1 _8062_/Q sky130_fd_sc_hd__dfxtp_1
X_4225_ _8376_/Q _4154_/X _4229_/S vssd1 vssd1 vccd1 vccd1 _4226_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4156_ _4156_/A vssd1 vssd1 vccd1 vccd1 _8400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4087_ _4087_/A vssd1 vssd1 vccd1 vccd1 _8415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6543__238 _6544__239/A vssd1 vssd1 vccd1 vccd1 _7916_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7915_ _7915_/CLK _7915_/D vssd1 vssd1 vccd1 vccd1 _7915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7846_ _7846_/CLK _7846_/D vssd1 vssd1 vccd1 vccd1 _7846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7777_ _7777_/CLK _7777_/D vssd1 vssd1 vccd1 vccd1 _7777_/Q sky130_fd_sc_hd__dfxtp_1
X_4989_ _4989_/A vssd1 vssd1 vccd1 vccd1 _8154_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6659_ _6659_/A vssd1 vssd1 vccd1 vccd1 _7999_/D sky130_fd_sc_hd__clkbuf_1
X_8587__234 vssd1 vssd1 vccd1 vccd1 _8587__234/HI manufacturerID[6] sky130_fd_sc_hd__conb_1
X_8329_ _8329_/CLK _8329_/D vssd1 vssd1 vccd1 vccd1 _8329_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3408_ _6878_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3408_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3656_ clkbuf_0__3656_/X vssd1 vssd1 vccd1 vccd1 _7493__25/A sky130_fd_sc_hd__clkbuf_4
X_6745__342 _6746__343/A vssd1 vssd1 vccd1 vccd1 _8052_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7073__512 _7073__512/A vssd1 vssd1 vccd1 vccd1 _8239_/CLK sky130_fd_sc_hd__inv_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput26 caravel_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 _6149_/A sky130_fd_sc_hd__clkbuf_4
Xinput15 caravel_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_4
Xinput37 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _5971_/A sky130_fd_sc_hd__buf_4
Xinput59 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _5975_/A sky130_fd_sc_hd__buf_4
Xinput48 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _5973_/A sky130_fd_sc_hd__buf_4
X_4010_ _8494_/Q vssd1 vssd1 vccd1 vccd1 _4280_/A sky130_fd_sc_hd__buf_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _5961_/A _5965_/B vssd1 vssd1 vccd1 vccd1 _5962_/A sky130_fd_sc_hd__or2_1
XFILLER_92_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ _7910_/Q _8082_/Q _4915_/S vssd1 vssd1 vccd1 vccd1 _4912_/X sky130_fd_sc_hd__mux2_1
X_7700_ _7700_/A vssd1 vssd1 vccd1 vccd1 _7701_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5892_ _6021_/A vssd1 vssd1 vccd1 vccd1 _6010_/A sky130_fd_sc_hd__clkbuf_2
X_7631_ _7631_/A _7637_/B _7640_/C vssd1 vssd1 vccd1 vccd1 _7632_/A sky130_fd_sc_hd__and3_1
X_4843_ _4794_/X _4841_/X _4842_/X _4782_/X vssd1 vssd1 vccd1 vccd1 _4843_/X sky130_fd_sc_hd__o211a_1
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4774_ _8170_/Q vssd1 vssd1 vccd1 vccd1 _4805_/A sky130_fd_sc_hd__buf_2
X_7562_ _7561_/Y _7542_/X _7555_/X _7522_/B vssd1 vssd1 vccd1 vccd1 _7563_/B sky130_fd_sc_hd__o22a_1
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6513_ _6513_/A vssd1 vssd1 vccd1 vccd1 _7897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6444_ _7201_/A _6452_/B _6444_/C vssd1 vssd1 vccd1 vccd1 _6444_/X sky130_fd_sc_hd__and3_1
XFILLER_106_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6375_ _7856_/Q _6328_/X _6374_/X vssd1 vssd1 vccd1 vccd1 _7856_/D sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1_0__3087_ clkbuf_0__3087_/X vssd1 vssd1 vccd1 vccd1 _6322_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5326_ _5350_/B _5304_/X _5311_/X _5325_/X vssd1 vssd1 vccd1 vccd1 _5326_/X sky130_fd_sc_hd__a31o_1
X_8114_ _8114_/CLK _8114_/D vssd1 vssd1 vccd1 vccd1 _8114_/Q sky130_fd_sc_hd__dfxtp_2
X_8045_ _8045_/CLK _8045_/D vssd1 vssd1 vccd1 vccd1 _8045_/Q sky130_fd_sc_hd__dfxtp_1
X_5257_ _5244_/A _5255_/X _5256_/X vssd1 vssd1 vccd1 vccd1 _5258_/C sky130_fd_sc_hd__o21a_1
X_4208_ _4208_/A vssd1 vssd1 vccd1 vccd1 _8383_/D sky130_fd_sc_hd__clkbuf_1
X_5188_ _5197_/A vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0__3441_ clkbuf_0__3441_/X vssd1 vssd1 vccd1 vccd1 _7011__462/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4139_ _4217_/A _8173_/Q vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7829_ _7829_/CLK _7829_/D vssd1 vssd1 vccd1 vccd1 _7829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7176__95 _7176__95/A vssd1 vssd1 vccd1 vccd1 _8322_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8561__259 vssd1 vssd1 vccd1 vccd1 partID[15] _8561__259/LO sky130_fd_sc_hd__conb_1
Xclkbuf_1_0_0__3639_ clkbuf_0__3639_/X vssd1 vssd1 vccd1 vccd1 _7426_/A sky130_fd_sc_hd__clkbuf_4
X_7651__30 _7651__30/A vssd1 vssd1 vccd1 vccd1 _8499_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7038__484 _7038__484/A vssd1 vssd1 vccd1 vccd1 _8211_/CLK sky130_fd_sc_hd__inv_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4490_ _4490_/A _5805_/A vssd1 vssd1 vccd1 vccd1 _4506_/S sky130_fd_sc_hd__or2_2
XFILLER_7_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6984__443 _6986__445/A vssd1 vssd1 vccd1 vccd1 _8168_/CLK sky130_fd_sc_hd__inv_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _7689_/A vssd1 vssd1 vccd1 vccd1 _7737_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5343_/A vssd1 vssd1 vccd1 vccd1 _5111_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6075_/X _6088_/X _6090_/X _6083_/X vssd1 vssd1 vccd1 vccd1 _6091_/X sky130_fd_sc_hd__o211a_1
XFILLER_97_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5042_ _5176_/A vssd1 vssd1 vccd1 vccd1 _5348_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3774_ clkbuf_0__3774_/X vssd1 vssd1 vccd1 vccd1 _7660__37/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6993_ _7058_/A vssd1 vssd1 vccd1 vccd1 _6993_/X sky130_fd_sc_hd__buf_1
X_5944_ _5944_/A vssd1 vssd1 vccd1 vccd1 _5944_/X sky130_fd_sc_hd__clkbuf_1
X_5875_ _4169_/X _7763_/Q _5875_/S vssd1 vssd1 vccd1 vccd1 _5876_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7614_ _7614_/A vssd1 vssd1 vccd1 vccd1 _7614_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4826_ _4435_/X _4629_/X _4825_/X _4690_/X vssd1 vssd1 vccd1 vccd1 _8182_/D sky130_fd_sc_hd__o211a_1
X_7545_ _7505_/A _7539_/C _7544_/Y vssd1 vssd1 vccd1 vccd1 _8460_/D sky130_fd_sc_hd__a21oi_1
X_4757_ _4739_/S _4756_/X _4886_/A vssd1 vssd1 vccd1 vccd1 _4757_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7476_ _7482_/A vssd1 vssd1 vccd1 vccd1 _7476_/X sky130_fd_sc_hd__buf_1
X_4688_ _4713_/A _8186_/Q _4947_/A _4686_/X _4712_/A vssd1 vssd1 vccd1 vccd1 _4688_/X
+ sky130_fd_sc_hd__a221o_1
X_6427_ _7864_/Q _6424_/X _6415_/X _6426_/X _6422_/X vssd1 vssd1 vccd1 vccd1 _7864_/D
+ sky130_fd_sc_hd__a221o_1
X_6358_ _6411_/A vssd1 vssd1 vccd1 vccd1 _6358_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5309_ _8269_/Q _5232_/X _5198_/X _8419_/Q vssd1 vssd1 vccd1 vccd1 _5309_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8028_ _8028_/CLK _8028_/D vssd1 vssd1 vccd1 vccd1 _8028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3424_ clkbuf_0__3424_/X vssd1 vssd1 vccd1 vccd1 _6937__410/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _8543_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7149__73 _7149__73/A vssd1 vssd1 vccd1 vccd1 _8300_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3990_ _3893_/X _8449_/Q _3996_/S vssd1 vssd1 vccd1 vccd1 _3991_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _5660_/A vssd1 vssd1 vccd1 vccd1 _7950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4611_ _4611_/A vssd1 vssd1 vccd1 vccd1 _8194_/D sky130_fd_sc_hd__clkbuf_1
X_5591_ _7985_/Q _5590_/X _5591_/S vssd1 vssd1 vccd1 vccd1 _5592_/A sky130_fd_sc_hd__mux2_1
X_4542_ _4542_/A vssd1 vssd1 vccd1 vccd1 _8224_/D sky130_fd_sc_hd__clkbuf_1
X_7330_ _8351_/Q _7318_/X _7326_/X _7329_/Y vssd1 vssd1 vccd1 vccd1 _7331_/B sky130_fd_sc_hd__o2bb2a_1
X_4473_ _4473_/A vssd1 vssd1 vccd1 vccd1 _8251_/D sky130_fd_sc_hd__clkbuf_1
X_7261_ _8542_/Q _7261_/B vssd1 vssd1 vccd1 vccd1 _7262_/D sky130_fd_sc_hd__xor2_1
X_6869__369 _6870__370/A vssd1 vssd1 vccd1 vccd1 _8083_/CLK sky130_fd_sc_hd__inv_2
X_6212_ _6208_/X _7999_/Q _6211_/X _6204_/X _7788_/Q vssd1 vssd1 vccd1 vccd1 _7788_/D
+ sky130_fd_sc_hd__o32a_1
X_7192_ _8361_/Q _8360_/Q _7356_/B _7298_/A vssd1 vssd1 vccd1 vccd1 _7350_/B sky130_fd_sc_hd__and4_1
X_6143_ _6143_/A _6151_/B vssd1 vssd1 vccd1 vccd1 _6143_/X sky130_fd_sc_hd__and2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6074_ _6056_/X _6072_/X _6073_/X _6063_/X vssd1 vssd1 vccd1 vccd1 _6074_/X sky130_fd_sc_hd__o211a_1
XFILLER_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_39 _6129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ _4435_/X _8138_/Q _5025_/S vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_17 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_28 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5927_ _5927_/A vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5858_ _5858_/A vssd1 vssd1 vccd1 vccd1 _7771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5789_ _7845_/Q _4275_/A _5797_/S vssd1 vssd1 vccd1 vccd1 _5790_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3656_ _7488_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3656_/X sky130_fd_sc_hd__clkbuf_16
X_4809_ _4809_/A vssd1 vssd1 vccd1 vccd1 _4955_/B sky130_fd_sc_hd__buf_2
XFILLER_119_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7528_ _7528_/A _7528_/B vssd1 vssd1 vccd1 vccd1 _7530_/C sky130_fd_sc_hd__or2_1
X_7423__143 _7425__145/A vssd1 vssd1 vccd1 vccd1 _8400_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3407_ clkbuf_0__3407_/X vssd1 vssd1 vccd1 vccd1 _6919_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3269_ clkbuf_0__3269_/X vssd1 vssd1 vccd1 vccd1 _6628__292/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6645__305 _6645__305/A vssd1 vssd1 vccd1 vccd1 _7991_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_110 _7640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6830_ _6830_/A _6830_/B vssd1 vssd1 vccd1 vccd1 _7565_/A sky130_fd_sc_hd__nand2_2
XINSDIODE2_121 _6269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6761_ _6761_/A vssd1 vssd1 vccd1 vccd1 _8063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8500_ _8500_/CLK _8500_/D vssd1 vssd1 vccd1 vccd1 _8500_/Q sky130_fd_sc_hd__dfxtp_1
X_5712_ _5712_/A vssd1 vssd1 vccd1 vccd1 _7927_/D sky130_fd_sc_hd__clkbuf_1
X_3973_ _8454_/Q _3972_/X _3973_/S vssd1 vssd1 vccd1 vccd1 _3974_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3473_ clkbuf_0__3473_/X vssd1 vssd1 vccd1 vccd1 _7170__90/A sky130_fd_sc_hd__clkbuf_4
X_6692_ _8014_/Q _5954_/A _6700_/S vssd1 vssd1 vccd1 vccd1 _6693_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5643_ _7957_/Q _5578_/X _5653_/S vssd1 vssd1 vccd1 vccd1 _5644_/A sky130_fd_sc_hd__mux2_1
X_8431_ _8431_/CLK _8431_/D vssd1 vssd1 vccd1 vccd1 _8431_/Q sky130_fd_sc_hd__dfxtp_1
X_5574_ _5574_/A vssd1 vssd1 vccd1 vccd1 _7991_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3441_ _7006_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3441_/X sky130_fd_sc_hd__clkbuf_16
X_8362_ _8368_/CLK _8362_/D vssd1 vssd1 vccd1 vccd1 _8362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4525_ _8231_/Q _4481_/X _4529_/S vssd1 vssd1 vccd1 vccd1 _4526_/A sky130_fd_sc_hd__mux2_1
X_7313_ _7321_/A _7313_/B vssd1 vssd1 vccd1 vccd1 _8345_/D sky130_fd_sc_hd__nor2_1
XFILLER_117_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8293_ _8293_/CLK _8293_/D vssd1 vssd1 vccd1 vccd1 _8293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7143__68 _7145__70/A vssd1 vssd1 vccd1 vccd1 _8295_/CLK sky130_fd_sc_hd__inv_2
X_4456_ _4456_/A vssd1 vssd1 vccd1 vccd1 _8257_/D sky130_fd_sc_hd__clkbuf_1
X_7244_ _8343_/Q vssd1 vssd1 vccd1 vccd1 _7302_/A sky130_fd_sc_hd__clkbuf_2
X_4387_ _4387_/A vssd1 vssd1 vccd1 vccd1 _8281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6126_ _6139_/A vssd1 vssd1 vccd1 vccd1 _6126_/X sky130_fd_sc_hd__clkbuf_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6057_ _6114_/A vssd1 vssd1 vccd1 vccd1 _6072_/S sky130_fd_sc_hd__buf_2
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6288__193 _6290__195/A vssd1 vssd1 vccd1 vccd1 _7823_/CLK sky130_fd_sc_hd__inv_2
X_5008_ _8145_/Q _4481_/X _5012_/S vssd1 vssd1 vccd1 vccd1 _5009_/A sky130_fd_sc_hd__mux2_1
X_6997__453 _6998__454/A vssd1 vssd1 vccd1 vccd1 _8178_/CLK sky130_fd_sc_hd__inv_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3639_ _7401_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3639_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_6_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6709__313 _6711__315/A vssd1 vssd1 vccd1 vccd1 _8023_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5290_ _8326_/Q _8047_/Q _5290_/S vssd1 vssd1 vccd1 vccd1 _5290_/X sky130_fd_sc_hd__mux2_1
X_4310_ _4286_/X _8313_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4311_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4241_ _4241_/A vssd1 vssd1 vccd1 vccd1 _8342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4172_ _8495_/Q vssd1 vssd1 vccd1 vccd1 _4172_/X sky130_fd_sc_hd__buf_2
XFILLER_83_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7931_ _7931_/CLK _7931_/D vssd1 vssd1 vccd1 vccd1 _7931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7862_ _8063_/CLK _7862_/D vssd1 vssd1 vccd1 vccd1 _7862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7793_ _8537_/CLK _7793_/D vssd1 vssd1 vccd1 vccd1 _7793_/Q sky130_fd_sc_hd__dfxtp_1
X_6813_ _7532_/B _7532_/C vssd1 vssd1 vccd1 vccd1 _6814_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3956_ _8133_/Q _3956_/B _4038_/A _5335_/A vssd1 vssd1 vccd1 vccd1 _5330_/A sky130_fd_sc_hd__and4_1
Xclkbuf_1_1_0__3456_ clkbuf_0__3456_/X vssd1 vssd1 vccd1 vccd1 _7087__524/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6675_ _6675_/A vssd1 vssd1 vccd1 vccd1 _8006_/D sky130_fd_sc_hd__clkbuf_1
X_5626_ _5626_/A vssd1 vssd1 vccd1 vccd1 _7965_/D sky130_fd_sc_hd__clkbuf_1
X_8414_ _8414_/CLK _8414_/D vssd1 vssd1 vccd1 vccd1 _8414_/Q sky130_fd_sc_hd__dfxtp_1
X_3887_ _3873_/X _3886_/Y _6247_/A vssd1 vssd1 vccd1 vccd1 _5109_/A sky130_fd_sc_hd__a21oi_4
X_5557_ _5554_/X _7997_/Q _5567_/S vssd1 vssd1 vccd1 vccd1 _5558_/A sky130_fd_sc_hd__mux2_1
X_8345_ _8345_/CLK _8345_/D vssd1 vssd1 vccd1 vccd1 _8345_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3424_ _6932_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3424_/X sky130_fd_sc_hd__clkbuf_16
X_5488_ _8051_/Q _4283_/A _5492_/S vssd1 vssd1 vccd1 vccd1 _5489_/A sky130_fd_sc_hd__mux2_1
X_8276_ _8276_/CLK _8276_/D vssd1 vssd1 vccd1 vccd1 _8276_/Q sky130_fd_sc_hd__dfxtp_1
X_4508_ _8175_/Q vssd1 vssd1 vccd1 vccd1 _5014_/C sky130_fd_sc_hd__buf_2
X_4439_ _4438_/X _8263_/Q _4445_/S vssd1 vssd1 vccd1 vccd1 _4440_/A sky130_fd_sc_hd__mux2_1
X_7227_ _7227_/A _7236_/A _7232_/B vssd1 vssd1 vccd1 vccd1 _7319_/A sky130_fd_sc_hd__nand3_1
XFILLER_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7089_ _7089_/A vssd1 vssd1 vccd1 vccd1 _7089_/X sky130_fd_sc_hd__buf_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _7796_/Q _6122_/A vssd1 vssd1 vccd1 vccd1 _6109_/X sky130_fd_sc_hd__or2_1
XFILLER_100_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7032__479 _7033__480/A vssd1 vssd1 vccd1 vccd1 _8206_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7436__153 _7436__153/A vssd1 vssd1 vccd1 vccd1 _8410_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4790_ _7929_/Q _4658_/B _4784_/X vssd1 vssd1 vccd1 vccd1 _4790_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1_0__3310_ clkbuf_0__3310_/X vssd1 vssd1 vccd1 vccd1 _6736__335/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6460_ _8534_/Q vssd1 vssd1 vccd1 vccd1 _7502_/A sky130_fd_sc_hd__inv_2
X_5411_ _5426_/S vssd1 vssd1 vccd1 vccd1 _5420_/S sky130_fd_sc_hd__buf_2
X_6391_ _7741_/A _7971_/Q _6352_/X _6364_/X vssd1 vssd1 vccd1 vccd1 _6391_/X sky130_fd_sc_hd__a31o_1
Xoutput125 _6025_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[24] sky130_fd_sc_hd__buf_2
Xoutput114 _6003_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[14] sky130_fd_sc_hd__buf_2
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5342_ _5106_/A _4038_/A _7680_/B _3956_/B vssd1 vssd1 vccd1 vccd1 _5343_/C sky130_fd_sc_hd__a31o_1
X_8130_ _8130_/CLK _8130_/D vssd1 vssd1 vccd1 vccd1 _8130_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput136 _5992_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[9] sky130_fd_sc_hd__buf_2
Xoutput158 _5964_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[28] sky130_fd_sc_hd__buf_2
Xoutput147 _5942_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[18] sky130_fd_sc_hd__buf_2
XFILLER_99_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8061_ _8061_/CLK _8061_/D vssd1 vssd1 vccd1 vccd1 _8061_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput169 _5922_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5273_ _8318_/Q _8055_/Q _5273_/S vssd1 vssd1 vccd1 vccd1 _5273_/X sky130_fd_sc_hd__mux2_1
X_4224_ _4224_/A vssd1 vssd1 vccd1 vccd1 _8377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4155_ _8400_/Q _4154_/X _4161_/S vssd1 vssd1 vccd1 vccd1 _4156_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4086_ _4019_/X _8415_/Q _4088_/S vssd1 vssd1 vccd1 vccd1 _4087_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7914_ _7914_/CLK _7914_/D vssd1 vssd1 vccd1 vccd1 _7914_/Q sky130_fd_sc_hd__dfxtp_1
X_7845_ _7845_/CLK _7845_/D vssd1 vssd1 vccd1 vccd1 _7845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7776_ _7776_/CLK _7776_/D vssd1 vssd1 vccd1 vccd1 _7776_/Q sky130_fd_sc_hd__dfxtp_1
X_4988_ _8154_/Q _4478_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__mux2_1
X_3939_ _3939_/A vssd1 vssd1 vccd1 vccd1 _8503_/D sky130_fd_sc_hd__clkbuf_1
X_6658_ _5921_/A _7999_/Q _6664_/S vssd1 vssd1 vccd1 vccd1 _6659_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3439_ clkbuf_0__3439_/X vssd1 vssd1 vccd1 vccd1 _6999__455/A sky130_fd_sc_hd__clkbuf_4
X_5609_ _5608_/X _7979_/Q _5614_/S vssd1 vssd1 vccd1 vccd1 _5610_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6589_ _6589_/A vssd1 vssd1 vccd1 vccd1 _6589_/X sky130_fd_sc_hd__buf_1
X_8328_ _8328_/CLK _8328_/D vssd1 vssd1 vccd1 vccd1 _8328_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3407_ _6877_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3407_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8259_ _8259_/CLK _8259_/D vssd1 vssd1 vccd1 vccd1 _8259_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3269_ _6626_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3269_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_86_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput27 caravel_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 _6151_/A sky130_fd_sc_hd__clkbuf_4
Xinput16 caravel_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 _6123_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput38 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 _5993_/A sky130_fd_sc_hd__buf_4
Xinput49 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _3866_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5960_ _5960_/A vssd1 vssd1 vccd1 vccd1 _5960_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5891_ _5891_/A vssd1 vssd1 vccd1 vccd1 _5891_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ _4955_/B _4909_/X _4910_/X vssd1 vssd1 vccd1 vccd1 _4911_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7630_ _7613_/A _7499_/X _7629_/X _7543_/X vssd1 vssd1 vccd1 vccd1 _8487_/D sky130_fd_sc_hd__o211a_1
X_4842_ _8397_/Q _4805_/Y _4806_/X _8373_/Q vssd1 vssd1 vccd1 vccd1 _4842_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4773_ _7993_/Q _8101_/Q _4873_/S vssd1 vssd1 vccd1 vccd1 _4773_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7561_ _8465_/Q vssd1 vssd1 vccd1 vccd1 _7561_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6512_ _8012_/Q _7897_/Q _6762_/S vssd1 vssd1 vccd1 vccd1 _6513_/A sky130_fd_sc_hd__mux2_1
X_6443_ _8536_/Q vssd1 vssd1 vccd1 vccd1 _7201_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6374_ _6331_/A _6371_/X _6373_/X _6367_/X vssd1 vssd1 vccd1 vccd1 _6374_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_1_1_0__3086_ clkbuf_0__3086_/X vssd1 vssd1 vccd1 vccd1 _6294__198/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5325_ _5235_/A _5314_/X _5317_/X _5324_/X _5047_/A vssd1 vssd1 vccd1 vccd1 _5325_/X
+ sky130_fd_sc_hd__o311a_1
X_8113_ _8531_/CLK _8113_/D vssd1 vssd1 vccd1 vccd1 _8113_/Q sky130_fd_sc_hd__dfxtp_4
X_8044_ _8044_/CLK _8044_/D vssd1 vssd1 vccd1 vccd1 _8044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5256_ _8413_/Q _5227_/A _5214_/A _8405_/Q _5091_/A vssd1 vssd1 vccd1 vccd1 _5256_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4207_ _8383_/Q _4184_/X _4209_/S vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3440_ clkbuf_0__3440_/X vssd1 vssd1 vccd1 vccd1 _7005__460/A sky130_fd_sc_hd__clkbuf_4
X_5187_ _8240_/Q _8256_/Q _5312_/S vssd1 vssd1 vccd1 vccd1 _5187_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4138_ _4622_/B _4135_/Y _4137_/X vssd1 vssd1 vccd1 vccd1 _4138_/Y sky130_fd_sc_hd__a21oi_1
X_4069_ _4069_/A vssd1 vssd1 vccd1 vccd1 _8422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7828_ _7828_/CLK _7828_/D vssd1 vssd1 vccd1 vccd1 _7828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7759_ _8550_/Q _7747_/Y _7758_/X vssd1 vssd1 vccd1 vccd1 _8550_/D sky130_fd_sc_hd__a21o_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3638_ clkbuf_0__3638_/X vssd1 vssd1 vccd1 vccd1 _7399__124/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _7791_/Q _6105_/B vssd1 vssd1 vccd1 vccd1 _6090_/X sky130_fd_sc_hd__or2_1
X_5110_ _6941_/B vssd1 vssd1 vccd1 vccd1 _5343_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A _7363_/A vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__nor2_1
XFILLER_97_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3773_ clkbuf_0__3773_/X vssd1 vssd1 vccd1 vccd1 _7656__34/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5943_ _5943_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5944_/A sky130_fd_sc_hd__or2_1
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5874_ _5874_/A vssd1 vssd1 vccd1 vccd1 _7764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7613_ _7613_/A vssd1 vssd1 vccd1 vccd1 _7613_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4825_ _4713_/X _8182_/Q _4712_/X _4824_/X vssd1 vssd1 vccd1 vccd1 _4825_/X sky130_fd_sc_hd__a211o_1
X_7544_ _7503_/C _7542_/X _7543_/X vssd1 vssd1 vccd1 vccd1 _7544_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4756_ _7767_/Q _7775_/Q _7850_/Q _7954_/Q _4729_/X _4716_/A vssd1 vssd1 vccd1 vccd1
+ _4756_/X sky130_fd_sc_hd__mux4_2
X_4687_ _8187_/Q _6605_/B vssd1 vssd1 vccd1 vccd1 _4712_/A sky130_fd_sc_hd__and2_1
XFILLER_104_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6426_ _7529_/A _6434_/B _6431_/C vssd1 vssd1 vccd1 vccd1 _6426_/X sky130_fd_sc_hd__and3_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6357_ _7742_/C _6398_/B vssd1 vssd1 vccd1 vccd1 _6411_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5308_ _8317_/Q _8054_/Q _5308_/S vssd1 vssd1 vccd1 vccd1 _5308_/X sky130_fd_sc_hd__mux2_1
X_5239_ _5319_/B vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8027_ _8027_/CLK _8027_/D vssd1 vssd1 vccd1 vccd1 _8027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3423_ clkbuf_0__3423_/X vssd1 vssd1 vccd1 vccd1 _6931__405/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6556__249 _6557__250/A vssd1 vssd1 vccd1 vccd1 _7927_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4610_ _8194_/Q _4181_/X _4614_/S vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5590_ _8109_/Q vssd1 vssd1 vccd1 vccd1 _5590_/X sky130_fd_sc_hd__buf_2
XFILLER_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7086__523 _7087__524/A vssd1 vssd1 vccd1 vccd1 _8250_/CLK sky130_fd_sc_hd__inv_2
X_4541_ _4388_/X _8224_/Q _4541_/S vssd1 vssd1 vccd1 vccd1 _4542_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4472_ _8251_/Q _4471_/X _4479_/S vssd1 vssd1 vccd1 vccd1 _4473_/A sky130_fd_sc_hd__mux2_1
X_7155__77 _7158__80/A vssd1 vssd1 vccd1 vccd1 _8304_/CLK sky130_fd_sc_hd__inv_2
X_7260_ _7210_/A _7210_/B _7218_/D _7329_/A _7259_/Y vssd1 vssd1 vccd1 vccd1 _7261_/B
+ sky130_fd_sc_hd__a32o_2
X_6211_ _6272_/A vssd1 vssd1 vccd1 vccd1 _6211_/X sky130_fd_sc_hd__clkbuf_2
X_7191_ _7385_/S vssd1 vssd1 vccd1 vccd1 _7286_/A sky130_fd_sc_hd__clkbuf_2
X_6142_ _6153_/B vssd1 vssd1 vccd1 vccd1 _6151_/B sky130_fd_sc_hd__clkbuf_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6073_ _7787_/Q _6086_/B vssd1 vssd1 vccd1 vccd1 _6073_/X sky130_fd_sc_hd__or2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_29 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_18 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5024_ _5024_/A vssd1 vssd1 vccd1 vccd1 _8139_/D sky130_fd_sc_hd__clkbuf_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6975_ _6975_/A vssd1 vssd1 vccd1 vccd1 _6975_/X sky130_fd_sc_hd__buf_1
XFILLER_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5926_ _5926_/A _5932_/B vssd1 vssd1 vccd1 vccd1 _5927_/A sky130_fd_sc_hd__or2_4
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5857_ _4169_/X _7771_/Q _5857_/S vssd1 vssd1 vccd1 vccd1 _5858_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5788_ _5803_/S vssd1 vssd1 vccd1 vccd1 _5797_/S sky130_fd_sc_hd__buf_2
Xclkbuf_0__3655_ _7482_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3655_/X sky130_fd_sc_hd__clkbuf_16
X_4808_ _4803_/X _4804_/X _4807_/X _4782_/X vssd1 vssd1 vccd1 vccd1 _4808_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4739_ _4736_/X _4738_/X _4739_/S vssd1 vssd1 vccd1 vccd1 _4739_/X sky130_fd_sc_hd__mux2_1
X_7527_ _7528_/A _7528_/B vssd1 vssd1 vccd1 vccd1 _7530_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6409_ _8543_/Q vssd1 vssd1 vccd1 vccd1 _6854_/A sky130_fd_sc_hd__clkbuf_4
X_7389_ _7389_/A vssd1 vssd1 vccd1 vccd1 _7389_/X sky130_fd_sc_hd__buf_1
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3406_ clkbuf_0__3406_/X vssd1 vssd1 vccd1 vccd1 _6876__375/A sky130_fd_sc_hd__clkbuf_4
X_6562__253 _6563__254/A vssd1 vssd1 vccd1 vccd1 _7931_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_111 _3896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_100 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_122 _7631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6760_ _6654_/A _6431_/C _6762_/S vssd1 vssd1 vccd1 vccd1 _6761_/A sky130_fd_sc_hd__mux2_1
X_5711_ _7927_/Q _5596_/X _5713_/S vssd1 vssd1 vccd1 vccd1 _5712_/A sky130_fd_sc_hd__mux2_1
X_3972_ _8491_/Q vssd1 vssd1 vccd1 vccd1 _3972_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3472_ clkbuf_0__3472_/X vssd1 vssd1 vccd1 vccd1 _7163__84/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6875__374 _6876__375/A vssd1 vssd1 vccd1 vccd1 _8088_/CLK sky130_fd_sc_hd__inv_2
X_6691_ _6706_/S vssd1 vssd1 vccd1 vccd1 _6700_/S sky130_fd_sc_hd__clkbuf_2
X_8430_ _8430_/CLK _8430_/D vssd1 vssd1 vccd1 vccd1 _8430_/Q sky130_fd_sc_hd__dfxtp_1
X_5642_ _5659_/S vssd1 vssd1 vccd1 vccd1 _5653_/S sky130_fd_sc_hd__buf_2
X_5573_ _5572_/X _7991_/Q _5576_/S vssd1 vssd1 vccd1 vccd1 _5574_/A sky130_fd_sc_hd__mux2_1
X_6916__393 _6918__395/A vssd1 vssd1 vccd1 vccd1 _8115_/CLK sky130_fd_sc_hd__inv_2
X_8361_ _8370_/CLK _8361_/D vssd1 vssd1 vccd1 vccd1 _8361_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3440_ _7000_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3440_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4524_ _4524_/A vssd1 vssd1 vccd1 vccd1 _8232_/D sky130_fd_sc_hd__clkbuf_1
X_7312_ _8345_/Q _7301_/X _7310_/X _7311_/Y vssd1 vssd1 vccd1 vccd1 _7313_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8292_ _8292_/CLK _8292_/D vssd1 vssd1 vccd1 vccd1 _8292_/Q sky130_fd_sc_hd__dfxtp_1
X_4455_ _4385_/X _8257_/Q _4457_/S vssd1 vssd1 vccd1 vccd1 _4456_/A sky130_fd_sc_hd__mux2_1
X_7243_ _7311_/A _7311_/B _6838_/A vssd1 vssd1 vccd1 vccd1 _7243_/Y sky130_fd_sc_hd__a21oi_1
X_4386_ _4385_/X _8281_/Q _4389_/S vssd1 vssd1 vccd1 vccd1 _4387_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6125_ _7875_/Q _6161_/C _7731_/A vssd1 vssd1 vccd1 vccd1 _6139_/A sky130_fd_sc_hd__a21bo_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6056_ _6075_/A vssd1 vssd1 vccd1 vccd1 _6056_/X sky130_fd_sc_hd__clkbuf_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5007_ _5007_/A vssd1 vssd1 vccd1 vccd1 _8146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5909_ _5909_/A vssd1 vssd1 vccd1 vccd1 _5909_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3638_ _7395_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3638_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_6_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6651__310 _6651__310/A vssd1 vssd1 vccd1 vccd1 _7996_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4240_ _8342_/Q _4114_/X _4248_/S vssd1 vssd1 vccd1 vccd1 _4241_/A sky130_fd_sc_hd__mux2_1
X_4171_ _4171_/A vssd1 vssd1 vccd1 vccd1 _8395_/D sky130_fd_sc_hd__clkbuf_1
X_6569__259 _6570__260/A vssd1 vssd1 vccd1 vccd1 _7937_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7930_ _7930_/CLK _7930_/D vssd1 vssd1 vccd1 vccd1 _7930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7861_ _8063_/CLK _7861_/D vssd1 vssd1 vccd1 vccd1 _7861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6812_ _6812_/A _6812_/B _6857_/D vssd1 vssd1 vccd1 vccd1 _7532_/C sky130_fd_sc_hd__or3b_4
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7792_ _8540_/CLK _7792_/D vssd1 vssd1 vccd1 vccd1 _7792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6743_ _6749_/A vssd1 vssd1 vccd1 vccd1 _6743_/X sky130_fd_sc_hd__buf_1
X_3955_ _4256_/A _5334_/A _4256_/C vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__nand3b_4
XFILLER_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3455_ clkbuf_0__3455_/X vssd1 vssd1 vccd1 vccd1 _7082__520/A sky130_fd_sc_hd__clkbuf_4
X_6674_ _5937_/A _8006_/Q _6682_/S vssd1 vssd1 vccd1 vccd1 _6675_/A sky130_fd_sc_hd__mux2_1
X_5625_ _5554_/X _7965_/Q _5633_/S vssd1 vssd1 vccd1 vccd1 _5626_/A sky130_fd_sc_hd__mux2_1
X_8413_ _8413_/CLK _8413_/D vssd1 vssd1 vccd1 vccd1 _8413_/Q sky130_fd_sc_hd__dfxtp_1
X_3886_ _6398_/A _6461_/B _6461_/C vssd1 vssd1 vccd1 vccd1 _3886_/Y sky130_fd_sc_hd__nor3_1
X_5556_ _5576_/S vssd1 vssd1 vccd1 vccd1 _5567_/S sky130_fd_sc_hd__clkbuf_2
X_8344_ _8370_/CLK _8344_/D vssd1 vssd1 vccd1 vccd1 _8344_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__3423_ _6926_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3423_/X sky130_fd_sc_hd__clkbuf_16
X_5487_ _5487_/A vssd1 vssd1 vccd1 vccd1 _8052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8275_ _8275_/CLK _8275_/D vssd1 vssd1 vccd1 vccd1 _8275_/Q sky130_fd_sc_hd__dfxtp_1
X_4507_ _4507_/A vssd1 vssd1 vccd1 vccd1 _8237_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4438_ _8108_/Q vssd1 vssd1 vccd1 vccd1 _4438_/X sky130_fd_sc_hd__buf_2
X_7226_ _7323_/A _7323_/B _7510_/A vssd1 vssd1 vccd1 vccd1 _7281_/A sky130_fd_sc_hd__a21o_1
XFILLER_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4369_ _4369_/A vssd1 vssd1 vccd1 vccd1 _8287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7099__533 _7099__533/A vssd1 vssd1 vccd1 vccd1 _8260_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ _6108_/A vssd1 vssd1 vccd1 vccd1 _6122_/A sky130_fd_sc_hd__clkbuf_2
X_6039_ _7854_/Q input3/X _6123_/B vssd1 vssd1 vccd1 vccd1 _6039_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8571__218 vssd1 vssd1 vccd1 vccd1 _8571__218/HI core0Index[5] sky130_fd_sc_hd__conb_1
Xclkbuf_1_0__f__3463_ clkbuf_0__3463_/X vssd1 vssd1 vccd1 vccd1 _7152_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5410_ _5661_/A _5733_/B vssd1 vssd1 vccd1 vccd1 _5426_/S sky130_fd_sc_hd__or2_2
X_6948__415 _6948__415/A vssd1 vssd1 vccd1 vccd1 _8139_/CLK sky130_fd_sc_hd__inv_2
X_6390_ _7522_/A _6362_/X _6410_/C _6397_/A vssd1 vssd1 vccd1 vccd1 _6390_/X sky130_fd_sc_hd__a31o_1
Xoutput115 _6005_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[15] sky130_fd_sc_hd__buf_2
X_5341_ _5334_/B _5334_/C _5340_/Y vssd1 vssd1 vccd1 vccd1 _8121_/D sky130_fd_sc_hd__a21oi_1
Xoutput126 _6027_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[25] sky130_fd_sc_hd__buf_2
Xoutput137 _5890_/B vssd1 vssd1 vccd1 vccd1 caravel_wb_cyc_o sky130_fd_sc_hd__buf_2
Xoutput159 _5966_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[29] sky130_fd_sc_hd__buf_2
Xoutput148 _5944_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[19] sky130_fd_sc_hd__buf_2
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8060_ _8060_/CLK _8060_/D vssd1 vssd1 vccd1 vccd1 _8060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5272_ _5356_/B _5269_/X _5271_/X vssd1 vssd1 vccd1 vccd1 _5272_/Y sky130_fd_sc_hd__o21ai_1
X_4223_ _8377_/Q _4151_/X _4229_/S vssd1 vssd1 vccd1 vccd1 _4224_/A sky130_fd_sc_hd__mux2_1
X_4154_ _8111_/Q vssd1 vssd1 vccd1 vccd1 _4154_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4085_ _4085_/A vssd1 vssd1 vccd1 vccd1 _8416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7913_ _7913_/CLK _7913_/D vssd1 vssd1 vccd1 vccd1 _7913_/Q sky130_fd_sc_hd__dfxtp_1
X_7844_ _7844_/CLK _7844_/D vssd1 vssd1 vccd1 vccd1 _7844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7775_ _7775_/CLK _7775_/D vssd1 vssd1 vccd1 vccd1 _7775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4987_ _4987_/A vssd1 vssd1 vccd1 vccd1 _8155_/D sky130_fd_sc_hd__clkbuf_1
X_3938_ _3831_/X _8503_/Q _3946_/S vssd1 vssd1 vccd1 vccd1 _3939_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3438_ clkbuf_0__3438_/X vssd1 vssd1 vccd1 vccd1 _7021_/A sky130_fd_sc_hd__clkbuf_4
X_6657_ _6657_/A vssd1 vssd1 vccd1 vccd1 _7998_/D sky130_fd_sc_hd__clkbuf_1
X_3869_ _3869_/A _3869_/B _3869_/C _3869_/D vssd1 vssd1 vccd1 vccd1 _3870_/C sky130_fd_sc_hd__or4_1
X_5608_ _8111_/Q vssd1 vssd1 vccd1 vccd1 _5608_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8327_ _8327_/CLK _8327_/D vssd1 vssd1 vccd1 vccd1 _8327_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3406_ _6871_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3406_/X sky130_fd_sc_hd__clkbuf_16
X_5539_ _5539_/A vssd1 vssd1 vccd1 vccd1 _8029_/D sky130_fd_sc_hd__clkbuf_1
X_6888__384 _6889__385/A vssd1 vssd1 vccd1 vccd1 _8098_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7107__540 _7107__540/A vssd1 vssd1 vccd1 vccd1 _8267_/CLK sky130_fd_sc_hd__inv_2
X_8258_ _8258_/CLK _8258_/D vssd1 vssd1 vccd1 vccd1 _8258_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3654_ clkbuf_0__3654_/X vssd1 vssd1 vccd1 vccd1 _7481__15/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8189_ _8189_/CLK _8189_/D vssd1 vssd1 vccd1 vccd1 _8189_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_15_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8473_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_7209_ _7232_/C vssd1 vssd1 vccd1 vccd1 _7210_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7663__40 _7663__40/A vssd1 vssd1 vccd1 vccd1 _8509_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 caravel_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 _6129_/A sky130_fd_sc_hd__clkbuf_4
Xinput28 caravel_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_4
X_6752__348 _6753__349/A vssd1 vssd1 vccd1 vccd1 _8058_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput39 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 _5995_/A sky130_fd_sc_hd__buf_4
X_7080__518 _7082__520/A vssd1 vssd1 vccd1 vccd1 _8245_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5890_ _6654_/A _5890_/B vssd1 vssd1 vccd1 vccd1 _5891_/A sky130_fd_sc_hd__and2_1
XFILLER_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4910_ _7926_/Q _4768_/A _4791_/X _7822_/Q _4755_/A vssd1 vssd1 vccd1 vccd1 _4910_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4841_ _7976_/Q _8263_/Q _4915_/S vssd1 vssd1 vccd1 vccd1 _4841_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4772_ _4866_/S vssd1 vssd1 vccd1 vccd1 _4873_/S sky130_fd_sc_hd__clkbuf_4
X_7560_ _7567_/A _7560_/B vssd1 vssd1 vccd1 vccd1 _8464_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6511_ _6511_/A vssd1 vssd1 vccd1 vccd1 _6762_/S sky130_fd_sc_hd__clkbuf_4
X_6442_ _6521_/A vssd1 vssd1 vccd1 vccd1 _6442_/X sky130_fd_sc_hd__clkbuf_2
X_8112_ _8486_/CLK _8112_/D vssd1 vssd1 vccd1 vccd1 _8112_/Q sky130_fd_sc_hd__dfxtp_4
X_6373_ _8527_/Q _6356_/X _6372_/X _6350_/X _6358_/X vssd1 vssd1 vccd1 vccd1 _6373_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5324_ _5250_/X _5320_/X _5323_/X _5083_/X vssd1 vssd1 vccd1 vccd1 _5324_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8043_ _8043_/CLK _8043_/D vssd1 vssd1 vccd1 vccd1 _8043_/Q sky130_fd_sc_hd__dfxtp_1
X_5255_ _8381_/Q _8389_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5255_/X sky130_fd_sc_hd__mux2_1
X_4206_ _4206_/A vssd1 vssd1 vccd1 vccd1 _8384_/D sky130_fd_sc_hd__clkbuf_1
X_5186_ _5318_/S vssd1 vssd1 vccd1 vccd1 _5312_/S sky130_fd_sc_hd__buf_4
XFILLER_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _4141_/A _4622_/C _4627_/B vssd1 vssd1 vccd1 vccd1 _4137_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4068_ _4023_/X _8422_/Q _4068_/S vssd1 vssd1 vccd1 vccd1 _4069_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8593__240 vssd1 vssd1 vccd1 vccd1 _8593__240/HI partID[3] sky130_fd_sc_hd__conb_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7827_ _7827_/CLK _7827_/D vssd1 vssd1 vccd1 vccd1 _7827_/Q sky130_fd_sc_hd__dfxtp_1
X_7758_ _7633_/A _7633_/B _6082_/A _7744_/X _7729_/A vssd1 vssd1 vccd1 vccd1 _7758_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7689_ _7689_/A vssd1 vssd1 vccd1 vccd1 _7719_/A sky130_fd_sc_hd__buf_2
XFILLER_20_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3637_ clkbuf_0__3637_/X vssd1 vssd1 vccd1 vccd1 _7392__118/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5041_/A vssd1 vssd1 vccd1 vccd1 _5040_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8577__224 vssd1 vssd1 vccd1 vccd1 _8577__224/HI core1Index[4] sky130_fd_sc_hd__conb_1
X_5942_ _5942_/A vssd1 vssd1 vccd1 vccd1 _5942_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5873_ _4166_/X _7764_/Q _5875_/S vssd1 vssd1 vccd1 vccd1 _5874_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6991__449 _6992__450/A vssd1 vssd1 vccd1 vccd1 _8174_/CLK sky130_fd_sc_hd__inv_2
X_7449__164 _7450__165/A vssd1 vssd1 vccd1 vccd1 _8421_/CLK sky130_fd_sc_hd__inv_2
X_4824_ _4802_/X _4822_/X _4948_/A vssd1 vssd1 vccd1 vccd1 _4824_/X sky130_fd_sc_hd__o21a_1
X_7612_ _7602_/Y _7610_/X _7611_/X vssd1 vssd1 vccd1 vccd1 _8479_/D sky130_fd_sc_hd__o21a_1
XFILLER_21_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4755_ _4755_/A _4755_/B vssd1 vssd1 vccd1 vccd1 _4755_/X sky130_fd_sc_hd__and2_1
X_7543_ _7552_/A vssd1 vssd1 vccd1 vccd1 _7543_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4686_ _4638_/X _4662_/X _4672_/X _4685_/X vssd1 vssd1 vccd1 vccd1 _4686_/X sky130_fd_sc_hd__a31o_1
X_6425_ _8541_/Q vssd1 vssd1 vccd1 vccd1 _7529_/A sky130_fd_sc_hd__clkbuf_4
X_6356_ _6356_/A vssd1 vssd1 vccd1 vccd1 _6356_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5307_ _8309_/Q _5270_/X _5207_/X _8301_/Q _5205_/S vssd1 vssd1 vccd1 vccd1 _5307_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8026_ _8026_/CLK _8026_/D vssd1 vssd1 vccd1 vccd1 _8026_/Q sky130_fd_sc_hd__dfxtp_1
X_5238_ _5264_/A _5236_/X _5237_/X vssd1 vssd1 vccd1 vccd1 _5243_/B sky130_fd_sc_hd__o21a_1
XFILLER_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5169_ _5169_/A _5169_/B vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__and2_1
XFILLER_68_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3422_ clkbuf_0__3422_/X vssd1 vssd1 vccd1 vccd1 _6932_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6302__204 _6303__205/A vssd1 vssd1 vccd1 vccd1 _7834_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _4540_/A vssd1 vssd1 vccd1 vccd1 _8225_/D sky130_fd_sc_hd__clkbuf_1
X_4471_ _8112_/Q vssd1 vssd1 vccd1 vccd1 _4471_/X sky130_fd_sc_hd__buf_4
X_6210_ _6210_/A vssd1 vssd1 vccd1 vccd1 _6272_/A sky130_fd_sc_hd__buf_4
X_7190_ _7633_/B _6284_/X _4122_/Y _7726_/A vssd1 vssd1 vccd1 vccd1 _7385_/S sky130_fd_sc_hd__a31oi_4
X_6141_ _7805_/Q _6138_/X _6139_/X _6140_/X _6136_/X vssd1 vssd1 vccd1 vccd1 _6141_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6072_ _7862_/Q input33/X _6072_/S vssd1 vssd1 vccd1 vccd1 _6072_/X sky130_fd_sc_hd__mux2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_19 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5023_ _4432_/X _8139_/Q _5025_/S vssd1 vssd1 vccd1 vccd1 _5024_/A sky130_fd_sc_hd__mux2_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7093__528 _7093__528/A vssd1 vssd1 vccd1 vccd1 _8255_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _5925_/A vssd1 vssd1 vccd1 vccd1 _5925_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5856_ _5856_/A vssd1 vssd1 vccd1 vccd1 _7772_/D sky130_fd_sc_hd__clkbuf_1
X_4807_ _8398_/Q _4805_/Y _4806_/X _8374_/Q vssd1 vssd1 vccd1 vccd1 _4807_/X sky130_fd_sc_hd__o22a_1
X_5787_ _5787_/A _5787_/B vssd1 vssd1 vccd1 vccd1 _5803_/S sky130_fd_sc_hd__nor2_2
Xclkbuf_0__3654_ _7476_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3654_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4738_ _8148_/Q _8103_/Q _7995_/Q _8340_/Q _4868_/S _4674_/X vssd1 vssd1 vccd1 vccd1
+ _4738_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7526_ _7727_/B _6800_/B _7525_/X vssd1 vssd1 vccd1 vccd1 _7535_/B sky130_fd_sc_hd__o21a_1
XFILLER_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7457_ _7457_/A vssd1 vssd1 vccd1 vccd1 _7457_/X sky130_fd_sc_hd__buf_1
X_4669_ _4683_/B _4669_/B vssd1 vssd1 vccd1 vccd1 _4740_/A sky130_fd_sc_hd__nor2_1
XFILLER_79_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6408_ _6444_/C _8167_/Q _6382_/A _7010_/B vssd1 vssd1 vccd1 vccd1 _6408_/X sky130_fd_sc_hd__a31o_1
X_6928__402 _6931__405/A vssd1 vssd1 vccd1 vccd1 _8124_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6339_ _7877_/Q _7885_/Q _7886_/Q vssd1 vssd1 vccd1 vccd1 _6348_/C sky130_fd_sc_hd__or3_1
XFILLER_103_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8009_ _8520_/CLK _8009_/D vssd1 vssd1 vccd1 vccd1 _8009_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7430__149 _7431__150/A vssd1 vssd1 vccd1 vccd1 _8406_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7160__81 _7164__85/A vssd1 vssd1 vccd1 vccd1 _8308_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_112 _3975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_101 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3971_ _3971_/A vssd1 vssd1 vccd1 vccd1 _8455_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_123 _4517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5710_ _5710_/A vssd1 vssd1 vccd1 vccd1 _7928_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3471_ clkbuf_0__3471_/X vssd1 vssd1 vccd1 vccd1 _7156__78/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6690_ _6690_/A _6690_/B vssd1 vssd1 vccd1 vccd1 _6706_/S sky130_fd_sc_hd__and2_4
X_5641_ _5641_/A _5859_/B vssd1 vssd1 vccd1 vccd1 _5659_/S sky130_fd_sc_hd__nor2_2
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5572_ _5572_/A vssd1 vssd1 vccd1 vccd1 _5572_/X sky130_fd_sc_hd__buf_2
X_8360_ _8370_/CLK _8360_/D vssd1 vssd1 vccd1 vccd1 _8360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4523_ _8232_/Q _4478_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4524_/A sky130_fd_sc_hd__mux2_1
X_7311_ _7311_/A _7311_/B vssd1 vssd1 vccd1 vccd1 _7311_/Y sky130_fd_sc_hd__nand2_1
X_8291_ _8291_/CLK _8291_/D vssd1 vssd1 vccd1 vccd1 _8291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7242_ _8549_/Q _7311_/A _7311_/B vssd1 vssd1 vccd1 vccd1 _7242_/X sky130_fd_sc_hd__and3_1
XFILLER_116_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4454_ _4454_/A vssd1 vssd1 vccd1 vccd1 _8258_/D sky130_fd_sc_hd__clkbuf_1
X_4385_ _8492_/Q vssd1 vssd1 vccd1 vccd1 _4385_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6124_ _6465_/B vssd1 vssd1 vccd1 vccd1 _7731_/A sky130_fd_sc_hd__clkbuf_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6882__379 _6883__380/A vssd1 vssd1 vccd1 vccd1 _8093_/CLK sky130_fd_sc_hd__inv_2
X_6055_ _6034_/X _6053_/X _6054_/X _6044_/X vssd1 vssd1 vccd1 vccd1 _6055_/X sky130_fd_sc_hd__o211a_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _8146_/Q _4478_/X _5006_/S vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__mux2_1
X_7101__535 _7101__535/A vssd1 vssd1 vccd1 vccd1 _8262_/CLK sky130_fd_sc_hd__inv_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5908_ _7637_/A _5910_/B vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__or2_1
X_5839_ _7822_/Q _5575_/A _5839_/S vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3637_ _7389_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3637_/X sky130_fd_sc_hd__clkbuf_16
X_7509_ _8544_/Q _7571_/A _7571_/B vssd1 vssd1 vccd1 vccd1 _7513_/A sky130_fd_sc_hd__and3b_1
XFILLER_30_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8489_ _8530_/CLK _8489_/D vssd1 vssd1 vccd1 vccd1 _8489_/Q sky130_fd_sc_hd__dfxtp_2
X_6295__199 _6296__200/A vssd1 vssd1 vccd1 vccd1 _7829_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3319_ clkbuf_0__3319_/X vssd1 vssd1 vccd1 vccd1 _6773__360/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6716__319 _6716__319/A vssd1 vssd1 vccd1 vccd1 _8029_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4170_ _8395_/Q _4169_/X _4170_/S vssd1 vssd1 vccd1 vccd1 _4171_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7860_ _8063_/CLK _7860_/D vssd1 vssd1 vccd1 vccd1 _7860_/Q sky130_fd_sc_hd__dfxtp_1
X_6168__177 _6170__179/A vssd1 vssd1 vccd1 vccd1 _7764_/CLK sky130_fd_sc_hd__inv_2
X_6811_ _8474_/Q vssd1 vssd1 vccd1 vccd1 _6812_/B sky130_fd_sc_hd__inv_2
XFILLER_51_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7791_ _8540_/CLK _7791_/D vssd1 vssd1 vccd1 vccd1 _7791_/Q sky130_fd_sc_hd__dfxtp_1
X_3954_ _8495_/Q vssd1 vssd1 vccd1 vccd1 _3954_/X sky130_fd_sc_hd__buf_4
XFILLER_16_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3454_ clkbuf_0__3454_/X vssd1 vssd1 vccd1 vccd1 _7073__512/A sky130_fd_sc_hd__clkbuf_4
X_6673_ _6688_/S vssd1 vssd1 vccd1 vccd1 _6682_/S sky130_fd_sc_hd__clkbuf_2
X_3885_ _7885_/Q _7886_/Q _7696_/A _7877_/Q vssd1 vssd1 vccd1 vccd1 _6461_/C sky130_fd_sc_hd__or4b_4
X_5624_ _5639_/S vssd1 vssd1 vccd1 vccd1 _5633_/S sky130_fd_sc_hd__clkbuf_2
X_8412_ _8412_/CLK _8412_/D vssd1 vssd1 vccd1 vccd1 _8412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__3422_ _6925_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3422_/X sky130_fd_sc_hd__clkbuf_16
X_8343_ _8370_/CLK _8343_/D vssd1 vssd1 vccd1 vccd1 _8343_/Q sky130_fd_sc_hd__dfxtp_1
X_5555_ _5555_/A _5769_/A vssd1 vssd1 vccd1 vccd1 _5576_/S sky130_fd_sc_hd__or2_2
X_5486_ _8052_/Q _4280_/A _5492_/S vssd1 vssd1 vccd1 vccd1 _5487_/A sky130_fd_sc_hd__mux2_1
X_4506_ _4397_/X _8237_/Q _4506_/S vssd1 vssd1 vccd1 vccd1 _4507_/A sky130_fd_sc_hd__mux2_1
X_8274_ _8274_/CLK _8274_/D vssd1 vssd1 vccd1 vccd1 _8274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4437_ _4437_/A vssd1 vssd1 vccd1 vccd1 _8264_/D sky130_fd_sc_hd__clkbuf_1
X_7225_ _7510_/A _7323_/A _7323_/B vssd1 vssd1 vccd1 vccd1 _7280_/A sky130_fd_sc_hd__nand3_1
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4368_ _4292_/X _8287_/Q _4372_/S vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__mux2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _7871_/Q input11/X _6111_/S vssd1 vssd1 vccd1 vccd1 _6107_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4299_ _4298_/X _8317_/Q _4299_/S vssd1 vssd1 vccd1 vccd1 _4300_/A sky130_fd_sc_hd__mux2_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6038_ _6114_/A vssd1 vssd1 vccd1 vccd1 _6123_/B sky130_fd_sc_hd__buf_4
XFILLER_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8557__255 vssd1 vssd1 vccd1 vccd1 partID[8] _8557__255/LO sky130_fd_sc_hd__conb_1
X_7989_ _7989_/CLK _7989_/D vssd1 vssd1 vccd1 vccd1 _7989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6575__264 _6576__265/A vssd1 vssd1 vccd1 vccd1 _7942_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7443__159 _7444__160/A vssd1 vssd1 vccd1 vccd1 _8416_/CLK sky130_fd_sc_hd__inv_2
Xoutput116 _6007_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[16] sky130_fd_sc_hd__buf_2
X_5340_ _5334_/B _5334_/C _5339_/X vssd1 vssd1 vccd1 vccd1 _5340_/Y sky130_fd_sc_hd__o21ai_1
Xoutput127 _6029_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput149 _5905_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput138 _5902_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[0] sky130_fd_sc_hd__buf_2
X_5271_ _8222_/Q _5270_/X _5207_/X _8206_/Q _5055_/A vssd1 vssd1 vccd1 vccd1 _5271_/X
+ sky130_fd_sc_hd__o221a_1
X_4222_ _4222_/A vssd1 vssd1 vccd1 vccd1 _8378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7010_ _7010_/A _7010_/B vssd1 vssd1 vccd1 vccd1 _8188_/D sky130_fd_sc_hd__nor2_1
XFILLER_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4153_ _4153_/A vssd1 vssd1 vccd1 vccd1 _8401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4084_ _4015_/X _8416_/Q _4088_/S vssd1 vssd1 vccd1 vccd1 _4085_/A sky130_fd_sc_hd__mux2_1
X_7912_ _7912_/CLK _7912_/D vssd1 vssd1 vccd1 vccd1 _7912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7843_ _7843_/CLK _7843_/D vssd1 vssd1 vccd1 vccd1 _7843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7774_ _7774_/CLK _7774_/D vssd1 vssd1 vccd1 vccd1 _7774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4986_ _8155_/Q _4520_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4987_/A sky130_fd_sc_hd__mux2_1
X_6725_ _6737_/A vssd1 vssd1 vccd1 vccd1 _6725_/X sky130_fd_sc_hd__buf_1
X_3937_ _3952_/S vssd1 vssd1 vccd1 vccd1 _3946_/S sky130_fd_sc_hd__buf_2
XFILLER_51_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3437_ clkbuf_0__3437_/X vssd1 vssd1 vccd1 vccd1 _6989__447/A sky130_fd_sc_hd__clkbuf_4
X_3868_ _3868_/A _3868_/B input57/X input58/X vssd1 vssd1 vccd1 vccd1 _3870_/B sky130_fd_sc_hd__or4bb_1
X_6656_ _5919_/A _7998_/Q _6664_/S vssd1 vssd1 vccd1 vccd1 _6657_/A sky130_fd_sc_hd__mux2_1
X_5607_ _5607_/A vssd1 vssd1 vccd1 vccd1 _7980_/D sky130_fd_sc_hd__clkbuf_1
X_8326_ _8326_/CLK _8326_/D vssd1 vssd1 vccd1 vccd1 _8326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5538_ _5361_/X _8029_/Q _5546_/S vssd1 vssd1 vccd1 vccd1 _5539_/A sky130_fd_sc_hd__mux2_1
X_8257_ _8257_/CLK _8257_/D vssd1 vssd1 vccd1 vccd1 _8257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5469_ _5469_/A vssd1 vssd1 vccd1 vccd1 _8060_/D sky130_fd_sc_hd__clkbuf_1
X_7208_ _7213_/A vssd1 vssd1 vccd1 vccd1 _7210_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_0_0__3653_ clkbuf_0__3653_/X vssd1 vssd1 vccd1 vccd1 _7472__7/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8188_ _8520_/CLK _8188_/D vssd1 vssd1 vccd1 vccd1 _8188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput18 caravel_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 _6131_/A sky130_fd_sc_hd__clkbuf_4
Xinput29 caravel_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4840_ _4673_/X _4829_/X _4832_/X _4839_/X _4949_/B vssd1 vssd1 vccd1 vccd1 _4840_/X
+ sky130_fd_sc_hd__o311a_1
X_6954__420 _6954__420/A vssd1 vssd1 vccd1 vccd1 _8144_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4771_ _4880_/S vssd1 vssd1 vccd1 vccd1 _4866_/S sky130_fd_sc_hd__buf_2
X_6510_ _6510_/A vssd1 vssd1 vccd1 vccd1 _7896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6441_ _7868_/Q _6424_/X _6437_/X _6440_/X _6435_/X vssd1 vssd1 vccd1 vccd1 _7868_/D
+ sky130_fd_sc_hd__a221o_1
X_6372_ _6362_/A _7968_/Q _6352_/X _6364_/X vssd1 vssd1 vccd1 vccd1 _6372_/X sky130_fd_sc_hd__a31o_1
X_5323_ _5230_/X _5321_/X _5322_/X vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__o21a_1
X_8111_ _8486_/CLK _8111_/D vssd1 vssd1 vccd1 vccd1 _8111_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8042_ _8042_/CLK _8042_/D vssd1 vssd1 vccd1 vccd1 _8042_/Q sky130_fd_sc_hd__dfxtp_1
X_6729__329 _6730__330/A vssd1 vssd1 vccd1 vccd1 _8039_/CLK sky130_fd_sc_hd__inv_2
X_5254_ _5230_/A _5252_/X _5253_/X _5100_/A vssd1 vssd1 vccd1 vccd1 _5258_/B sky130_fd_sc_hd__o211a_1
XFILLER_87_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4205_ _8384_/Q _4181_/X _4209_/S vssd1 vssd1 vccd1 vccd1 _4206_/A sky130_fd_sc_hd__mux2_1
X_5185_ _5230_/A vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__buf_2
XFILLER_96_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4136_ _8176_/Q _8171_/Q vssd1 vssd1 vccd1 vccd1 _4622_/C sky130_fd_sc_hd__and2b_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ _4067_/A vssd1 vssd1 vccd1 vccd1 _8423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7826_ _7826_/CLK _7826_/D vssd1 vssd1 vccd1 vccd1 _7826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4969_ _8162_/Q _4478_/X _4969_/S vssd1 vssd1 vccd1 vccd1 _4970_/A sky130_fd_sc_hd__mux2_1
X_7757_ _6838_/A _7747_/Y _7756_/X vssd1 vssd1 vccd1 vccd1 _8549_/D sky130_fd_sc_hd__a21o_1
X_7688_ _7688_/A vssd1 vssd1 vccd1 vccd1 _8527_/D sky130_fd_sc_hd__clkbuf_1
X_6639_ _6755_/A vssd1 vssd1 vccd1 vccd1 _6639_/X sky130_fd_sc_hd__buf_1
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8309_ _8309_/CLK _8309_/D vssd1 vssd1 vccd1 vccd1 _8309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3319_ _6768_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3319_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_94_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6526__225 _6526__225/A vssd1 vssd1 vccd1 vccd1 _7903_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7167__87 _7169__89/A vssd1 vssd1 vccd1 vccd1 _8314_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5941_ _5941_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5942_/A sky130_fd_sc_hd__or2_1
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5872_ _5872_/A vssd1 vssd1 vccd1 vccd1 _7765_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_0_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _8370_/CLK sky130_fd_sc_hd__clkbuf_16
X_7611_ _8479_/Q _7597_/X _7552_/A vssd1 vssd1 vccd1 vccd1 _7611_/X sky130_fd_sc_hd__o21a_1
X_4823_ _4823_/A vssd1 vssd1 vccd1 vccd1 _4948_/A sky130_fd_sc_hd__buf_2
X_4754_ _7826_/Q _7946_/Q _7962_/Q _7930_/Q _4729_/X _4716_/A vssd1 vssd1 vccd1 vccd1
+ _4755_/B sky130_fd_sc_hd__mux4_2
X_7542_ _7588_/A vssd1 vssd1 vccd1 vccd1 _7542_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4685_ _4673_/X _4677_/X _4682_/X _4684_/X vssd1 vssd1 vccd1 vccd1 _4685_/X sky130_fd_sc_hd__o211a_2
X_6424_ _6521_/A vssd1 vssd1 vccd1 vccd1 _6424_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6355_ _6355_/A _6355_/B vssd1 vssd1 vccd1 vccd1 _6356_/A sky130_fd_sc_hd__nor2_1
X_5306_ _5306_/A _5306_/B vssd1 vssd1 vccd1 vccd1 _5306_/X sky130_fd_sc_hd__or2_1
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6286_ _7359_/A _6282_/X _7308_/A _7360_/B vssd1 vssd1 vccd1 vccd1 _7821_/D sky130_fd_sc_hd__a211o_4
XFILLER_102_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5237_ _8311_/Q _5270_/A _5319_/B _8303_/Q _5125_/A vssd1 vssd1 vccd1 vccd1 _5237_/X
+ sky130_fd_sc_hd__o221a_1
X_8025_ _8025_/CLK _8025_/D vssd1 vssd1 vccd1 vccd1 _8025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5168_ _8508_/Q _8257_/Q _8241_/Q _8281_/Q _5087_/X _5061_/A vssd1 vssd1 vccd1 vccd1
+ _5169_/B sky130_fd_sc_hd__mux4_2
XFILLER_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3421_ clkbuf_0__3421_/X vssd1 vssd1 vccd1 vccd1 _6924__400/A sky130_fd_sc_hd__clkbuf_4
X_6629__293 _6631__295/A vssd1 vssd1 vccd1 vccd1 _7979_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5099_ _8426_/Q _8324_/Q _8061_/Q _8276_/Q _5080_/A _5308_/S vssd1 vssd1 vccd1 vccd1
+ _5099_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4119_ _8174_/Q vssd1 vssd1 vccd1 vccd1 _4217_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7809_ _8487_/CLK _7809_/D vssd1 vssd1 vccd1 vccd1 _7809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7051__495 _7051__495/A vssd1 vssd1 vccd1 vccd1 _8222_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4470_ _4470_/A vssd1 vssd1 vccd1 vccd1 _8252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6140_ _6140_/A _6140_/B vssd1 vssd1 vccd1 vccd1 _6140_/X sky130_fd_sc_hd__and2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6071_ _6056_/X _6068_/X _6070_/X _6063_/X vssd1 vssd1 vccd1 vccd1 _6071_/X sky130_fd_sc_hd__o211a_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5022_/A vssd1 vssd1 vccd1 vccd1 _8140_/D sky130_fd_sc_hd__clkbuf_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5924_ _5924_/A _5932_/B vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__or2_4
XFILLER_110_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5855_ _4166_/X _7772_/Q _5857_/S vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3653_ _7470_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3653_/X sky130_fd_sc_hd__clkbuf_16
X_4806_ _4806_/A vssd1 vssd1 vccd1 vccd1 _4806_/X sky130_fd_sc_hd__buf_2
XFILLER_21_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5786_ _5786_/A vssd1 vssd1 vccd1 vccd1 _7846_/D sky130_fd_sc_hd__clkbuf_1
X_4737_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4868_/S sky130_fd_sc_hd__clkbuf_4
X_7525_ _8540_/Q _7525_/B vssd1 vssd1 vccd1 vccd1 _7525_/X sky130_fd_sc_hd__xor2_1
X_4668_ _8378_/Q _8268_/Q _7981_/Q _8402_/Q _4666_/X _4667_/X vssd1 vssd1 vccd1 vccd1
+ _4668_/X sky130_fd_sc_hd__mux4_2
X_6407_ _8063_/Q vssd1 vssd1 vccd1 vccd1 _6444_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4599_ _4599_/A vssd1 vssd1 vccd1 vccd1 _8199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6338_ _6517_/A _6417_/A vssd1 vssd1 vccd1 vccd1 _6341_/A sky130_fd_sc_hd__or2b_1
XFILLER_88_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6269_ _7820_/Q _7819_/Q _6269_/C vssd1 vssd1 vccd1 vccd1 _6272_/C sky130_fd_sc_hd__or3_1
X_8008_ _8520_/CLK _8008_/D vssd1 vssd1 vccd1 vccd1 _8008_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7398__123 _7399__124/A vssd1 vssd1 vccd1 vccd1 _8380_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_102 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_124 _4517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _8455_/Q _3969_/X _3973_/S vssd1 vssd1 vccd1 vccd1 _3971_/A sky130_fd_sc_hd__mux2_1
XINSDIODE2_113 _3981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3470_ clkbuf_0__3470_/X vssd1 vssd1 vccd1 vccd1 _7177_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5640_ _5640_/A vssd1 vssd1 vccd1 vccd1 _7958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6539__235 _6539__235/A vssd1 vssd1 vccd1 vccd1 _7913_/CLK sky130_fd_sc_hd__inv_2
X_5571_ _5571_/A vssd1 vssd1 vccd1 vccd1 _7992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4522_ _4522_/A vssd1 vssd1 vccd1 vccd1 _8233_/D sky130_fd_sc_hd__clkbuf_1
X_7310_ _7310_/A vssd1 vssd1 vccd1 vccd1 _7310_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_8290_ _8290_/CLK _8290_/D vssd1 vssd1 vccd1 vccd1 _8290_/Q sky130_fd_sc_hd__dfxtp_1
X_4453_ _4382_/X _8258_/Q _4457_/S vssd1 vssd1 vccd1 vccd1 _4454_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7241_ _8344_/Q _8343_/Q _8345_/Q vssd1 vssd1 vccd1 vccd1 _7311_/B sky130_fd_sc_hd__a21o_1
X_4384_ _4384_/A vssd1 vssd1 vccd1 vccd1 _8282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6123_/A _6123_/B vssd1 vssd1 vccd1 vccd1 _6123_/X sky130_fd_sc_hd__and2_1
XFILLER_105_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6054_ _7782_/Q _6066_/B vssd1 vssd1 vccd1 vccd1 _6054_/X sky130_fd_sc_hd__or2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5005_ _5005_/A vssd1 vssd1 vccd1 vccd1 _8147_/D sky130_fd_sc_hd__clkbuf_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6923__399 _6923__399/A vssd1 vssd1 vccd1 vccd1 _8121_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5907_ _5907_/A vssd1 vssd1 vccd1 vccd1 _5907_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7466__2 _7466__2/A vssd1 vssd1 vccd1 vccd1 _8434_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5838_ _5838_/A vssd1 vssd1 vccd1 vccd1 _7823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5769_ _5769_/A _5859_/B vssd1 vssd1 vccd1 vccd1 _5785_/S sky130_fd_sc_hd__or2_2
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7508_ _8542_/Q _7514_/B _7506_/X _7507_/Y vssd1 vssd1 vccd1 vccd1 _7524_/A sky130_fd_sc_hd__a211o_1
XFILLER_107_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8488_ _8527_/CLK _8488_/D vssd1 vssd1 vccd1 vccd1 _8488_/Q sky130_fd_sc_hd__dfxtp_2
X_7439_ _7439_/A vssd1 vssd1 vccd1 vccd1 _7439_/X sky130_fd_sc_hd__buf_1
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3249_ clkbuf_0__3249_/X vssd1 vssd1 vccd1 vccd1 _6554__247/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6315__215 _6315__215/A vssd1 vssd1 vccd1 vccd1 _7845_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7133__60 _7133__60/A vssd1 vssd1 vccd1 vccd1 _8287_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6810_ _8475_/Q vssd1 vssd1 vccd1 vccd1 _6812_/A sky130_fd_sc_hd__inv_2
X_7790_ _8540_/CLK _7790_/D vssd1 vssd1 vccd1 vccd1 _7790_/Q sky130_fd_sc_hd__dfxtp_1
X_3953_ _3953_/A vssd1 vssd1 vccd1 vccd1 _8496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3453_ clkbuf_0__3453_/X vssd1 vssd1 vccd1 vccd1 _7069__509/A sky130_fd_sc_hd__clkbuf_4
X_6672_ _6672_/A _6690_/B vssd1 vssd1 vccd1 vccd1 _6688_/S sky130_fd_sc_hd__nand2_2
X_3884_ _7878_/Q _6348_/B vssd1 vssd1 vccd1 vccd1 _6461_/B sky130_fd_sc_hd__or2_2
X_8411_ _8411_/CLK _8411_/D vssd1 vssd1 vccd1 vccd1 _8411_/Q sky130_fd_sc_hd__dfxtp_1
X_5623_ _5769_/A _5823_/B vssd1 vssd1 vccd1 vccd1 _5639_/S sky130_fd_sc_hd__or2_2
X_8342_ _8342_/CLK _8342_/D vssd1 vssd1 vccd1 vccd1 _8342_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3421_ _6919_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3421_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5554_ _5554_/A vssd1 vssd1 vccd1 vccd1 _5554_/X sky130_fd_sc_hd__buf_2
X_5485_ _5485_/A vssd1 vssd1 vccd1 vccd1 _8053_/D sky130_fd_sc_hd__clkbuf_1
X_8273_ _8273_/CLK _8273_/D vssd1 vssd1 vccd1 vccd1 _8273_/Q sky130_fd_sc_hd__dfxtp_1
X_4505_ _4505_/A vssd1 vssd1 vccd1 vccd1 _8238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4436_ _4435_/X _8264_/Q _4436_/S vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__mux2_1
X_7224_ _8348_/Q _8347_/Q _7236_/B _8349_/Q vssd1 vssd1 vccd1 vccd1 _7323_/B sky130_fd_sc_hd__a31o_1
XFILLER_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7675__50 _7675__50/A vssd1 vssd1 vccd1 vccd1 _8519_/CLK sky130_fd_sc_hd__inv_2
X_4367_ _4367_/A vssd1 vssd1 vccd1 vccd1 _8288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6106_ _6095_/X _6104_/X _6105_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6106_/X sky130_fd_sc_hd__o211a_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4298_/A vssd1 vssd1 vccd1 vccd1 _4298_/X sky130_fd_sc_hd__clkbuf_2
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6037_ _6466_/B vssd1 vssd1 vccd1 vccd1 _6114_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7988_ _7988_/CLK _7988_/D vssd1 vssd1 vccd1 vccd1 _7988_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6939_ _7646_/C vssd1 vssd1 vccd1 vccd1 _7640_/C sky130_fd_sc_hd__clkbuf_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6722__324 _6723__325/A vssd1 vssd1 vccd1 vccd1 _8034_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7649__28 _7651__30/A vssd1 vssd1 vccd1 vccd1 _8497_/CLK sky130_fd_sc_hd__inv_2
Xoutput128 _6031_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[27] sky130_fd_sc_hd__buf_2
Xoutput117 _6009_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[17] sky130_fd_sc_hd__buf_2
Xoutput139 _5925_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[10] sky130_fd_sc_hd__buf_2
X_5270_ _5270_/A vssd1 vssd1 vccd1 vccd1 _5270_/X sky130_fd_sc_hd__buf_2
X_4221_ _8378_/Q _4114_/X _4229_/S vssd1 vssd1 vccd1 vccd1 _4222_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6174__182 _6175__183/A vssd1 vssd1 vccd1 vccd1 _7769_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4152_ _8401_/Q _4151_/X _4161_/S vssd1 vssd1 vccd1 vccd1 _4153_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4083_ _4083_/A vssd1 vssd1 vccd1 vccd1 _8417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7911_ _7911_/CLK _7911_/D vssd1 vssd1 vccd1 vccd1 _7911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7842_ _7842_/CLK _7842_/D vssd1 vssd1 vccd1 vccd1 _7842_/Q sky130_fd_sc_hd__dfxtp_1
X_6623__288 _6625__290/A vssd1 vssd1 vccd1 vccd1 _7974_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7773_ _7773_/CLK _7773_/D vssd1 vssd1 vccd1 vccd1 _7773_/Q sky130_fd_sc_hd__dfxtp_1
X_4985_ _4985_/A vssd1 vssd1 vccd1 vccd1 _8156_/D sky130_fd_sc_hd__clkbuf_1
X_6724_ _6755_/A vssd1 vssd1 vccd1 vccd1 _6724_/X sky130_fd_sc_hd__buf_1
X_3936_ _5500_/A _5428_/A vssd1 vssd1 vccd1 vccd1 _3952_/S sky130_fd_sc_hd__or2_2
XFILLER_51_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3436_ clkbuf_0__3436_/X vssd1 vssd1 vccd1 vccd1 _6986__445/A sky130_fd_sc_hd__clkbuf_4
X_6655_ _6670_/S vssd1 vssd1 vccd1 vccd1 _6664_/S sky130_fd_sc_hd__clkbuf_2
X_3867_ _3867_/A _3867_/B input69/X vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__or3b_1
XFILLER_31_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5606_ _5559_/X _7980_/Q _5614_/S vssd1 vssd1 vccd1 vccd1 _5607_/A sky130_fd_sc_hd__mux2_1
X_8325_ _8325_/CLK _8325_/D vssd1 vssd1 vccd1 vccd1 _8325_/Q sky130_fd_sc_hd__dfxtp_1
X_5537_ _5552_/S vssd1 vssd1 vccd1 vccd1 _5546_/S sky130_fd_sc_hd__buf_2
XFILLER_117_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8256_ _8256_/CLK _8256_/D vssd1 vssd1 vccd1 vccd1 _8256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5468_ _3963_/X _8060_/Q _5474_/S vssd1 vssd1 vccd1 vccd1 _5469_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7207_ _7207_/A _7277_/C _7207_/C vssd1 vssd1 vccd1 vccd1 _7263_/B sky130_fd_sc_hd__and3_1
Xclkbuf_1_0_0__3652_ clkbuf_0__3652_/X vssd1 vssd1 vccd1 vccd1 _7469__5/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5399_ _5399_/A vssd1 vssd1 vccd1 vccd1 _5399_/X sky130_fd_sc_hd__clkbuf_4
X_8187_ _8520_/CLK _8187_/D vssd1 vssd1 vccd1 vccd1 _8187_/Q sky130_fd_sc_hd__dfxtp_1
X_4419_ _4929_/A _4944_/A _4931_/B vssd1 vssd1 vccd1 vccd1 _5841_/A sky130_fd_sc_hd__or3_4
XFILLER_101_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 caravel_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 _6133_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4770_ _4809_/A vssd1 vssd1 vccd1 vccd1 _4770_/X sky130_fd_sc_hd__buf_2
XFILLER_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6440_ _6440_/A _6452_/B _6444_/C vssd1 vssd1 vccd1 vccd1 _6440_/X sky130_fd_sc_hd__and3_1
X_6371_ _6838_/A _6362_/X _6336_/X _6343_/X vssd1 vssd1 vccd1 vccd1 _6371_/X sky130_fd_sc_hd__a31o_1
XFILLER_114_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5322_ _8411_/Q _5270_/A _5319_/B _8403_/Q _5125_/A vssd1 vssd1 vccd1 vccd1 _5322_/X
+ sky130_fd_sc_hd__o221a_1
X_8110_ _8480_/CLK _8110_/D vssd1 vssd1 vccd1 vccd1 _8110_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8041_ _8041_/CLK _8041_/D vssd1 vssd1 vccd1 vccd1 _8041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5253_ _8445_/Q _5232_/A _5214_/A _8437_/Q vssd1 vssd1 vccd1 vccd1 _5253_/X sky130_fd_sc_hd__o22a_1
X_4204_ _4204_/A vssd1 vssd1 vccd1 vccd1 _8385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5184_ _5192_/A vssd1 vssd1 vccd1 vccd1 _5230_/A sky130_fd_sc_hd__clkbuf_2
X_7419__140 _7419__140/A vssd1 vssd1 vccd1 vccd1 _8397_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4135_ _4627_/B _4141_/A vssd1 vssd1 vccd1 vccd1 _4135_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ _4019_/X _8423_/Q _4068_/S vssd1 vssd1 vccd1 vccd1 _4067_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7825_ _7825_/CLK _7825_/D vssd1 vssd1 vccd1 vccd1 _7825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4968_ _4968_/A vssd1 vssd1 vccd1 vccd1 _8163_/D sky130_fd_sc_hd__clkbuf_1
X_7756_ _7635_/A _7702_/X _7743_/X _7729_/A vssd1 vssd1 vccd1 vccd1 _7756_/X sky130_fd_sc_hd__a31o_1
X_4899_ _8395_/Q _4805_/Y _4777_/X _8371_/Q _4677_/S vssd1 vssd1 vccd1 vccd1 _4899_/X
+ sky130_fd_sc_hd__o221a_1
X_6707_ _6707_/A vssd1 vssd1 vccd1 vccd1 _8021_/D sky130_fd_sc_hd__clkbuf_1
X_7687_ _7687_/A _8521_/Q vssd1 vssd1 vccd1 vccd1 _7688_/A sky130_fd_sc_hd__and2_1
X_3919_ _3831_/X _8511_/Q _3927_/S vssd1 vssd1 vccd1 vccd1 _3920_/A sky130_fd_sc_hd__mux2_1
X_6638_ _6961_/A vssd1 vssd1 vccd1 vccd1 _6638_/X sky130_fd_sc_hd__buf_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8308_ _8308_/CLK _8308_/D vssd1 vssd1 vccd1 vccd1 _8308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8239_ _8239_/CLK _8239_/D vssd1 vssd1 vccd1 vccd1 _8239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3249_ _6552_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3249_/X sky130_fd_sc_hd__clkbuf_16
X_7392__118 _7392__118/A vssd1 vssd1 vccd1 vccd1 _8375_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8602__249 vssd1 vssd1 vccd1 vccd1 _8602__249/HI versionID[3] sky130_fd_sc_hd__conb_1
XFILLER_101_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5940_ _5940_/A vssd1 vssd1 vccd1 vccd1 _5940_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5871_ _4163_/X _7765_/Q _5875_/S vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__mux2_1
X_7610_ _8479_/Q _7606_/B _7609_/Y vssd1 vssd1 vccd1 vccd1 _7610_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4822_ _4740_/X _4808_/X _4813_/X _4821_/X _4638_/X vssd1 vssd1 vccd1 vccd1 _4822_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_119_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6735__334 _6736__335/A vssd1 vssd1 vccd1 vccd1 _8044_/CLK sky130_fd_sc_hd__inv_2
X_4753_ _4953_/B _4750_/X _4752_/X vssd1 vssd1 vccd1 vccd1 _4753_/X sky130_fd_sc_hd__a21o_1
X_7541_ _7541_/A vssd1 vssd1 vccd1 vccd1 _7588_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4684_ _4801_/A vssd1 vssd1 vccd1 vccd1 _4684_/X sky130_fd_sc_hd__clkbuf_2
X_6423_ _7863_/Q _6388_/X _6415_/X _6420_/X _6422_/X vssd1 vssd1 vccd1 vccd1 _7863_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7063__504 _7063__504/A vssd1 vssd1 vccd1 vccd1 _8231_/CLK sky130_fd_sc_hd__inv_2
X_6354_ _7741_/A _7966_/Q _6352_/X _6395_/A vssd1 vssd1 vccd1 vccd1 _6354_/X sky130_fd_sc_hd__a31o_1
XFILLER_88_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5305_ _8285_/Q _8293_/Q _5305_/S vssd1 vssd1 vccd1 vccd1 _5306_/B sky130_fd_sc_hd__mux2_1
X_6285_ _5903_/A _6284_/X _4122_/Y _6466_/A vssd1 vssd1 vccd1 vccd1 _7360_/B sky130_fd_sc_hd__a31o_4
XFILLER_102_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6588__275 _6588__275/A vssd1 vssd1 vccd1 vccd1 _7953_/CLK sky130_fd_sc_hd__inv_2
X_5236_ _8287_/Q _8295_/Q _5312_/S vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__mux2_1
X_8024_ _8024_/CLK _8024_/D vssd1 vssd1 vccd1 vccd1 _8024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5167_ _5165_/X _5166_/X _5167_/S vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5098_ _5318_/S vssd1 vssd1 vccd1 vccd1 _5308_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4118_ _4466_/B _4933_/C _5622_/A vssd1 vssd1 vccd1 vccd1 _5602_/A sky130_fd_sc_hd__or3b_4
XFILLER_17_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4049_ _4023_/X _8430_/Q _4049_/S vssd1 vssd1 vccd1 vccd1 _4050_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7808_ _8487_/CLK _7808_/D vssd1 vssd1 vccd1 vccd1 _7808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7739_ _5919_/A _7731_/X _7723_/X vssd1 vssd1 vccd1 vccd1 _7739_/X sky130_fd_sc_hd__a21bo_1
XFILLER_4_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7172__91 _7173__92/A vssd1 vssd1 vccd1 vccd1 _8318_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7400__125 _7400__125/A vssd1 vssd1 vccd1 vccd1 _8382_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8583__230 vssd1 vssd1 vccd1 vccd1 _8583__230/HI manufacturerID[2] sky130_fd_sc_hd__conb_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _7786_/Q _6086_/B vssd1 vssd1 vccd1 vccd1 _6070_/X sky130_fd_sc_hd__or2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5021_ _4428_/X _8140_/Q _5025_/S vssd1 vssd1 vccd1 vccd1 _5022_/A sky130_fd_sc_hd__mux2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5923_ _5956_/A vssd1 vssd1 vccd1 vccd1 _5932_/B sky130_fd_sc_hd__clkbuf_2
X_5854_ _5854_/A vssd1 vssd1 vccd1 vccd1 _7773_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3652_ _7464_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3652_/X sky130_fd_sc_hd__clkbuf_16
X_4805_ _4805_/A vssd1 vssd1 vccd1 vccd1 _4805_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5785_ _5575_/X _7846_/Q _5785_/S vssd1 vssd1 vccd1 vccd1 _5786_/A sky130_fd_sc_hd__mux2_1
X_7524_ _7524_/A _7524_/B _7524_/C _7524_/D vssd1 vssd1 vccd1 vccd1 _7524_/X sky130_fd_sc_hd__or4_1
X_4736_ _8250_/Q _8035_/Q _7987_/Q _7939_/Q _4729_/X _4716_/A vssd1 vssd1 vccd1 vccd1
+ _4736_/X sky130_fd_sc_hd__mux4_2
XFILLER_107_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4667_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4667_/X sky130_fd_sc_hd__buf_2
X_6406_ _6331_/X _6404_/X _6405_/X vssd1 vssd1 vccd1 vccd1 _7861_/D sky130_fd_sc_hd__a21o_1
X_7386_ _7386_/A vssd1 vssd1 vccd1 vccd1 _8370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4598_ _4438_/X _8199_/Q _4602_/S vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6337_ _6337_/A vssd1 vssd1 vccd1 vccd1 _7742_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6268_ _7820_/Q _7819_/Q vssd1 vssd1 vccd1 vccd1 _6270_/B sky130_fd_sc_hd__nand2_1
X_5219_ _5227_/A _8076_/Q _7841_/Q _5214_/A _5125_/A vssd1 vssd1 vccd1 vccd1 _5219_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6199_ _6367_/A vssd1 vssd1 vccd1 vccd1 _6235_/A sky130_fd_sc_hd__clkbuf_2
X_8007_ _8520_/CLK _8007_/D vssd1 vssd1 vccd1 vccd1 _8007_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6974__435 _6974__435/A vssd1 vssd1 vccd1 vccd1 _8159_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6935__408 _6936__409/A vssd1 vssd1 vccd1 vccd1 _8130_/CLK sky130_fd_sc_hd__inv_2
X_6603__286 _6604__287/A vssd1 vssd1 vccd1 vccd1 _7964_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8567__214 vssd1 vssd1 vccd1 vccd1 _8567__214/HI core0Index[1] sky130_fd_sc_hd__conb_1
XFILLER_4_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_103 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_114 _4517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5570_ _5569_/X _7992_/Q _5576_/S vssd1 vssd1 vccd1 vccd1 _5571_/A sky130_fd_sc_hd__mux2_1
X_4521_ _8233_/Q _4520_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4522_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4452_ _4452_/A vssd1 vssd1 vccd1 vccd1 _8259_/D sky130_fd_sc_hd__clkbuf_1
X_7240_ _7754_/A _7240_/B vssd1 vssd1 vccd1 vccd1 _7280_/C sky130_fd_sc_hd__xor2_1
XFILLER_116_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7171_ _7177_/A vssd1 vssd1 vccd1 vccd1 _7171_/X sky130_fd_sc_hd__buf_1
X_4383_ _4382_/X _8282_/Q _4389_/S vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6122_/A vssd1 vssd1 vccd1 vccd1 _6122_/X sky130_fd_sc_hd__clkbuf_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _7857_/Q input28/X _6123_/B vssd1 vssd1 vccd1 vccd1 _6053_/X sky130_fd_sc_hd__mux2_1
X_5004_ _8147_/Q _4520_/X _5006_/S vssd1 vssd1 vccd1 vccd1 _5005_/A sky130_fd_sc_hd__mux2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _6955_/A vssd1 vssd1 vccd1 vccd1 _6955_/X sky130_fd_sc_hd__buf_1
X_5906_ _7635_/A _5910_/B vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__or2_1
XFILLER_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5837_ _7823_/Q _5572_/A _5839_/S vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5768_ _5768_/A vssd1 vssd1 vccd1 vccd1 _7902_/D sky130_fd_sc_hd__clkbuf_1
X_4719_ _8218_/Q _8202_/Q _8164_/Q _8234_/Q _4915_/S _4649_/X vssd1 vssd1 vccd1 vccd1
+ _4719_/X sky130_fd_sc_hd__mux4_1
X_7507_ _7576_/A _7576_/B _6854_/A vssd1 vssd1 vccd1 vccd1 _7507_/Y sky130_fd_sc_hd__a21boi_1
X_8487_ _8487_/CLK _8487_/D vssd1 vssd1 vccd1 vccd1 _8487_/Q sky130_fd_sc_hd__dfxtp_1
X_5699_ _7933_/Q _5578_/X _5707_/S vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7369_ _8125_/Q _7679_/B _7366_/X _7368_/X _7286_/X vssd1 vssd1 vccd1 vccd1 _8362_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7002__457 _7002__457/A vssd1 vssd1 vccd1 vccd1 _8182_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3248_ clkbuf_0__3248_/X vssd1 vssd1 vccd1 vccd1 _6551__245/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6545__240 _6545__240/A vssd1 vssd1 vccd1 vccd1 _7918_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7413__135 _7413__135/A vssd1 vssd1 vccd1 vccd1 _8392_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3952_ _3911_/X _8496_/Q _3952_/S vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3452_ clkbuf_0__3452_/X vssd1 vssd1 vccd1 vccd1 _7063__504/A sky130_fd_sc_hd__clkbuf_4
X_6671_ _6671_/A vssd1 vssd1 vccd1 vccd1 _8005_/D sky130_fd_sc_hd__clkbuf_1
X_3883_ _7696_/A _7696_/B _7696_/C _7696_/D vssd1 vssd1 vccd1 vccd1 _6348_/B sky130_fd_sc_hd__or4_1
X_8410_ _8410_/CLK _8410_/D vssd1 vssd1 vccd1 vccd1 _8410_/Q sky130_fd_sc_hd__dfxtp_1
X_5622_ _5622_/A _8175_/Q _4466_/B vssd1 vssd1 vccd1 vccd1 _5823_/B sky130_fd_sc_hd__or3b_4
X_8341_ _8341_/CLK _8341_/D vssd1 vssd1 vccd1 vccd1 _8341_/Q sky130_fd_sc_hd__dfxtp_1
X_5553_ _5553_/A vssd1 vssd1 vccd1 vccd1 _8022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4504_ _4394_/X _8238_/Q _4506_/S vssd1 vssd1 vccd1 vccd1 _4505_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5484_ _8053_/Q _4275_/A _5492_/S vssd1 vssd1 vccd1 vccd1 _5485_/A sky130_fd_sc_hd__mux2_1
X_8272_ _8272_/CLK _8272_/D vssd1 vssd1 vccd1 vccd1 _8272_/Q sky130_fd_sc_hd__dfxtp_1
X_7223_ _8349_/Q _7227_/A _7236_/A _7232_/B vssd1 vssd1 vccd1 vccd1 _7323_/A sky130_fd_sc_hd__nand4_2
X_4435_ _8109_/Q vssd1 vssd1 vccd1 vccd1 _4435_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4366_ _4289_/X _8288_/Q _4366_/S vssd1 vssd1 vccd1 vccd1 _4367_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _7795_/Q _6105_/B vssd1 vssd1 vccd1 vccd1 _6105_/X sky130_fd_sc_hd__or2_1
X_4297_ _4297_/A vssd1 vssd1 vccd1 vccd1 _8318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6465_/B _5878_/B _5879_/X _7762_/Q vssd1 vssd1 vccd1 vccd1 _6466_/B sky130_fd_sc_hd__a31oi_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7987_ _7987_/CLK _7987_/D vssd1 vssd1 vccd1 vccd1 _7987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ _6941_/B _6938_/B vssd1 vssd1 vccd1 vccd1 _7646_/C sky130_fd_sc_hd__and2_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8539_ _8540_/CLK _8539_/D vssd1 vssd1 vccd1 vccd1 _8539_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6321__220 _6321__220/A vssd1 vssd1 vccd1 vccd1 _7850_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput118 _6012_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput129 _5976_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[2] sky130_fd_sc_hd__buf_2
X_4220_ _4235_/S vssd1 vssd1 vccd1 vccd1 _4229_/S sky130_fd_sc_hd__buf_2
X_4151_ _8112_/Q vssd1 vssd1 vccd1 vccd1 _4151_/X sky130_fd_sc_hd__clkbuf_4
X_4082_ _4011_/X _8417_/Q _4088_/S vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7910_ _7910_/CLK _7910_/D vssd1 vssd1 vccd1 vccd1 _7910_/Q sky130_fd_sc_hd__dfxtp_1
X_7841_ _7841_/CLK _7841_/D vssd1 vssd1 vccd1 vccd1 _7841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7772_ _7772_/CLK _7772_/D vssd1 vssd1 vccd1 vccd1 _7772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4984_ _8156_/Q _4517_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4985_/A sky130_fd_sc_hd__mux2_1
X_3935_ _3956_/B _4038_/A _5345_/B _5109_/A vssd1 vssd1 vccd1 vccd1 _5428_/A sky130_fd_sc_hd__or4b_4
Xclkbuf_1_1_0__3435_ clkbuf_0__3435_/X vssd1 vssd1 vccd1 vccd1 _6979__439/A sky130_fd_sc_hd__clkbuf_4
X_6654_ _6654_/A _6690_/B vssd1 vssd1 vccd1 vccd1 _6670_/S sky130_fd_sc_hd__nand2_2
X_5605_ _5605_/A vssd1 vssd1 vccd1 vccd1 _7981_/D sky130_fd_sc_hd__clkbuf_1
X_3866_ _3866_/A _3866_/B _3866_/C _3866_/D vssd1 vssd1 vccd1 vccd1 _3871_/C sky130_fd_sc_hd__or4_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8324_ _8324_/CLK _8324_/D vssd1 vssd1 vccd1 vccd1 _8324_/Q sky130_fd_sc_hd__dfxtp_1
X_5536_ _5661_/A _5751_/B vssd1 vssd1 vccd1 vccd1 _5552_/S sky130_fd_sc_hd__or2_2
XFILLER_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5467_ _5467_/A vssd1 vssd1 vccd1 vccd1 _8061_/D sky130_fd_sc_hd__clkbuf_1
X_8255_ _8255_/CLK _8255_/D vssd1 vssd1 vccd1 vccd1 _8255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7206_ _8537_/Q _7344_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _7207_/C sky130_fd_sc_hd__nand3b_1
X_4418_ _8113_/Q vssd1 vssd1 vccd1 vccd1 _4418_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0_0__3651_ clkbuf_0__3651_/X vssd1 vssd1 vccd1 vccd1 _7482_/A sky130_fd_sc_hd__clkbuf_4
X_8186_ _8186_/CLK _8186_/D vssd1 vssd1 vccd1 vccd1 _8186_/Q sky130_fd_sc_hd__dfxtp_1
X_5398_ _5398_/A vssd1 vssd1 vccd1 vccd1 _8095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4349_ _4349_/A vssd1 vssd1 vccd1 vccd1 _8296_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6019_ _8012_/Q _6019_/B vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__and2_1
X_6641__301 _6643__303/A vssd1 vssd1 vccd1 vccd1 _7987_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7179__97 _7179__97/A vssd1 vssd1 vccd1 vccd1 _8324_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7654__32 _7656__34/A vssd1 vssd1 vccd1 vccd1 _8501_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7187__103 _7189__105/A vssd1 vssd1 vccd1 vccd1 _8330_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6370_ _8549_/Q vssd1 vssd1 vccd1 vccd1 _6838_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5321_ _8379_/Q _8387_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8040_ _8040_/CLK _8040_/D vssd1 vssd1 vccd1 vccd1 _8040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5252_ _7832_/Q _8429_/Q _5252_/S vssd1 vssd1 vccd1 vccd1 _5252_/X sky130_fd_sc_hd__mux2_1
X_4203_ _8385_/Q _4178_/X _4209_/S vssd1 vssd1 vccd1 vccd1 _4204_/A sky130_fd_sc_hd__mux2_1
X_5183_ _5183_/A _5197_/A vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__nand2_1
XFILLER_110_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4134_ _8175_/Q _4217_/A _8173_/Q vssd1 vssd1 vccd1 vccd1 _4141_/A sky130_fd_sc_hd__nand3_2
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4065_ _4065_/A vssd1 vssd1 vccd1 vccd1 _8424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7824_ _7824_/CLK _7824_/D vssd1 vssd1 vccd1 vccd1 _7824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4967_ _8163_/Q _4520_/X _4969_/S vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7755_ _3873_/X _7747_/Y _7754_/X _7687_/A vssd1 vssd1 vccd1 vccd1 _8548_/D sky130_fd_sc_hd__o211a_1
X_4898_ _7974_/Q _8261_/Q _4901_/S vssd1 vssd1 vccd1 vccd1 _4898_/X sky130_fd_sc_hd__mux2_1
X_3918_ _3933_/S vssd1 vssd1 vccd1 vccd1 _3927_/S sky130_fd_sc_hd__clkbuf_2
X_6706_ _8021_/Q _5969_/A _6706_/S vssd1 vssd1 vccd1 vccd1 _6707_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7686_ _7686_/A vssd1 vssd1 vccd1 vccd1 _8526_/D sky130_fd_sc_hd__clkbuf_1
X_3849_ _5035_/A _3849_/B vssd1 vssd1 vccd1 vccd1 _3860_/B sky130_fd_sc_hd__and2b_1
XFILLER_118_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7479__13 _7479__13/A vssd1 vssd1 vccd1 vccd1 _8445_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5519_ _5534_/S vssd1 vssd1 vccd1 vccd1 _5528_/S sky130_fd_sc_hd__buf_2
X_8307_ _8307_/CLK _8307_/D vssd1 vssd1 vccd1 vccd1 _8307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6499_ _6499_/A vssd1 vssd1 vccd1 vccd1 _7891_/D sky130_fd_sc_hd__clkbuf_1
X_8238_ _8238_/CLK _8238_/D vssd1 vssd1 vccd1 vccd1 _8238_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3248_ _6546_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3248_/X sky130_fd_sc_hd__clkbuf_16
X_8169_ _8169_/CLK _8169_/D vssd1 vssd1 vccd1 vccd1 _8169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6648__307 _6651__310/A vssd1 vssd1 vccd1 vccd1 _7993_/CLK sky130_fd_sc_hd__inv_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _5870_/A vssd1 vssd1 vccd1 vccd1 _7766_/D sky130_fd_sc_hd__clkbuf_1
X_4821_ _4886_/A _4821_/B _4821_/C vssd1 vssd1 vccd1 vccd1 _4821_/X sky130_fd_sc_hd__or3_1
XFILLER_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4752_ _4654_/X _4751_/X _4951_/B vssd1 vssd1 vccd1 vccd1 _4752_/X sky130_fd_sc_hd__a21o_1
X_7540_ _7540_/A vssd1 vssd1 vccd1 vccd1 _8459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4683_ _8172_/Q _4683_/B vssd1 vssd1 vccd1 vccd1 _4801_/A sky130_fd_sc_hd__xnor2_1
XFILLER_119_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6422_ _6435_/A vssd1 vssd1 vccd1 vccd1 _6422_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6353_ _6398_/B _6461_/D vssd1 vssd1 vccd1 vccd1 _6395_/A sky130_fd_sc_hd__or2_1
XFILLER_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5304_ _5299_/X _5300_/X _5352_/B _5303_/X vssd1 vssd1 vccd1 vccd1 _5304_/X sky130_fd_sc_hd__a211o_1
X_6284_ _6465_/B vssd1 vssd1 vccd1 vccd1 _6284_/X sky130_fd_sc_hd__buf_2
XFILLER_115_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5235_ _5235_/A _5235_/B _5235_/C vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__or3_1
X_8023_ _8023_/CLK _8023_/D vssd1 vssd1 vccd1 vccd1 _8023_/Q sky130_fd_sc_hd__dfxtp_1
X_6781__366 _6782__367/A vssd1 vssd1 vccd1 vccd1 _8079_/CLK sky130_fd_sc_hd__inv_2
X_5166_ _8305_/Q _8297_/Q _8289_/Q _8313_/Q _5095_/X _5080_/A vssd1 vssd1 vccd1 vccd1
+ _5166_/X sky130_fd_sc_hd__mux4_1
X_5097_ _5215_/S vssd1 vssd1 vccd1 vccd1 _5318_/S sky130_fd_sc_hd__buf_2
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4117_ _8177_/Q vssd1 vssd1 vccd1 vccd1 _5622_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4048_ _4048_/A vssd1 vssd1 vccd1 vccd1 _8431_/D sky130_fd_sc_hd__clkbuf_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _6010_/A vssd1 vssd1 vccd1 vccd1 _6008_/B sky130_fd_sc_hd__clkbuf_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7807_ _8486_/CLK _7807_/D vssd1 vssd1 vccd1 vccd1 _7807_/Q sky130_fd_sc_hd__dfxtp_1
X_7738_ _7514_/A _7717_/A _7736_/X _7737_/X vssd1 vssd1 vccd1 vccd1 _8542_/D sky130_fd_sc_hd__o211a_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6636__299 _6637__300/A vssd1 vssd1 vccd1 vccd1 _7985_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5020_/A vssd1 vssd1 vccd1 vccd1 _8141_/D sky130_fd_sc_hd__clkbuf_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5922_ _5922_/A vssd1 vssd1 vccd1 vccd1 _5922_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5853_ _4163_/X _7773_/Q _5857_/S vssd1 vssd1 vccd1 vccd1 _5854_/A sky130_fd_sc_hd__mux2_1
X_5784_ _5784_/A vssd1 vssd1 vccd1 vccd1 _7847_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3651_ _7463_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3651_/X sky130_fd_sc_hd__clkbuf_16
X_4804_ _7977_/Q _8264_/Q _4915_/S vssd1 vssd1 vccd1 vccd1 _4804_/X sky130_fd_sc_hd__mux2_1
X_4735_ _4739_/S _4734_/X _4694_/X vssd1 vssd1 vccd1 vccd1 _4735_/X sky130_fd_sc_hd__a21o_1
X_7523_ _7523_/A _7523_/B _7523_/C _7523_/D vssd1 vssd1 vccd1 vccd1 _7524_/D sky130_fd_sc_hd__or4_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7462__175 _7462__175/A vssd1 vssd1 vccd1 vccd1 _8432_/CLK sky130_fd_sc_hd__inv_2
X_4666_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4666_/X sky130_fd_sc_hd__clkbuf_4
X_4597_ _4597_/A vssd1 vssd1 vccd1 vccd1 _8200_/D sky130_fd_sc_hd__clkbuf_1
X_6405_ _7861_/Q _6328_/A _6233_/X vssd1 vssd1 vccd1 vccd1 _6405_/X sky130_fd_sc_hd__a21o_1
X_7385_ _8370_/Q _7366_/A _7385_/S vssd1 vssd1 vccd1 vccd1 _7386_/A sky130_fd_sc_hd__mux2_1
X_6336_ _6382_/A vssd1 vssd1 vccd1 vccd1 _6336_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6267_ _7820_/Q _6266_/X _7737_/A vssd1 vssd1 vccd1 vccd1 _6273_/B sky130_fd_sc_hd__o21a_1
X_5218_ _8328_/Q _8049_/Q _5321_/S vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6198_ _6188_/X _7813_/Q _6191_/X _6195_/X _7781_/Q vssd1 vssd1 vccd1 vccd1 _7781_/D
+ sky130_fd_sc_hd__o32a_1
X_8006_ _8548_/CLK _8006_/D vssd1 vssd1 vccd1 vccd1 _8006_/Q sky130_fd_sc_hd__dfxtp_4
X_5149_ _8509_/Q _8258_/Q _8242_/Q _8282_/Q _5087_/X _5061_/A vssd1 vssd1 vccd1 vccd1
+ _5150_/B sky130_fd_sc_hd__mux4_2
XFILLER_72_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7145__70 _7145__70/A vssd1 vssd1 vccd1 vccd1 _8297_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_104 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_115 _4755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4520_ _8110_/Q vssd1 vssd1 vccd1 vccd1 _4520_/X sky130_fd_sc_hd__buf_4
X_4451_ _4379_/X _8259_/Q _4457_/S vssd1 vssd1 vccd1 vccd1 _4452_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4382_ _8493_/Q vssd1 vssd1 vccd1 vccd1 _4382_/X sky130_fd_sc_hd__buf_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ _6075_/A _6118_/X _6119_/X _6120_/X vssd1 vssd1 vccd1 vccd1 _6121_/X sky130_fd_sc_hd__o211a_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6052_ _6034_/X _6049_/X _6051_/X _6044_/X vssd1 vssd1 vccd1 vccd1 _6052_/X sky130_fd_sc_hd__o211a_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5003_ _5003_/A vssd1 vssd1 vccd1 vccd1 _8148_/D sky130_fd_sc_hd__clkbuf_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5905_ _5905_/A vssd1 vssd1 vccd1 vccd1 _5905_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5836_ _5836_/A vssd1 vssd1 vccd1 vccd1 _7824_/D sky130_fd_sc_hd__clkbuf_1
X_5767_ _7902_/Q _5575_/A _5767_/S vssd1 vssd1 vccd1 vccd1 _5768_/A sky130_fd_sc_hd__mux2_1
X_5698_ _5713_/S vssd1 vssd1 vccd1 vccd1 _5707_/S sky130_fd_sc_hd__buf_2
X_4718_ _4876_/A vssd1 vssd1 vccd1 vccd1 _4915_/S sky130_fd_sc_hd__buf_4
X_7506_ _6854_/A _7576_/A _7576_/B vssd1 vssd1 vccd1 vccd1 _7506_/X sky130_fd_sc_hd__and3b_1
X_8486_ _8486_/CLK _8486_/D vssd1 vssd1 vccd1 vccd1 _8486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4649_ _4649_/A vssd1 vssd1 vccd1 vccd1 _4649_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7368_ _8362_/Q _7377_/B vssd1 vssd1 vccd1 vccd1 _7368_/X sky130_fd_sc_hd__or2_1
XFILLER_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6748__345 _6748__345/A vssd1 vssd1 vccd1 vccd1 _8055_/CLK sky130_fd_sc_hd__inv_2
X_6980__440 _6980__440/A vssd1 vssd1 vccd1 vccd1 _8164_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7299_ _8534_/Q _7299_/B vssd1 vssd1 vccd1 vccd1 _7303_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8063_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7076__515 _7076__515/A vssd1 vssd1 vccd1 vccd1 _8242_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3247_ clkbuf_0__3247_/X vssd1 vssd1 vccd1 vccd1 _6544__239/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3951_ _3951_/A vssd1 vssd1 vccd1 vccd1 _8497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3451_ clkbuf_0__3451_/X vssd1 vssd1 vccd1 vccd1 _7083_/A sky130_fd_sc_hd__clkbuf_4
X_6670_ _5935_/A _8005_/Q _6670_/S vssd1 vssd1 vccd1 vccd1 _6671_/A sky130_fd_sc_hd__mux2_1
X_3882_ _7888_/Q _7889_/Q _7890_/Q _7887_/Q vssd1 vssd1 vccd1 vccd1 _7696_/D sky130_fd_sc_hd__or4b_1
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5621_ _5621_/A vssd1 vssd1 vccd1 vccd1 _7974_/D sky130_fd_sc_hd__clkbuf_1
X_8340_ _8340_/CLK _8340_/D vssd1 vssd1 vccd1 vccd1 _8340_/Q sky130_fd_sc_hd__dfxtp_1
X_5552_ _5387_/X _8022_/Q _5552_/S vssd1 vssd1 vccd1 vccd1 _5553_/A sky130_fd_sc_hd__mux2_1
X_8271_ _8271_/CLK _8271_/D vssd1 vssd1 vccd1 vccd1 _8271_/Q sky130_fd_sc_hd__dfxtp_1
X_4503_ _4503_/A vssd1 vssd1 vccd1 vccd1 _8239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5483_ _5498_/S vssd1 vssd1 vccd1 vccd1 _5492_/S sky130_fd_sc_hd__buf_2
XFILLER_117_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4434_ _4434_/A vssd1 vssd1 vccd1 vccd1 _8265_/D sky130_fd_sc_hd__clkbuf_1
X_7222_ _8545_/Q vssd1 vssd1 vccd1 vccd1 _7510_/A sky130_fd_sc_hd__inv_2
X_7153_ _7165_/A vssd1 vssd1 vccd1 vccd1 _7153_/X sky130_fd_sc_hd__buf_1
X_4365_ _4365_/A vssd1 vssd1 vccd1 vccd1 _8289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _7870_/Q input10/X _6111_/S vssd1 vssd1 vccd1 vccd1 _6104_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4296_ _4295_/X _8318_/Q _4299_/S vssd1 vssd1 vccd1 vccd1 _4297_/A sky130_fd_sc_hd__mux2_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6035_/A vssd1 vssd1 vccd1 vccd1 _6465_/B sky130_fd_sc_hd__clkbuf_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7986_ _7986_/CLK _7986_/D vssd1 vssd1 vccd1 vccd1 _7986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3649_ clkbuf_0__3649_/X vssd1 vssd1 vccd1 vccd1 _7456__170/A sky130_fd_sc_hd__clkbuf_4
X_5819_ _3978_/X _7831_/Q _5821_/S vssd1 vssd1 vccd1 vccd1 _5820_/A sky130_fd_sc_hd__mux2_1
X_8538_ _8540_/CLK _8538_/D vssd1 vssd1 vccd1 vccd1 _8538_/Q sky130_fd_sc_hd__dfxtp_1
X_6799_ _6802_/B _6799_/B vssd1 vssd1 vccd1 vccd1 _6800_/B sky130_fd_sc_hd__nand2_2
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8469_ _8473_/CLK _8469_/D vssd1 vssd1 vccd1 vccd1 _8469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3314_ clkbuf_0__3314_/X vssd1 vssd1 vccd1 vccd1 _6871_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_60_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput119 _6014_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[19] sky130_fd_sc_hd__buf_2
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput108 _7821_/Q vssd1 vssd1 vccd1 vccd1 caravel_uart_tx sky130_fd_sc_hd__buf_2
XFILLER_114_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4150_ _4150_/A vssd1 vssd1 vccd1 vccd1 _8402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4081_ _4081_/A vssd1 vssd1 vccd1 vccd1 _8418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7840_ _7840_/CLK _7840_/D vssd1 vssd1 vccd1 vccd1 _7840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7771_ _7771_/CLK _7771_/D vssd1 vssd1 vccd1 vccd1 _7771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4983_ _4983_/A vssd1 vssd1 vccd1 vccd1 _8157_/D sky130_fd_sc_hd__clkbuf_1
X_3934_ _3934_/A vssd1 vssd1 vccd1 vccd1 _8504_/D sky130_fd_sc_hd__clkbuf_1
X_6181__188 _6183__190/A vssd1 vssd1 vccd1 vccd1 _7775_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3434_ clkbuf_0__3434_/X vssd1 vssd1 vccd1 vccd1 _6974__435/A sky130_fd_sc_hd__clkbuf_4
X_3865_ _6417_/A _6517_/A vssd1 vssd1 vccd1 vccd1 _6326_/A sky130_fd_sc_hd__and2b_1
XFILLER_32_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5604_ _5554_/X _7981_/Q _5614_/S vssd1 vssd1 vccd1 vccd1 _5605_/A sky130_fd_sc_hd__mux2_1
X_8323_ _8323_/CLK _8323_/D vssd1 vssd1 vccd1 vccd1 _8323_/Q sky130_fd_sc_hd__dfxtp_1
X_5535_ _5535_/A vssd1 vssd1 vccd1 vccd1 _8030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5466_ _3954_/X _8061_/Q _5474_/S vssd1 vssd1 vccd1 vccd1 _5467_/A sky130_fd_sc_hd__mux2_1
X_8254_ _8254_/CLK _8254_/D vssd1 vssd1 vccd1 vccd1 _8254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3650_ clkbuf_0__3650_/X vssd1 vssd1 vccd1 vccd1 _7460__173/A sky130_fd_sc_hd__clkbuf_4
X_4417_ _4417_/A vssd1 vssd1 vccd1 vccd1 _8269_/D sky130_fd_sc_hd__clkbuf_1
X_7205_ _8538_/Q _7205_/B vssd1 vssd1 vccd1 vccd1 _7277_/C sky130_fd_sc_hd__xor2_1
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8185_ _8185_/CLK _8185_/D vssd1 vssd1 vccd1 vccd1 _8185_/Q sky130_fd_sc_hd__dfxtp_1
X_5397_ _5396_/X _8095_/Q _5402_/S vssd1 vssd1 vccd1 vccd1 _5398_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4348_ _4289_/X _8296_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4349_/A sky130_fd_sc_hd__mux2_1
X_4279_ _4279_/A vssd1 vssd1 vccd1 vccd1 _8324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6018_ _6018_/A vssd1 vssd1 vccd1 vccd1 _6018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7969_ _8527_/CLK _7969_/D vssd1 vssd1 vccd1 vccd1 _7969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7047__491 _7049__493/A vssd1 vssd1 vccd1 vccd1 _8218_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5320_ _8443_/Q _5232_/X _5230_/A _5318_/X _5319_/X vssd1 vssd1 vccd1 vccd1 _5320_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5251_ _5264_/A _5248_/X _5249_/X _5250_/X vssd1 vssd1 vccd1 vccd1 _5251_/X sky130_fd_sc_hd__o211a_1
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4202_ _4202_/A vssd1 vssd1 vccd1 vccd1 _8386_/D sky130_fd_sc_hd__clkbuf_1
X_5182_ _8115_/Q _5182_/B vssd1 vssd1 vccd1 vccd1 _5197_/A sky130_fd_sc_hd__or2_1
XFILLER_110_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4133_ _8177_/Q _8172_/Q vssd1 vssd1 vccd1 vccd1 _4627_/B sky130_fd_sc_hd__xnor2_2
X_4064_ _4015_/X _8424_/Q _4068_/S vssd1 vssd1 vccd1 vccd1 _4065_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7823_ _7823_/CLK _7823_/D vssd1 vssd1 vccd1 vccd1 _7823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7754_ _7754_/A _7754_/B vssd1 vssd1 vccd1 vccd1 _7754_/X sky130_fd_sc_hd__or2_1
X_4966_ _4966_/A vssd1 vssd1 vccd1 vccd1 _8164_/D sky130_fd_sc_hd__clkbuf_1
X_6705_ _6705_/A vssd1 vssd1 vccd1 vccd1 _8020_/D sky130_fd_sc_hd__clkbuf_1
X_4897_ _7934_/Q _4768_/A _4896_/X vssd1 vssd1 vccd1 vccd1 _4897_/Y sky130_fd_sc_hd__o21ai_1
X_3917_ _5787_/A _4490_/A vssd1 vssd1 vccd1 vccd1 _3933_/S sky130_fd_sc_hd__or2_2
X_7685_ _7687_/A _8520_/Q vssd1 vssd1 vccd1 vccd1 _7686_/A sky130_fd_sc_hd__and2_1
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3848_ _8121_/Q _8120_/Q _8119_/Q vssd1 vssd1 vccd1 vccd1 _3849_/B sky130_fd_sc_hd__and3_1
XFILLER_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5518_ _5661_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _5534_/S sky130_fd_sc_hd__or2_2
X_8306_ _8306_/CLK _8306_/D vssd1 vssd1 vccd1 vccd1 _8306_/Q sky130_fd_sc_hd__dfxtp_1
X_6498_ _8006_/Q _7891_/Q _6498_/S vssd1 vssd1 vccd1 vccd1 _6499_/A sky130_fd_sc_hd__mux2_1
X_5449_ _5449_/A vssd1 vssd1 vccd1 vccd1 _8072_/D sky130_fd_sc_hd__clkbuf_1
X_8237_ _8237_/CLK _8237_/D vssd1 vssd1 vccd1 vccd1 _8237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3247_ _6540_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3247_/X sky130_fd_sc_hd__clkbuf_16
X_8168_ _8168_/CLK _8168_/D vssd1 vssd1 vccd1 vccd1 _8168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8099_ _8099_/CLK _8099_/D vssd1 vssd1 vccd1 vccd1 _8099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4820_ _8093_/Q _4781_/A _4782_/A _4819_/X vssd1 vssd1 vccd1 vccd1 _4821_/C sky130_fd_sc_hd__o211a_1
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _8139_/Q _8026_/Q _7922_/Q _7906_/Q _4655_/X _4656_/X vssd1 vssd1 vccd1 vccd1
+ _4751_/X sky130_fd_sc_hd__mux4_1
X_7470_ _7482_/A vssd1 vssd1 vccd1 vccd1 _7470_/X sky130_fd_sc_hd__buf_1
X_4682_ _4654_/X _4678_/X _4681_/X vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__a21o_1
X_6421_ _7742_/B _7010_/B _6397_/X _7726_/A vssd1 vssd1 vccd1 vccd1 _6435_/A sky130_fd_sc_hd__a31o_2
XFILLER_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6352_ _6352_/A vssd1 vssd1 vccd1 vccd1 _6352_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5303_ _5306_/A _5301_/X _5302_/X _5250_/X vssd1 vssd1 vccd1 vccd1 _5303_/X sky130_fd_sc_hd__o211a_1
X_6283_ _8334_/Q _8333_/Q vssd1 vssd1 vccd1 vccd1 _7308_/A sky130_fd_sc_hd__nor2_2
X_5234_ _5230_/X _5231_/X _5233_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _5235_/C sky130_fd_sc_hd__o211a_1
X_8022_ _8022_/CLK _8022_/D vssd1 vssd1 vccd1 vccd1 _8022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5165_ _8423_/Q _8321_/Q _8058_/Q _8273_/Q _5129_/A _5305_/S vssd1 vssd1 vccd1 vccd1
+ _5165_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4116_ _8175_/Q vssd1 vssd1 vccd1 vccd1 _4933_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5096_ _8308_/Q _8300_/Q _8292_/Q _8316_/Q _5095_/X _5088_/X vssd1 vssd1 vccd1 vccd1
+ _5096_/X sky130_fd_sc_hd__mux4_1
X_4047_ _4019_/X _8431_/Q _4049_/S vssd1 vssd1 vccd1 vccd1 _4048_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7806_ _8486_/CLK _7806_/D vssd1 vssd1 vccd1 vccd1 _7806_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5998_/A vssd1 vssd1 vccd1 vccd1 _5998_/X sky130_fd_sc_hd__clkbuf_1
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7737_ _7737_/A vssd1 vssd1 vccd1 vccd1 _7737_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4949_ _4955_/A _4949_/B vssd1 vssd1 vccd1 vccd1 _4949_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6619_ _8185_/Q _6621_/B vssd1 vssd1 vccd1 vccd1 _6620_/A sky130_fd_sc_hd__and2_1
X_7599_ _6857_/A _7588_/X _7597_/X _7598_/X vssd1 vssd1 vccd1 vccd1 _7600_/B sky130_fd_sc_hd__o22a_1
XFILLER_106_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6944__411 _6946__413/A vssd1 vssd1 vccd1 vccd1 _8135_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5921_ _5921_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__or2_1
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5852_ _5852_/A vssd1 vssd1 vccd1 vccd1 _7774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5783_ _5572_/X _7847_/Q _5785_/S vssd1 vssd1 vccd1 vccd1 _5784_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3650_ _7457_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3650_/X sky130_fd_sc_hd__clkbuf_16
X_4803_ _4803_/A vssd1 vssd1 vccd1 vccd1 _4803_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4734_ _7768_/Q _7776_/Q _7851_/Q _7955_/Q _4666_/X _4667_/X vssd1 vssd1 vccd1 vccd1
+ _4734_/X sky130_fd_sc_hd__mux4_2
X_7522_ _7522_/A _7522_/B vssd1 vssd1 vccd1 vccd1 _7523_/D sky130_fd_sc_hd__and2_1
XFILLER_9_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4665_ _8220_/Q _8204_/Q _8166_/Q _8236_/Q _4810_/S _4649_/X vssd1 vssd1 vccd1 vccd1
+ _4665_/X sky130_fd_sc_hd__mux4_1
X_4596_ _4435_/X _8200_/Q _4596_/S vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__mux2_1
X_6404_ _7216_/A _6398_/Y _6403_/X _6397_/X vssd1 vssd1 vccd1 vccd1 _6404_/X sky130_fd_sc_hd__a22o_1
X_7384_ _8132_/Q _7364_/A _7366_/A _7383_/X _7286_/A vssd1 vssd1 vccd1 vccd1 _8369_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_115_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6335_ _6352_/A vssd1 vssd1 vccd1 vccd1 _6382_/A sky130_fd_sc_hd__buf_2
XFILLER_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6266_ _6095_/A _6465_/A _6082_/A _7819_/Q vssd1 vssd1 vccd1 vccd1 _6266_/X sky130_fd_sc_hd__a31o_1
X_8005_ _8537_/CLK _8005_/D vssd1 vssd1 vccd1 vccd1 _8005_/Q sky130_fd_sc_hd__dfxtp_4
X_5217_ _8515_/Q _5214_/X _5100_/A _5216_/X vssd1 vssd1 vccd1 vccd1 _5221_/B sky130_fd_sc_hd__o211a_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6197_ _6188_/X _7812_/Q _6191_/X _6195_/X _7780_/Q vssd1 vssd1 vccd1 vccd1 _7780_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5148_ _5146_/X _5147_/X _5205_/S vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5079_ _5250_/A vssd1 vssd1 vccd1 vccd1 _5079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_105 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_116 _5879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4450_ _4450_/A vssd1 vssd1 vccd1 vccd1 _8260_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4381_ _4381_/A vssd1 vssd1 vccd1 vccd1 _8283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6120_ _7633_/C vssd1 vssd1 vccd1 vccd1 _6120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _7781_/Q _6066_/B vssd1 vssd1 vccd1 vccd1 _6051_/X sky130_fd_sc_hd__or2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _8148_/Q _4517_/X _5006_/S vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__mux2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5904_ _7633_/B _5910_/B vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__or2_1
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6884_ _6890_/A vssd1 vssd1 vccd1 vccd1 _6884_/X sky130_fd_sc_hd__buf_1
X_5835_ _7824_/Q _5569_/A _5839_/S vssd1 vssd1 vccd1 vccd1 _5836_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5766_ _5766_/A vssd1 vssd1 vccd1 vccd1 _7903_/D sky130_fd_sc_hd__clkbuf_1
X_4717_ _8376_/Q _8266_/Q _7979_/Q _8400_/Q _4646_/X _4716_/X vssd1 vssd1 vccd1 vccd1
+ _4717_/X sky130_fd_sc_hd__mux4_2
X_5697_ _5751_/A _5823_/B vssd1 vssd1 vccd1 vccd1 _5713_/S sky130_fd_sc_hd__nor2_2
X_7505_ _7505_/A _8459_/Q vssd1 vssd1 vccd1 vccd1 _7505_/Y sky130_fd_sc_hd__nand2_1
X_8485_ _8486_/CLK _8485_/D vssd1 vssd1 vccd1 vccd1 _8485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4648_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4649_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4579_ _3975_/X _8207_/Q _4583_/S vssd1 vssd1 vccd1 vccd1 _4580_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7367_ _7383_/B vssd1 vssd1 vccd1 vccd1 _7377_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7298_ _7298_/A _8333_/Q vssd1 vssd1 vccd1 vccd1 _7299_/B sky130_fd_sc_hd__or2_2
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6249_ _6264_/S vssd1 vssd1 vccd1 vccd1 _6258_/S sky130_fd_sc_hd__buf_2
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7041__486 _7043__488/A vssd1 vssd1 vccd1 vccd1 _8213_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3315_ clkbuf_0__3315_/X vssd1 vssd1 vccd1 vccd1 _6766__354/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3246_ clkbuf_0__3246_/X vssd1 vssd1 vccd1 vccd1 _6539__235/A sky130_fd_sc_hd__clkbuf_4
X_8573__220 vssd1 vssd1 vccd1 vccd1 _8573__220/HI core0Index[7] sky130_fd_sc_hd__conb_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3950_ _3908_/X _8497_/Q _3952_/S vssd1 vssd1 vccd1 vccd1 _3951_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3450_ clkbuf_0__3450_/X vssd1 vssd1 vccd1 vccd1 _7057__500/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3881_ _7895_/Q _7896_/Q _7897_/Q _7898_/Q vssd1 vssd1 vccd1 vccd1 _7696_/C sky130_fd_sc_hd__or4_2
XFILLER_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5620_ _5575_/X _7974_/Q _5620_/S vssd1 vssd1 vccd1 vccd1 _5621_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5551_ _5551_/A vssd1 vssd1 vccd1 vccd1 _8023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4502_ _4391_/X _8239_/Q _4506_/S vssd1 vssd1 vccd1 vccd1 _4503_/A sky130_fd_sc_hd__mux2_1
X_8270_ _8270_/CLK _8270_/D vssd1 vssd1 vccd1 vccd1 _8270_/Q sky130_fd_sc_hd__dfxtp_1
X_5482_ _5482_/A _5787_/B vssd1 vssd1 vccd1 vccd1 _5498_/S sky130_fd_sc_hd__nor2_2
XFILLER_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7221_ _8541_/Q _7221_/B vssd1 vssd1 vccd1 vccd1 _7251_/B sky130_fd_sc_hd__xor2_1
X_4433_ _4432_/X _8265_/Q _4436_/S vssd1 vssd1 vccd1 vccd1 _4434_/A sky130_fd_sc_hd__mux2_1
X_7124__52 _7124__52/A vssd1 vssd1 vccd1 vccd1 _8279_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7152_ _7152_/A vssd1 vssd1 vccd1 vccd1 _7152_/X sky130_fd_sc_hd__buf_1
X_4364_ _4286_/X _8289_/Q _4366_/S vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4295_ _4295_/A vssd1 vssd1 vccd1 vccd1 _4295_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7083_ _7083_/A vssd1 vssd1 vccd1 vccd1 _7083_/X sky130_fd_sc_hd__buf_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6095_/X _6100_/X _6101_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6103_/X sky130_fd_sc_hd__o211a_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6075_/A vssd1 vssd1 vccd1 vccd1 _6034_/X sky130_fd_sc_hd__clkbuf_2
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7985_ _7985_/CLK _7985_/D vssd1 vssd1 vccd1 vccd1 _7985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3648_ clkbuf_0__3648_/X vssd1 vssd1 vccd1 vccd1 _7447__162/A sky130_fd_sc_hd__clkbuf_4
X_6867_ _7568_/A _7613_/A _6867_/C vssd1 vssd1 vccd1 vccd1 _8081_/D sky130_fd_sc_hd__nor3_1
X_5818_ _5818_/A vssd1 vssd1 vccd1 vccd1 _7832_/D sky130_fd_sc_hd__clkbuf_1
X_6798_ _8471_/Q _6804_/A _6830_/A _6824_/B _8472_/Q vssd1 vssd1 vccd1 vccd1 _6799_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6754__350 _6754__350/A vssd1 vssd1 vccd1 vccd1 _8060_/CLK sky130_fd_sc_hd__inv_2
X_5749_ _7910_/Q _5575_/A _5749_/S vssd1 vssd1 vccd1 vccd1 _5750_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8537_ _8537_/CLK _8537_/D vssd1 vssd1 vccd1 vccd1 _8537_/Q sky130_fd_sc_hd__dfxtp_2
X_8468_ _8473_/CLK _8468_/D vssd1 vssd1 vccd1 vccd1 _8468_/Q sky130_fd_sc_hd__dfxtp_1
X_8399_ _8399_/CLK _8399_/D vssd1 vssd1 vccd1 vccd1 _8399_/Q sky130_fd_sc_hd__dfxtp_1
X_7082__520 _7082__520/A vssd1 vssd1 vccd1 vccd1 _8247_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7666__42 _7666__42/A vssd1 vssd1 vccd1 vccd1 _8511_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6529__226 _6530__227/A vssd1 vssd1 vccd1 vccd1 _7904_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput109 _5972_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[0] sky130_fd_sc_hd__buf_2
XFILLER_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4080_ _4005_/X _8418_/Q _4088_/S vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7770_ _7770_/CLK _7770_/D vssd1 vssd1 vccd1 vccd1 _7770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4982_ _8157_/Q _4471_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4983_/A sky130_fd_sc_hd__mux2_1
X_3933_ _3911_/X _8504_/Q _3933_/S vssd1 vssd1 vccd1 vccd1 _3934_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _8530_/CLK sky130_fd_sc_hd__clkbuf_16
X_6652_ _6652_/A vssd1 vssd1 vccd1 vccd1 _6652_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3433_ clkbuf_0__3433_/X vssd1 vssd1 vccd1 vccd1 _6964__426/A sky130_fd_sc_hd__clkbuf_4
X_3864_ _7899_/Q vssd1 vssd1 vccd1 vccd1 _6517_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5603_ _5620_/S vssd1 vssd1 vccd1 vccd1 _5614_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6583_ _6583_/A vssd1 vssd1 vccd1 vccd1 _6583_/X sky130_fd_sc_hd__buf_1
X_8322_ _8322_/CLK _8322_/D vssd1 vssd1 vccd1 vccd1 _8322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5534_ _5387_/X _8030_/Q _5534_/S vssd1 vssd1 vccd1 vccd1 _5535_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5465_ _5480_/S vssd1 vssd1 vccd1 vccd1 _5474_/S sky130_fd_sc_hd__clkbuf_2
X_8253_ _8253_/CLK _8253_/D vssd1 vssd1 vccd1 vccd1 _8253_/Q sky130_fd_sc_hd__dfxtp_1
X_4416_ _4397_/X _8269_/Q _4416_/S vssd1 vssd1 vccd1 vccd1 _4417_/A sky130_fd_sc_hd__mux2_1
X_7204_ _8356_/Q _7257_/A vssd1 vssd1 vccd1 vccd1 _7205_/B sky130_fd_sc_hd__xnor2_1
X_8184_ _8184_/CLK _8184_/D vssd1 vssd1 vccd1 vccd1 _8184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5396_ _5396_/A vssd1 vssd1 vccd1 vccd1 _5396_/X sky130_fd_sc_hd__buf_4
XFILLER_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4347_ _4347_/A vssd1 vssd1 vccd1 vccd1 _8297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4278_ _4275_/X _8324_/Q _4290_/S vssd1 vssd1 vccd1 vccd1 _4279_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6017_ _8011_/Q _6019_/B vssd1 vssd1 vccd1 vccd1 _6018_/A sky130_fd_sc_hd__and2_1
XFILLER_67_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6305__206 _6306__207/A vssd1 vssd1 vccd1 vccd1 _7836_/CLK sky130_fd_sc_hd__inv_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7968_ _8527_/CLK _7968_/D vssd1 vssd1 vccd1 vccd1 _7968_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6919_ _6919_/A vssd1 vssd1 vccd1 vccd1 _6919_/X sky130_fd_sc_hd__buf_1
X_7899_ _8551_/CLK _7899_/D vssd1 vssd1 vccd1 vccd1 _7899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5250_ _5250_/A vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__buf_2
X_4201_ _8386_/Q _4172_/X _4209_/S vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5181_ _5181_/A _5182_/B vssd1 vssd1 vccd1 vccd1 _5183_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4132_ _8171_/Q _8176_/Q vssd1 vssd1 vccd1 vccd1 _4622_/B sky130_fd_sc_hd__and2b_1
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4063_ _4063_/A vssd1 vssd1 vccd1 vccd1 _8425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7660__37 _7660__37/A vssd1 vssd1 vccd1 vccd1 _8506_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7822_ _7822_/CLK _7822_/D vssd1 vssd1 vccd1 vccd1 _7822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4965_ _8164_/Q _4517_/X _4969_/S vssd1 vssd1 vccd1 vccd1 _4966_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7753_ _8547_/Q _7743_/X _7752_/X _7737_/X vssd1 vssd1 vccd1 vccd1 _8547_/D sky130_fd_sc_hd__o211a_1
X_3916_ _4301_/A _4076_/A _4301_/B vssd1 vssd1 vccd1 vccd1 _4490_/A sky130_fd_sc_hd__or3b_1
X_6704_ _8020_/Q _5967_/A _6706_/S vssd1 vssd1 vccd1 vccd1 _6705_/A sky130_fd_sc_hd__mux2_1
X_4896_ _8245_/Q _4781_/X _4803_/X _4895_/X _4782_/X vssd1 vssd1 vccd1 vccd1 _4896_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7684_ _7684_/A vssd1 vssd1 vccd1 vccd1 _8525_/D sky130_fd_sc_hd__clkbuf_1
X_3847_ _4057_/B _3845_/Y _3846_/Y vssd1 vssd1 vccd1 vccd1 _5035_/A sky130_fd_sc_hd__o21ai_1
X_5517_ _5517_/A vssd1 vssd1 vccd1 vccd1 _8038_/D sky130_fd_sc_hd__clkbuf_1
X_8305_ _8305_/CLK _8305_/D vssd1 vssd1 vccd1 vccd1 _8305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3315_ _6756_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3315_/X sky130_fd_sc_hd__clkbuf_16
X_8236_ _8236_/CLK _8236_/D vssd1 vssd1 vccd1 vccd1 _8236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6497_ _6497_/A vssd1 vssd1 vccd1 vccd1 _7890_/D sky130_fd_sc_hd__clkbuf_1
X_5448_ _8072_/Q _4172_/X _5456_/S vssd1 vssd1 vccd1 vccd1 _5449_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5379_ _5569_/A vssd1 vssd1 vccd1 vccd1 _5379_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__3246_ _6534_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3246_/X sky130_fd_sc_hd__clkbuf_16
X_8167_ _8527_/CLK _8167_/D vssd1 vssd1 vccd1 vccd1 _8167_/Q sky130_fd_sc_hd__dfxtp_1
X_8098_ _8098_/CLK _8098_/D vssd1 vssd1 vccd1 vccd1 _8098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7485__18 _7485__18/A vssd1 vssd1 vccd1 vccd1 _8450_/CLK sky130_fd_sc_hd__inv_2
XFILLER_88_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7095__530 _7095__530/A vssd1 vssd1 vccd1 vccd1 _8257_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8553__251 vssd1 vssd1 vccd1 vccd1 partID[0] _8553__251/LO sky130_fd_sc_hd__conb_1
XFILLER_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4750_ _8094_/Q _8086_/Q _7914_/Q _8155_/Q _4646_/X _4716_/X vssd1 vssd1 vccd1 vccd1
+ _4750_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4681_ _4677_/S _4679_/X _4886_/A vssd1 vssd1 vccd1 vccd1 _4681_/X sky130_fd_sc_hd__a21o_1
X_6420_ _7514_/A _6434_/B _6431_/C vssd1 vssd1 vccd1 vccd1 _6420_/X sky130_fd_sc_hd__and3_1
X_6351_ _8062_/Q vssd1 vssd1 vccd1 vccd1 _7741_/A sky130_fd_sc_hd__clkbuf_2
X_5302_ _8277_/Q _5180_/X _5198_/X _8504_/Q vssd1 vssd1 vccd1 vccd1 _5302_/X sky130_fd_sc_hd__o22a_1
XFILLER_6_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6282_ _8361_/Q _6278_/X _6280_/X _7355_/A vssd1 vssd1 vccd1 vccd1 _6282_/X sky130_fd_sc_hd__a211o_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5233_ _8279_/Q _5232_/X _5214_/X _8506_/Q vssd1 vssd1 vccd1 vccd1 _5233_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8021_ _8486_/CLK _8021_/D vssd1 vssd1 vccd1 vccd1 _8021_/Q sky130_fd_sc_hd__dfxtp_1
X_5164_ _5055_/A _5161_/X _5163_/X vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__a21o_1
X_7104__537 _7107__540/A vssd1 vssd1 vccd1 vccd1 _8264_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4115_ _8176_/Q vssd1 vssd1 vccd1 vccd1 _4466_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5095_ _5215_/S vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__clkbuf_4
X_4046_ _4046_/A vssd1 vssd1 vccd1 vccd1 _8432_/D sky130_fd_sc_hd__clkbuf_1
X_7469__5 _7469__5/A vssd1 vssd1 vccd1 vccd1 _8437_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7805_ _8487_/CLK _7805_/D vssd1 vssd1 vccd1 vccd1 _7805_/Q sky130_fd_sc_hd__dfxtp_1
X_5997_ _5997_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5998_/A sky130_fd_sc_hd__and2_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7736_ _5921_/A _7731_/X _7723_/X vssd1 vssd1 vccd1 vccd1 _7736_/X sky130_fd_sc_hd__a21bo_1
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4948_ _4948_/A vssd1 vssd1 vccd1 vccd1 _4955_/A sky130_fd_sc_hd__clkbuf_2
X_4879_ _4803_/X _4877_/X _4878_/X _4782_/X vssd1 vssd1 vccd1 vccd1 _4879_/X sky130_fd_sc_hd__o211a_1
X_6618_ _6618_/A vssd1 vssd1 vccd1 vccd1 _7971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7598_ _7598_/A _7588_/A vssd1 vssd1 vccd1 vccd1 _7598_/X sky130_fd_sc_hd__or2b_1
XFILLER_118_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8219_ _8219_/CLK _8219_/D vssd1 vssd1 vccd1 vccd1 _8219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3477_ clkbuf_0__3477_/X vssd1 vssd1 vccd1 vccd1 _7186__102/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7409__131 _7411__133/A vssd1 vssd1 vccd1 vccd1 _8388_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5920_ _5920_/A vssd1 vssd1 vccd1 vccd1 _5920_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5851_ _4160_/X _7774_/Q _5851_/S vssd1 vssd1 vccd1 vccd1 _5852_/A sky130_fd_sc_hd__mux2_1
X_8590__237 vssd1 vssd1 vccd1 vccd1 _8590__237/HI manufacturerID[9] sky130_fd_sc_hd__conb_1
X_5782_ _5782_/A vssd1 vssd1 vccd1 vccd1 _7848_/D sky130_fd_sc_hd__clkbuf_1
X_4802_ _4673_/X _4779_/X _4789_/X _4800_/X _4949_/B vssd1 vssd1 vccd1 vccd1 _4802_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4733_ _4733_/A vssd1 vssd1 vccd1 vccd1 _4739_/S sky130_fd_sc_hd__clkbuf_2
X_7521_ _8547_/Q _7521_/B vssd1 vssd1 vccd1 vccd1 _7523_/C sky130_fd_sc_hd__xnor2_1
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4664_ _4760_/S vssd1 vssd1 vccd1 vccd1 _4664_/X sky130_fd_sc_hd__clkbuf_2
X_6403_ _7747_/A _7973_/Q _6410_/C _7010_/B vssd1 vssd1 vccd1 vccd1 _6403_/X sky130_fd_sc_hd__a31o_1
X_4595_ _4595_/A vssd1 vssd1 vccd1 vccd1 _8201_/D sky130_fd_sc_hd__clkbuf_1
X_7383_ _8369_/Q _7383_/B vssd1 vssd1 vccd1 vccd1 _7383_/X sky130_fd_sc_hd__or2_1
X_6334_ _6362_/A vssd1 vssd1 vccd1 vccd1 _7747_/A sky130_fd_sc_hd__clkbuf_2
X_7471__6 _7472__7/A vssd1 vssd1 vccd1 vccd1 _8438_/CLK sky130_fd_sc_hd__inv_2
X_6265_ _6265_/A vssd1 vssd1 vccd1 vccd1 _7818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5216_ _8499_/Q _5063_/B _5215_/X _5192_/A vssd1 vssd1 vccd1 vccd1 _5216_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8004_ _8537_/CLK _8004_/D vssd1 vssd1 vccd1 vccd1 _8004_/Q sky130_fd_sc_hd__dfxtp_1
X_6196_ _6188_/X _7811_/Q _6191_/X _6195_/X _7779_/Q vssd1 vssd1 vccd1 vccd1 _7779_/D
+ sky130_fd_sc_hd__o32a_1
X_5147_ _8306_/Q _8298_/Q _8290_/Q _8314_/Q _5095_/X _5088_/X vssd1 vssd1 vccd1 vccd1
+ _5147_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5078_ _8410_/Q _8394_/Q _8386_/Q _8418_/Q _5273_/S _5068_/X vssd1 vssd1 vccd1 vccd1
+ _5078_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4029_ _4029_/A vssd1 vssd1 vccd1 vccd1 _8437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7719_ _7719_/A vssd1 vssd1 vccd1 vccd1 _7719_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6764__352 _6767__355/A vssd1 vssd1 vccd1 vccd1 _8065_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_106 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_117 _6367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6578__266 _6579__267/A vssd1 vssd1 vccd1 vccd1 _7944_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4380_ _4379_/X _8283_/Q _4389_/S vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7151__75 _7151__75/A vssd1 vssd1 vccd1 vccd1 _8302_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6138_/A vssd1 vssd1 vccd1 vccd1 _6066_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5001_/A vssd1 vssd1 vccd1 vccd1 _8149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5903_ _5903_/A vssd1 vssd1 vccd1 vccd1 _7633_/B sky130_fd_sc_hd__buf_6
X_5834_ _5834_/A vssd1 vssd1 vccd1 vccd1 _7825_/D sky130_fd_sc_hd__clkbuf_1
X_5765_ _7903_/Q _5572_/A _5767_/S vssd1 vssd1 vccd1 vccd1 _5766_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4716_ _4716_/A vssd1 vssd1 vccd1 vccd1 _4716_/X sky130_fd_sc_hd__buf_4
X_5696_ _5696_/A vssd1 vssd1 vccd1 vccd1 _7934_/D sky130_fd_sc_hd__clkbuf_1
X_7504_ _7609_/A _7609_/B _7499_/X _7541_/A _7503_/X vssd1 vssd1 vccd1 vccd1 _7504_/X
+ sky130_fd_sc_hd__o221a_1
X_8484_ _8486_/CLK _8484_/D vssd1 vssd1 vccd1 vccd1 _8484_/Q sky130_fd_sc_hd__dfxtp_1
X_4647_ _4767_/A vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__buf_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7366_ _7366_/A vssd1 vssd1 vccd1 vccd1 _7366_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4578_ _4578_/A vssd1 vssd1 vccd1 vccd1 _8208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6248_ _6248_/A _6690_/B vssd1 vssd1 vccd1 vccd1 _6264_/S sky130_fd_sc_hd__nand2_1
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3245_ clkbuf_0__3245_/X vssd1 vssd1 vccd1 vccd1 _6533__230/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6957__422 _6957__422/A vssd1 vssd1 vccd1 vccd1 _8146_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3880_ _7891_/Q _7892_/Q _7893_/Q _7894_/Q vssd1 vssd1 vccd1 vccd1 _7696_/B sky130_fd_sc_hd__or4_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5550_ _5383_/X _8023_/Q _5552_/S vssd1 vssd1 vccd1 vccd1 _5551_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5481_ _5481_/A vssd1 vssd1 vccd1 vccd1 _8054_/D sky130_fd_sc_hd__clkbuf_1
X_4501_ _4501_/A vssd1 vssd1 vccd1 vccd1 _8240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4432_ _5399_/A vssd1 vssd1 vccd1 vccd1 _4432_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7220_ _7220_/A _7220_/B vssd1 vssd1 vccd1 vccd1 _7221_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6964__426 _6964__426/A vssd1 vssd1 vccd1 vccd1 _8150_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4363_ _4363_/A vssd1 vssd1 vccd1 vccd1 _8290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4294_ _4294_/A vssd1 vssd1 vccd1 vccd1 _8319_/D sky130_fd_sc_hd__clkbuf_1
X_6102_ _7633_/C vssd1 vssd1 vccd1 vccd1 _6102_/X sky130_fd_sc_hd__clkbuf_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _6095_/A vssd1 vssd1 vccd1 vccd1 _6075_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8596__243 vssd1 vssd1 vccd1 vccd1 _8596__243/HI partID[9] sky130_fd_sc_hd__conb_1
XFILLER_82_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7984_ _7984_/CLK _7984_/D vssd1 vssd1 vccd1 vccd1 _7984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3647_ clkbuf_0__3647_/X vssd1 vssd1 vccd1 vccd1 _7444__160/A sky130_fd_sc_hd__clkbuf_4
X_7388__115 _7388__115/A vssd1 vssd1 vccd1 vccd1 _8372_/CLK sky130_fd_sc_hd__inv_2
X_6897__391 _6897__391/A vssd1 vssd1 vccd1 vccd1 _8105_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6866_ _8479_/Q _7606_/B vssd1 vssd1 vccd1 vccd1 _6867_/C sky130_fd_sc_hd__nand2_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5817_ _3975_/X _7832_/Q _5821_/S vssd1 vssd1 vccd1 vccd1 _5818_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6797_ _8470_/Q _8469_/Q vssd1 vssd1 vccd1 vccd1 _6804_/A sky130_fd_sc_hd__and2_1
X_5748_ _5748_/A vssd1 vssd1 vccd1 vccd1 _7911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8536_ _8537_/CLK _8536_/D vssd1 vssd1 vccd1 vccd1 _8536_/Q sky130_fd_sc_hd__dfxtp_1
X_5679_ _5751_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _5695_/S sky130_fd_sc_hd__nor2_2
X_8467_ _8473_/CLK _8467_/D vssd1 vssd1 vccd1 vccd1 _8467_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3477_ _7184_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3477_/X sky130_fd_sc_hd__clkbuf_16
X_8398_ _8398_/CLK _8398_/D vssd1 vssd1 vccd1 vccd1 _8398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7349_ _7356_/B vssd1 vssd1 vccd1 vccd1 _7354_/A sky130_fd_sc_hd__inv_2
XFILLER_103_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _4981_/A vssd1 vssd1 vccd1 vccd1 _8158_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__3655_ clkbuf_0__3655_/X vssd1 vssd1 vccd1 vccd1 _7485__18/A sky130_fd_sc_hd__clkbuf_16
X_3932_ _3932_/A vssd1 vssd1 vccd1 vccd1 _8505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3432_ clkbuf_0__3432_/X vssd1 vssd1 vccd1 vccd1 _6975_/A sky130_fd_sc_hd__clkbuf_4
X_3863_ _7900_/Q vssd1 vssd1 vccd1 vccd1 _6417_/A sky130_fd_sc_hd__clkbuf_1
X_5602_ _5602_/A _5769_/A vssd1 vssd1 vccd1 vccd1 _5620_/S sky130_fd_sc_hd__or2_2
X_6296__200 _6296__200/A vssd1 vssd1 vccd1 vccd1 _7830_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5533_ _5533_/A vssd1 vssd1 vccd1 vccd1 _8031_/D sky130_fd_sc_hd__clkbuf_1
X_8321_ _8321_/CLK _8321_/D vssd1 vssd1 vccd1 vccd1 _8321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8252_ _8252_/CLK _8252_/D vssd1 vssd1 vccd1 vccd1 _8252_/Q sky130_fd_sc_hd__dfxtp_1
X_5464_ _5464_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _5480_/S sky130_fd_sc_hd__or2_2
X_4415_ _4415_/A vssd1 vssd1 vccd1 vccd1 _8270_/D sky130_fd_sc_hd__clkbuf_1
X_7203_ _7199_/A _7344_/B _8537_/Q vssd1 vssd1 vccd1 vccd1 _7207_/A sky130_fd_sc_hd__a21bo_1
X_5395_ _5395_/A vssd1 vssd1 vccd1 vccd1 _8096_/D sky130_fd_sc_hd__clkbuf_1
X_8183_ _8183_/CLK _8183_/D vssd1 vssd1 vccd1 vccd1 _8183_/Q sky130_fd_sc_hd__dfxtp_1
X_4346_ _4286_/X _8297_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__mux2_1
X_7134_ _7146_/A vssd1 vssd1 vccd1 vccd1 _7134_/X sky130_fd_sc_hd__buf_1
XFILLER_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4277_ _4299_/S vssd1 vssd1 vccd1 vccd1 _4290_/S sky130_fd_sc_hd__clkbuf_2
X_7065_ _7077_/A vssd1 vssd1 vccd1 vccd1 _7065_/X sky130_fd_sc_hd__buf_1
X_6016_ _6016_/A vssd1 vssd1 vccd1 vccd1 _6016_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7967_ _8527_/CLK _7967_/D vssd1 vssd1 vccd1 vccd1 _7967_/Q sky130_fd_sc_hd__dfxtp_1
X_7898_ _8531_/CLK _7898_/D vssd1 vssd1 vccd1 vccd1 _7898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6849_ _8465_/Q _6849_/B vssd1 vssd1 vccd1 vccd1 _7522_/B sky130_fd_sc_hd__xnor2_4
XFILLER_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8519_ _8519_/CLK _8519_/D vssd1 vssd1 vccd1 vccd1 _8519_/Q sky130_fd_sc_hd__dfxtp_1
X_6535__231 _6539__235/A vssd1 vssd1 vccd1 vccd1 _7909_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7403__126 _7405__128/A vssd1 vssd1 vccd1 vccd1 _8383_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7054__497 _7054__497/A vssd1 vssd1 vccd1 vccd1 _8224_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4200_ _4215_/S vssd1 vssd1 vccd1 vccd1 _4209_/S sky130_fd_sc_hd__buf_2
X_5180_ _5232_/A vssd1 vssd1 vccd1 vccd1 _5180_/X sky130_fd_sc_hd__buf_2
X_7458__171 _7460__173/A vssd1 vssd1 vccd1 vccd1 _8428_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4131_ _4627_/C _4131_/B _4125_/A vssd1 vssd1 vccd1 vccd1 _4131_/X sky130_fd_sc_hd__or3b_1
XFILLER_110_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4062_ _4011_/X _8425_/Q _4068_/S vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7821_ _8486_/CLK _7821_/D vssd1 vssd1 vccd1 vccd1 _7821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7752_ _7640_/A _7702_/A _7744_/X vssd1 vssd1 vccd1 vccd1 _7752_/X sky130_fd_sc_hd__a21bo_1
X_4964_ _4964_/A vssd1 vssd1 vccd1 vccd1 _8165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3915_ _4057_/B vssd1 vssd1 vccd1 vccd1 _4301_/B sky130_fd_sc_hd__clkbuf_2
X_6703_ _6703_/A vssd1 vssd1 vccd1 vccd1 _8019_/D sky130_fd_sc_hd__clkbuf_1
X_4895_ _7982_/Q _8030_/Q _4901_/S vssd1 vssd1 vccd1 vccd1 _4895_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7683_ _7687_/A _8167_/Q vssd1 vssd1 vccd1 vccd1 _7684_/A sky130_fd_sc_hd__and2_1
X_3846_ _8123_/Q _8118_/Q vssd1 vssd1 vccd1 vccd1 _3846_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6565_ _6571_/A vssd1 vssd1 vccd1 vccd1 _6565_/X sky130_fd_sc_hd__buf_1
XFILLER_118_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5516_ _8038_/Q _4298_/A _5516_/S vssd1 vssd1 vccd1 vccd1 _5517_/A sky130_fd_sc_hd__mux2_1
X_8304_ _8304_/CLK _8304_/D vssd1 vssd1 vccd1 vccd1 _8304_/Q sky130_fd_sc_hd__dfxtp_1
X_6496_ _8005_/Q _7890_/Q _6498_/S vssd1 vssd1 vccd1 vccd1 _6497_/A sky130_fd_sc_hd__mux2_1
X_5447_ _5462_/S vssd1 vssd1 vccd1 vccd1 _5456_/S sky130_fd_sc_hd__buf_2
Xclkbuf_0__3314_ _6755_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3314_/X sky130_fd_sc_hd__clkbuf_16
X_8235_ _8235_/CLK _8235_/D vssd1 vssd1 vccd1 vccd1 _8235_/Q sky130_fd_sc_hd__dfxtp_1
X_5378_ _8108_/Q vssd1 vssd1 vccd1 vccd1 _5569_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3245_ _6528_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3245_/X sky130_fd_sc_hd__clkbuf_16
X_8166_ _8166_/CLK _8166_/D vssd1 vssd1 vccd1 vccd1 _8166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6311__211 _6312__212/A vssd1 vssd1 vccd1 vccd1 _7841_/CLK sky130_fd_sc_hd__inv_2
X_4329_ _4329_/A vssd1 vssd1 vccd1 vccd1 _8305_/D sky130_fd_sc_hd__clkbuf_1
X_8097_ _8097_/CLK _8097_/D vssd1 vssd1 vccd1 vccd1 _8097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ _4694_/A vssd1 vssd1 vccd1 vccd1 _4886_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6350_ _6397_/B vssd1 vssd1 vccd1 vccd1 _6350_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5301_ _8237_/Q _8253_/Q _5315_/S vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__mux2_1
X_6281_ _8333_/Q vssd1 vssd1 vccd1 vccd1 _7355_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5232_ _5232_/A vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__buf_2
X_8020_ _8486_/CLK _8020_/D vssd1 vssd1 vccd1 vccd1 _8020_/Q sky130_fd_sc_hd__dfxtp_1
X_5163_ _5079_/X _5162_/X _5131_/X vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4114_ _8113_/Q vssd1 vssd1 vccd1 vccd1 _4114_/X sky130_fd_sc_hd__buf_2
XFILLER_83_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5094_ _5092_/X _5093_/X _5221_/A vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4045_ _4015_/X _8432_/Q _4049_/S vssd1 vssd1 vccd1 vccd1 _4046_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7804_ _8487_/CLK _7804_/D vssd1 vssd1 vccd1 vccd1 _7804_/Q sky130_fd_sc_hd__dfxtp_1
X_5996_ _5996_/A vssd1 vssd1 vccd1 vccd1 _5996_/X sky130_fd_sc_hd__clkbuf_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7735_ _7529_/A _7717_/X _7734_/X _7719_/X vssd1 vssd1 vccd1 vccd1 _8541_/D sky130_fd_sc_hd__o211a_1
X_4947_ _4947_/A vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__clkbuf_2
X_4878_ _8396_/Q _4805_/Y _4806_/X _8372_/Q vssd1 vssd1 vccd1 vccd1 _4878_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6617_ _8184_/Q _6621_/B vssd1 vssd1 vccd1 vccd1 _6618_/A sky130_fd_sc_hd__and2_1
X_7597_ _7505_/A _6860_/X _7550_/C vssd1 vssd1 vccd1 vccd1 _7597_/X sky130_fd_sc_hd__o21ba_1
X_6479_ _5986_/A _7882_/Q _6487_/S vssd1 vssd1 vccd1 vccd1 _6480_/A sky130_fd_sc_hd__mux2_1
X_8218_ _8218_/CLK _8218_/D vssd1 vssd1 vccd1 vccd1 _8218_/Q sky130_fd_sc_hd__dfxtp_1
X_8149_ _8149_/CLK _8149_/D vssd1 vssd1 vccd1 vccd1 _8149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_0 _7821_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7490__22 _7490__22/A vssd1 vssd1 vccd1 vccd1 _8454_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3476_ clkbuf_0__3476_/X vssd1 vssd1 vccd1 vccd1 _7395_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6951__417 _6952__418/A vssd1 vssd1 vccd1 vccd1 _8141_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6318__217 _6318__217/A vssd1 vssd1 vccd1 vccd1 _7847_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7163__84 _7163__84/A vssd1 vssd1 vccd1 vccd1 _8311_/CLK sky130_fd_sc_hd__inv_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5850_ _5850_/A vssd1 vssd1 vccd1 vccd1 _7775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5781_ _5569_/X _7848_/Q _5785_/S vssd1 vssd1 vccd1 vccd1 _5782_/A sky130_fd_sc_hd__mux2_1
X_4801_ _4801_/A vssd1 vssd1 vccd1 vccd1 _4949_/B sky130_fd_sc_hd__buf_2
X_6891__386 _6892__387/A vssd1 vssd1 vccd1 vccd1 _8100_/CLK sky130_fd_sc_hd__inv_2
X_4732_ _4732_/A vssd1 vssd1 vccd1 vccd1 _4733_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7520_ _7522_/A _7522_/B vssd1 vssd1 vccd1 vccd1 _7523_/B sky130_fd_sc_hd__nor2_1
X_7451_ _7457_/A vssd1 vssd1 vccd1 vccd1 _7451_/X sky130_fd_sc_hd__buf_1
X_7110__542 _7113__545/A vssd1 vssd1 vccd1 vccd1 _8269_/CLK sky130_fd_sc_hd__inv_2
X_4663_ _4663_/A vssd1 vssd1 vccd1 vccd1 _4760_/S sky130_fd_sc_hd__clkbuf_4
X_6402_ _8544_/Q vssd1 vssd1 vccd1 vccd1 _7216_/A sky130_fd_sc_hd__buf_2
X_4594_ _4432_/X _8201_/Q _4596_/S vssd1 vssd1 vccd1 vccd1 _4595_/A sky130_fd_sc_hd__mux2_1
X_7382_ _8131_/Q _7364_/A _7366_/A _7381_/X _7286_/A vssd1 vssd1 vccd1 vccd1 _8368_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6333_ _8062_/Q vssd1 vssd1 vccd1 vccd1 _6362_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6264_ _7646_/A _7818_/Q _6264_/S vssd1 vssd1 vccd1 vccd1 _6265_/A sky130_fd_sc_hd__mux2_1
X_5215_ _8041_/Q _8068_/Q _5215_/S vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__mux2_1
X_8003_ _8540_/CLK _8003_/D vssd1 vssd1 vccd1 vccd1 _8003_/Q sky130_fd_sc_hd__dfxtp_1
X_6195_ _6213_/A vssd1 vssd1 vccd1 vccd1 _6195_/X sky130_fd_sc_hd__clkbuf_2
X_5146_ _8424_/Q _8322_/Q _8059_/Q _8274_/Q _5129_/A _5305_/S vssd1 vssd1 vccd1 vccd1
+ _5146_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5077_ _5321_/S vssd1 vssd1 vccd1 vccd1 _5273_/S sky130_fd_sc_hd__buf_4
XFILLER_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4028_ _4027_/X _8437_/Q _4036_/S vssd1 vssd1 vccd1 vccd1 _4029_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5979_ _5979_/A vssd1 vssd1 vccd1 vccd1 _5979_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7718_ _5935_/A _7710_/X _7717_/A vssd1 vssd1 vccd1 vccd1 _7718_/X sky130_fd_sc_hd__a21bo_1
XFILLER_100_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7011__462 _7011__462/A vssd1 vssd1 vccd1 vccd1 _8189_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_107 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_0__3459_ clkbuf_0__3459_/X vssd1 vssd1 vccd1 vccd1 _7099__533/A sky130_fd_sc_hd__clkbuf_4
XINSDIODE2_118 _6202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7136__62 _7136__62/A vssd1 vssd1 vccd1 vccd1 _8289_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _8149_/Q _4471_/X _5006_/S vssd1 vssd1 vccd1 vccd1 _5001_/A sky130_fd_sc_hd__mux2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5902_ _5902_/A vssd1 vssd1 vccd1 vccd1 _5902_/X sky130_fd_sc_hd__clkbuf_1
X_5833_ _7825_/Q _5566_/A _5833_/S vssd1 vssd1 vccd1 vccd1 _5834_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5764_ _5764_/A vssd1 vssd1 vccd1 vccd1 _7904_/D sky130_fd_sc_hd__clkbuf_1
X_7503_ _8460_/Q _8459_/Q _7503_/C vssd1 vssd1 vccd1 vccd1 _7503_/X sky130_fd_sc_hd__or3_1
X_4715_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__buf_2
X_5695_ _7934_/Q _5599_/X _5695_/S vssd1 vssd1 vccd1 vccd1 _5696_/A sky130_fd_sc_hd__mux2_1
X_8483_ _8486_/CLK _8483_/D vssd1 vssd1 vccd1 vccd1 _8483_/Q sky130_fd_sc_hd__dfxtp_1
X_4646_ _4646_/A vssd1 vssd1 vccd1 vccd1 _4646_/X sky130_fd_sc_hd__buf_4
X_4577_ _3972_/X _8208_/Q _4577_/S vssd1 vssd1 vccd1 vccd1 _4578_/A sky130_fd_sc_hd__mux2_1
X_7365_ _7365_/A vssd1 vssd1 vccd1 vccd1 _7366_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6316_ _6322_/A vssd1 vssd1 vccd1 vccd1 _6316_/X sky130_fd_sc_hd__buf_1
XFILLER_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6247_ _6247_/A _6272_/B vssd1 vssd1 vccd1 vccd1 _6690_/B sky130_fd_sc_hd__nor2_4
X_6178_ _6184_/A vssd1 vssd1 vccd1 vccd1 _6178_/X sky130_fd_sc_hd__buf_1
XFILLER_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5129_ _5129_/A vssd1 vssd1 vccd1 vccd1 _5129_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3313_ clkbuf_0__3313_/X vssd1 vssd1 vccd1 vccd1 _6753__349/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3244_ clkbuf_0__3244_/X vssd1 vssd1 vccd1 vccd1 _6540_/A sky130_fd_sc_hd__clkbuf_4
X_7117__548 _7118__549/A vssd1 vssd1 vccd1 vccd1 _8275_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6584__271 _6584__271/A vssd1 vssd1 vccd1 vccd1 _7949_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7452__166 _7453__167/A vssd1 vssd1 vccd1 vccd1 _8423_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6625__290 _6625__290/A vssd1 vssd1 vccd1 vccd1 _7976_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7018__468 _7019__469/A vssd1 vssd1 vccd1 vccd1 _8195_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5480_ _3981_/X _8054_/Q _5480_/S vssd1 vssd1 vccd1 vccd1 _5481_/A sky130_fd_sc_hd__mux2_1
X_4500_ _4388_/X _8240_/Q _4500_/S vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4431_ _8110_/Q vssd1 vssd1 vccd1 vccd1 _5399_/A sky130_fd_sc_hd__buf_4
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4362_ _4283_/X _8290_/Q _4366_/S vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4293_ _4292_/X _8319_/Q _4299_/S vssd1 vssd1 vccd1 vccd1 _4294_/A sky130_fd_sc_hd__mux2_1
X_6101_ _7794_/Q _6105_/B vssd1 vssd1 vccd1 vccd1 _6101_/X sky130_fd_sc_hd__or2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6108_/A vssd1 vssd1 vccd1 vccd1 _6095_/A sky130_fd_sc_hd__clkinv_2
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7983_ _7983_/CLK _7983_/D vssd1 vssd1 vccd1 vccd1 _7983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3646_ clkbuf_0__3646_/X vssd1 vssd1 vccd1 vccd1 _7436__153/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6865_ _6865_/A _6865_/B vssd1 vssd1 vccd1 vccd1 _7606_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5816_ _5816_/A vssd1 vssd1 vccd1 vccd1 _7833_/D sky130_fd_sc_hd__clkbuf_1
X_6796_ _6796_/A _6830_/A _6824_/B vssd1 vssd1 vccd1 vccd1 _6802_/B sky130_fd_sc_hd__nand3_4
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5747_ _7911_/Q _5572_/A _5749_/S vssd1 vssd1 vccd1 vccd1 _5748_/A sky130_fd_sc_hd__mux2_1
X_8535_ _8548_/CLK _8535_/D vssd1 vssd1 vccd1 vccd1 _8535_/Q sky130_fd_sc_hd__dfxtp_1
X_8466_ _8473_/CLK _8466_/D vssd1 vssd1 vccd1 vccd1 _8466_/Q sky130_fd_sc_hd__dfxtp_1
X_5678_ _5678_/A vssd1 vssd1 vccd1 vccd1 _7942_/D sky130_fd_sc_hd__clkbuf_1
X_8397_ _8397_/CLK _8397_/D vssd1 vssd1 vccd1 vccd1 _8397_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3476_ _7183_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3476_/X sky130_fd_sc_hd__clkbuf_16
X_4629_ _4764_/B vssd1 vssd1 vccd1 vccd1 _4629_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7348_ _7348_/A _7348_/B vssd1 vssd1 vccd1 vccd1 _8358_/D sky130_fd_sc_hd__nor2_1
X_7279_ _7344_/A _7344_/B _6440_/A vssd1 vssd1 vccd1 vccd1 _7279_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7130__57 _7130__57/A vssd1 vssd1 vccd1 vccd1 _8284_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3089_ clkbuf_0__3089_/X vssd1 vssd1 vccd1 vccd1 _6306__207/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6924__400 _6924__400/A vssd1 vssd1 vccd1 vccd1 _8122_/CLK sky130_fd_sc_hd__inv_2
X_7672__47 _7672__47/A vssd1 vssd1 vccd1 vccd1 _8516_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _8158_/Q _4465_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4981_/A sky130_fd_sc_hd__mux2_1
X_6777__363 _6777__363/A vssd1 vssd1 vccd1 vccd1 _8076_/CLK sky130_fd_sc_hd__inv_2
X_3931_ _3908_/X _8505_/Q _3933_/S vssd1 vssd1 vccd1 vccd1 _3932_/A sky130_fd_sc_hd__mux2_1
X_6738__336 _6742__340/A vssd1 vssd1 vccd1 vccd1 _8046_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3431_ clkbuf_0__3431_/X vssd1 vssd1 vccd1 vccd1 _7058_/A sky130_fd_sc_hd__clkbuf_4
X_6970__431 _6973__434/A vssd1 vssd1 vccd1 vccd1 _8155_/CLK sky130_fd_sc_hd__inv_2
X_3862_ _5345_/A _5345_/B vssd1 vssd1 vccd1 vccd1 _5346_/A sky130_fd_sc_hd__or2_1
X_5601_ _5601_/A vssd1 vssd1 vccd1 vccd1 _7982_/D sky130_fd_sc_hd__clkbuf_1
X_8320_ _8320_/CLK _8320_/D vssd1 vssd1 vccd1 vccd1 _8320_/Q sky130_fd_sc_hd__dfxtp_1
X_5532_ _5383_/X _8031_/Q _5534_/S vssd1 vssd1 vccd1 vccd1 _5533_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7066__506 _7069__509/A vssd1 vssd1 vccd1 vccd1 _8233_/CLK sky130_fd_sc_hd__inv_2
X_8251_ _8251_/CLK _8251_/D vssd1 vssd1 vccd1 vccd1 _8251_/Q sky130_fd_sc_hd__dfxtp_1
X_5463_ _5463_/A vssd1 vssd1 vccd1 vccd1 _8065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4414_ _4394_/X _8270_/Q _4416_/S vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__mux2_1
X_7202_ _8356_/Q _7257_/A _8357_/Q vssd1 vssd1 vccd1 vccd1 _7344_/B sky130_fd_sc_hd__a21o_1
X_5394_ _5367_/X _8096_/Q _5402_/S vssd1 vssd1 vccd1 vccd1 _5395_/A sky130_fd_sc_hd__mux2_1
X_8182_ _8182_/CLK _8182_/D vssd1 vssd1 vccd1 vccd1 _8182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8563__210 vssd1 vssd1 vccd1 vccd1 _8563__210/HI caravel_irq[1] sky130_fd_sc_hd__conb_1
X_4345_ _4345_/A vssd1 vssd1 vccd1 vccd1 _8298_/D sky130_fd_sc_hd__clkbuf_1
X_7394__120 _7394__120/A vssd1 vssd1 vccd1 vccd1 _8377_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4276_ _5500_/B _5464_/B vssd1 vssd1 vccd1 vccd1 _4299_/S sky130_fd_sc_hd__or2_2
X_6015_ _8010_/Q _6019_/B vssd1 vssd1 vccd1 vccd1 _6016_/A sky130_fd_sc_hd__and2_1
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _8526_/CLK _7966_/D vssd1 vssd1 vccd1 vccd1 _7966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7897_ _8531_/CLK _7897_/D vssd1 vssd1 vccd1 vccd1 _7897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6848_ _7754_/A _7521_/B vssd1 vssd1 vccd1 vccd1 _6848_/X sky130_fd_sc_hd__xor2_1
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8518_ _8518_/CLK _8518_/D vssd1 vssd1 vccd1 vccd1 _8518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8449_ _8449_/CLK _8449_/D vssd1 vssd1 vccd1 vccd1 _8449_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3459_ _7096_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3459_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3776_ clkbuf_0__3776_/X vssd1 vssd1 vccd1 vccd1 _7672__47/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_11_wb_clk_i clkbuf_1_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _8531_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4130_ _4929_/A _4622_/A vssd1 vssd1 vccd1 vccd1 _4131_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4061_ _4061_/A vssd1 vssd1 vccd1 vccd1 _8426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7820_ _8355_/CLK _7820_/D vssd1 vssd1 vccd1 vccd1 _7820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7751_ _7522_/A _7743_/X _7750_/X _7737_/X vssd1 vssd1 vccd1 vccd1 _8546_/D sky130_fd_sc_hd__o211a_1
XFILLER_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4963_ _8165_/Q _4471_/X _4969_/S vssd1 vssd1 vccd1 vccd1 _4964_/A sky130_fd_sc_hd__mux2_1
X_3914_ _4567_/A vssd1 vssd1 vccd1 vccd1 _5787_/A sky130_fd_sc_hd__buf_2
X_6702_ _8019_/Q _5965_/A _6706_/S vssd1 vssd1 vccd1 vccd1 _6703_/A sky130_fd_sc_hd__mux2_1
X_7682_ _7682_/A vssd1 vssd1 vccd1 vccd1 _8524_/D sky130_fd_sc_hd__clkbuf_1
X_6597__281 _6600__284/A vssd1 vssd1 vccd1 vccd1 _7959_/CLK sky130_fd_sc_hd__inv_2
X_4894_ _4955_/B _4892_/X _4893_/X vssd1 vssd1 vccd1 vccd1 _4894_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3845_ _8117_/Q vssd1 vssd1 vccd1 vccd1 _3845_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5515_ _5515_/A vssd1 vssd1 vccd1 vccd1 _8039_/D sky130_fd_sc_hd__clkbuf_1
X_8303_ _8303_/CLK _8303_/D vssd1 vssd1 vccd1 vccd1 _8303_/Q sky130_fd_sc_hd__dfxtp_1
X_6495_ _6495_/A vssd1 vssd1 vccd1 vccd1 _7889_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3313_ _6749_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3313_/X sky130_fd_sc_hd__clkbuf_16
X_5446_ _5500_/A _5482_/A vssd1 vssd1 vccd1 vccd1 _5462_/S sky130_fd_sc_hd__nor2_2
X_8234_ _8234_/CLK _8234_/D vssd1 vssd1 vccd1 vccd1 _8234_/Q sky130_fd_sc_hd__dfxtp_1
X_5377_ _5377_/A vssd1 vssd1 vccd1 vccd1 _8101_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3244_ _6527_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3244_/X sky130_fd_sc_hd__clkbuf_16
X_8165_ _8165_/CLK _8165_/D vssd1 vssd1 vccd1 vccd1 _8165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4328_ _4286_/X _8305_/Q _4330_/S vssd1 vssd1 vccd1 vccd1 _4329_/A sky130_fd_sc_hd__mux2_1
X_8096_ _8096_/CLK _8096_/D vssd1 vssd1 vccd1 vccd1 _8096_/Q sky130_fd_sc_hd__dfxtp_1
X_4259_ _8332_/Q _4172_/X _4267_/S vssd1 vssd1 vccd1 vccd1 _4260_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6977__437 _6979__439/A vssd1 vssd1 vccd1 vccd1 _8161_/CLK sky130_fd_sc_hd__inv_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7949_ _7949_/CLK _7949_/D vssd1 vssd1 vccd1 vccd1 _7949_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7297__113 _7297__113/A vssd1 vssd1 vccd1 vccd1 _8342_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5300_ _8221_/Q _5270_/X _5207_/X _8205_/Q _5092_/X vssd1 vssd1 vccd1 vccd1 _5300_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6280_ _8361_/Q _6280_/B vssd1 vssd1 vccd1 vccd1 _6280_/X sky130_fd_sc_hd__and2b_1
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5231_ _8239_/Q _8255_/Q _5231_/S vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__mux2_1
X_5162_ _8516_/Q _8069_/Q _8042_/Q _8500_/Q _5290_/S _5129_/X vssd1 vssd1 vccd1 vccd1
+ _5162_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4113_ _4113_/A vssd1 vssd1 vccd1 vccd1 _8403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5093_ _8212_/Q _8196_/Q _8458_/Q _8228_/Q _5087_/X _5061_/A vssd1 vssd1 vccd1 vccd1
+ _5093_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4044_ _4044_/A vssd1 vssd1 vccd1 vccd1 _8433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7803_ _8531_/CLK _7803_/D vssd1 vssd1 vccd1 vccd1 _7803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6937__410 _6937__410/A vssd1 vssd1 vccd1 vccd1 _8132_/CLK sky130_fd_sc_hd__inv_2
X_5995_ _5995_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5996_/A sky130_fd_sc_hd__and2_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7734_ _5924_/A _7731_/X _7723_/X vssd1 vssd1 vccd1 vccd1 _7734_/X sky130_fd_sc_hd__a21bo_1
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4946_ _4946_/A vssd1 vssd1 vccd1 vccd1 _8173_/D sky130_fd_sc_hd__clkbuf_1
X_4877_ _7975_/Q _8262_/Q _4901_/S vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__mux2_1
X_7596_ _7600_/A _7596_/B vssd1 vssd1 vccd1 vccd1 _8475_/D sky130_fd_sc_hd__nor2_1
X_6616_ _6616_/A vssd1 vssd1 vccd1 vccd1 _7970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3259_ clkbuf_0__3259_/X vssd1 vssd1 vccd1 vccd1 _6604__287/A sky130_fd_sc_hd__clkbuf_4
X_6478_ _6511_/A vssd1 vssd1 vccd1 vccd1 _6487_/S sky130_fd_sc_hd__clkbuf_2
X_5429_ _5444_/S vssd1 vssd1 vccd1 vccd1 _5438_/S sky130_fd_sc_hd__buf_2
X_8217_ _8217_/CLK _8217_/D vssd1 vssd1 vccd1 vccd1 _8217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8148_ _8148_/CLK _8148_/D vssd1 vssd1 vccd1 vccd1 _8148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_1 _7821_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8079_ _8079_/CLK _8079_/D vssd1 vssd1 vccd1 vccd1 _8079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3089_ _6304_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3089_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3475_ clkbuf_0__3475_/X vssd1 vssd1 vccd1 vccd1 _7179__97/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6548__242 _6549__243/A vssd1 vssd1 vccd1 vccd1 _7920_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7416__137 _7416__137/A vssd1 vssd1 vccd1 vccd1 _8394_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4800_ _4790_/X _4793_/X _4694_/X _4799_/X vssd1 vssd1 vccd1 vccd1 _4800_/X sky130_fd_sc_hd__a211o_1
XFILLER_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5780_ _5780_/A vssd1 vssd1 vccd1 vccd1 _7849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4755_/A _4731_/B vssd1 vssd1 vccd1 vccd1 _4731_/X sky130_fd_sc_hd__and2_1
XFILLER_9_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4662_ _4714_/A _4650_/X _4661_/X vssd1 vssd1 vccd1 vccd1 _4662_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6401_ _6331_/X _6399_/X _6400_/X vssd1 vssd1 vccd1 vccd1 _7860_/D sky130_fd_sc_hd__a21o_1
XFILLER_115_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4593_ _4593_/A vssd1 vssd1 vccd1 vccd1 _8202_/D sky130_fd_sc_hd__clkbuf_1
X_7381_ _8368_/Q _7383_/B vssd1 vssd1 vccd1 vccd1 _7381_/X sky130_fd_sc_hd__or2_1
X_6332_ _8551_/Q vssd1 vssd1 vccd1 vccd1 _7247_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6263_ _6263_/A vssd1 vssd1 vccd1 vccd1 _7817_/D sky130_fd_sc_hd__clkbuf_1
X_5214_ _5214_/A vssd1 vssd1 vccd1 vccd1 _5214_/X sky130_fd_sc_hd__clkbuf_2
X_8002_ _8540_/CLK _8002_/D vssd1 vssd1 vccd1 vccd1 _8002_/Q sky130_fd_sc_hd__dfxtp_1
X_6194_ _6239_/A vssd1 vssd1 vccd1 vccd1 _6213_/A sky130_fd_sc_hd__buf_4
X_5145_ _5258_/A vssd1 vssd1 vccd1 vccd1 _5293_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5215_/S vssd1 vssd1 vccd1 vccd1 _5321_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4027_ _4292_/A vssd1 vssd1 vccd1 vccd1 _4027_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5978_ _5978_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _5979_/A sky130_fd_sc_hd__and2_1
XFILLER_13_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3776_ _7670_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3776_/X sky130_fd_sc_hd__clkbuf_16
X_7717_ _7717_/A vssd1 vssd1 vccd1 vccd1 _7717_/X sky130_fd_sc_hd__clkbuf_2
X_4929_ _4929_/A _4945_/B vssd1 vssd1 vccd1 vccd1 _4943_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7579_ _6853_/A _7570_/X _7575_/X _7514_/B vssd1 vssd1 vccd1 vccd1 _7580_/B sky130_fd_sc_hd__o22a_1
XFILLER_109_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_108 _5969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3458_ clkbuf_0__3458_/X vssd1 vssd1 vccd1 vccd1 _7095__530/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_119 _7247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6324__222 _6325__223/A vssd1 vssd1 vccd1 vccd1 _7852_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6771__358 _6772__359/A vssd1 vssd1 vccd1 vccd1 _8071_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6177__185 _6177__185/A vssd1 vssd1 vccd1 vccd1 _7772_/CLK sky130_fd_sc_hd__inv_2
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5901_ _7631_/A _5910_/B vssd1 vssd1 vccd1 vccd1 _5902_/A sky130_fd_sc_hd__or2_1
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5832_ _5832_/A vssd1 vssd1 vccd1 vccd1 _7826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5763_ _7904_/Q _5569_/A _5767_/S vssd1 vssd1 vccd1 vccd1 _5764_/A sky130_fd_sc_hd__mux2_1
X_8551_ _8551_/CLK _8551_/D vssd1 vssd1 vccd1 vccd1 _8551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4714_ _4714_/A vssd1 vssd1 vccd1 vccd1 _4953_/B sky130_fd_sc_hd__clkbuf_2
X_7502_ _7502_/A input1/X vssd1 vssd1 vccd1 vccd1 _7503_/C sky130_fd_sc_hd__nor2_1
X_5694_ _5694_/A vssd1 vssd1 vccd1 vccd1 _7935_/D sky130_fd_sc_hd__clkbuf_1
X_8482_ _8486_/CLK _8482_/D vssd1 vssd1 vccd1 vccd1 _8482_/Q sky130_fd_sc_hd__dfxtp_1
X_7433_ _7439_/A vssd1 vssd1 vccd1 vccd1 _7433_/X sky130_fd_sc_hd__buf_1
X_4645_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4646_/A sky130_fd_sc_hd__buf_2
X_4576_ _4576_/A vssd1 vssd1 vccd1 vccd1 _8209_/D sky130_fd_sc_hd__clkbuf_1
X_7364_ _7364_/A vssd1 vssd1 vccd1 vccd1 _7679_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3027_ clkbuf_0__3027_/X vssd1 vssd1 vccd1 vccd1 _6185__191/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6246_ _8021_/Q _6188_/X _6202_/A _6213_/A _7810_/Q vssd1 vssd1 vccd1 vccd1 _7810_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5128_ _5169_/A _5128_/B vssd1 vssd1 vccd1 vccd1 _5128_/X sky130_fd_sc_hd__and2_1
Xclkbuf_1_0_0__3312_ clkbuf_0__3312_/X vssd1 vssd1 vccd1 vccd1 _6748__345/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5059_ _5181_/A vssd1 vssd1 vccd1 vccd1 _5129_/A sky130_fd_sc_hd__buf_2
XFILLER_38_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8580__227 vssd1 vssd1 vccd1 vccd1 _8580__227/HI core1Index[7] sky130_fd_sc_hd__conb_1
XFILLER_88_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6591__276 _6595__280/A vssd1 vssd1 vccd1 vccd1 _7954_/CLK sky130_fd_sc_hd__inv_2
X_4430_ _4430_/A vssd1 vssd1 vccd1 vccd1 _8266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6100_ _7869_/Q input9/X _6111_/S vssd1 vssd1 vccd1 vccd1 _6100_/X sky130_fd_sc_hd__mux2_1
X_4361_ _4361_/A vssd1 vssd1 vccd1 vccd1 _8291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4292_ _4292_/A vssd1 vssd1 vccd1 vccd1 _4292_/X sky130_fd_sc_hd__clkbuf_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _6031_/A vssd1 vssd1 vccd1 vccd1 _6031_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7982_ _7982_/CLK _7982_/D vssd1 vssd1 vccd1 vccd1 _7982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3645_ clkbuf_0__3645_/X vssd1 vssd1 vccd1 vccd1 _7439_/A sky130_fd_sc_hd__clkbuf_4
X_6864_ _8477_/Q vssd1 vssd1 vccd1 vccd1 _6865_/B sky130_fd_sc_hd__inv_2
X_5815_ _3972_/X _7833_/Q _5815_/S vssd1 vssd1 vccd1 vccd1 _5816_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6795_ _6795_/A vssd1 vssd1 vccd1 vccd1 _6824_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5746_ _5746_/A vssd1 vssd1 vccd1 vccd1 _7912_/D sky130_fd_sc_hd__clkbuf_1
X_8534_ _8548_/CLK _8534_/D vssd1 vssd1 vccd1 vccd1 _8534_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5677_ _5575_/X _7942_/Q _5677_/S vssd1 vssd1 vccd1 vccd1 _5678_/A sky130_fd_sc_hd__mux2_1
X_8465_ _8487_/CLK _8465_/D vssd1 vssd1 vccd1 vccd1 _8465_/Q sky130_fd_sc_hd__dfxtp_2
X_4628_ _8187_/Q _6605_/B vssd1 vssd1 vccd1 vccd1 _4764_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8396_ _8396_/CLK _8396_/D vssd1 vssd1 vccd1 vccd1 _8396_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3475_ _7177_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3475_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4559_ _4435_/X _8216_/Q _4559_/S vssd1 vssd1 vccd1 vccd1 _4560_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7347_ _8358_/Q _7334_/A _7310_/A _7201_/B vssd1 vssd1 vccd1 vccd1 _7348_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7278_ _8537_/Q _7344_/A _7344_/B vssd1 vssd1 vccd1 vccd1 _7278_/X sky130_fd_sc_hd__and3_1
XFILLER_106_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6229_ _6239_/A vssd1 vssd1 vccd1 vccd1 _6229_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7291__108 _7293__110/A vssd1 vssd1 vccd1 vccd1 _8337_/CLK sky130_fd_sc_hd__inv_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3088_ clkbuf_0__3088_/X vssd1 vssd1 vccd1 vccd1 _6303__205/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7024__473 _7026__475/A vssd1 vssd1 vccd1 vccd1 _8200_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3930_ _3930_/A vssd1 vssd1 vccd1 vccd1 _8506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3430_ clkbuf_0__3430_/X vssd1 vssd1 vccd1 vccd1 _6960__425/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _8133_/Q _5335_/A vssd1 vssd1 vccd1 vccd1 _5345_/B sky130_fd_sc_hd__nand2_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5600_ _7982_/Q _5599_/X _5600_/S vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__mux2_1
X_6931__405 _6931__405/A vssd1 vssd1 vccd1 vccd1 _8127_/CLK sky130_fd_sc_hd__inv_2
X_5531_ _5531_/A vssd1 vssd1 vccd1 vccd1 _8032_/D sky130_fd_sc_hd__clkbuf_1
X_8250_ _8250_/CLK _8250_/D vssd1 vssd1 vccd1 vccd1 _8250_/Q sky130_fd_sc_hd__dfxtp_1
X_5462_ _8065_/Q _4196_/X _5462_/S vssd1 vssd1 vccd1 vccd1 _5463_/A sky130_fd_sc_hd__mux2_1
X_7201_ _7201_/A _7201_/B vssd1 vssd1 vccd1 vccd1 _7284_/B sky130_fd_sc_hd__xor2_1
X_4413_ _4413_/A vssd1 vssd1 vccd1 vccd1 _8271_/D sky130_fd_sc_hd__clkbuf_1
X_8181_ _8181_/CLK _8181_/D vssd1 vssd1 vccd1 vccd1 _8181_/Q sky130_fd_sc_hd__dfxtp_1
X_5393_ _5393_/A vssd1 vssd1 vccd1 vccd1 _8097_/D sky130_fd_sc_hd__clkbuf_1
X_4344_ _4283_/X _8298_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4345_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6014_ _6014_/A vssd1 vssd1 vccd1 vccd1 _6014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4275_ _4275_/A vssd1 vssd1 vccd1 vccd1 _4275_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7965_ _7965_/CLK _7965_/D vssd1 vssd1 vccd1 vccd1 _7965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7896_ _8520_/CLK _7896_/D vssd1 vssd1 vccd1 vccd1 _7896_/Q sky130_fd_sc_hd__dfxtp_1
X_6847_ _6847_/A _7556_/A vssd1 vssd1 vccd1 vccd1 _7521_/B sky130_fd_sc_hd__xnor2_2
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8517_ _8517_/CLK _8517_/D vssd1 vssd1 vccd1 vccd1 _8517_/Q sky130_fd_sc_hd__dfxtp_1
X_5729_ _7919_/Q _5596_/X _5731_/S vssd1 vssd1 vccd1 vccd1 _5730_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8448_ _8448_/CLK _8448_/D vssd1 vssd1 vccd1 vccd1 _8448_/Q sky130_fd_sc_hd__dfxtp_1
X_8379_ _8379_/CLK _8379_/D vssd1 vssd1 vccd1 vccd1 _8379_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3458_ _7090_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3458_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3775_ clkbuf_0__3775_/X vssd1 vssd1 vccd1 vccd1 _7666__42/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6542__237 _6544__239/A vssd1 vssd1 vccd1 vccd1 _7915_/CLK sky130_fd_sc_hd__inv_2
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8586__233 vssd1 vssd1 vccd1 vccd1 _8586__233/HI manufacturerID[5] sky130_fd_sc_hd__conb_1
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6744__341 _6746__343/A vssd1 vssd1 vccd1 vccd1 _8051_/CLK sky130_fd_sc_hd__inv_2
X_4060_ _4005_/X _8426_/Q _4068_/S vssd1 vssd1 vccd1 vccd1 _4061_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7072__511 _7073__512/A vssd1 vssd1 vccd1 vccd1 _8238_/CLK sky130_fd_sc_hd__inv_2
X_7750_ _7642_/A _7702_/A _7744_/X vssd1 vssd1 vccd1 vccd1 _7750_/X sky130_fd_sc_hd__a21bo_1
X_4962_ _4962_/A vssd1 vssd1 vccd1 vccd1 _8166_/D sky130_fd_sc_hd__clkbuf_1
X_3913_ _3913_/A vssd1 vssd1 vccd1 vccd1 _8512_/D sky130_fd_sc_hd__clkbuf_1
X_4893_ _8335_/Q _4811_/X _8143_/Q _4781_/X _4739_/S vssd1 vssd1 vccd1 vccd1 _4893_/X
+ sky130_fd_sc_hd__o221a_1
X_6701_ _6701_/A vssd1 vssd1 vccd1 vccd1 _8018_/D sky130_fd_sc_hd__clkbuf_1
X_7681_ _8124_/Q _7737_/A vssd1 vssd1 vccd1 vccd1 _7682_/A sky130_fd_sc_hd__and2_1
X_6632_ _6632_/A vssd1 vssd1 vccd1 vccd1 _6632_/X sky130_fd_sc_hd__buf_1
XFILLER_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3844_ _5034_/C _5034_/D _5034_/B vssd1 vssd1 vccd1 vccd1 _3860_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5514_ _8039_/Q _4295_/A _5516_/S vssd1 vssd1 vccd1 vccd1 _5515_/A sky130_fd_sc_hd__mux2_1
X_8302_ _8302_/CLK _8302_/D vssd1 vssd1 vccd1 vccd1 _8302_/Q sky130_fd_sc_hd__dfxtp_1
X_6494_ _6002_/A _7889_/Q _6498_/S vssd1 vssd1 vccd1 vccd1 _6495_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3312_ _6743_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3312_/X sky130_fd_sc_hd__clkbuf_16
X_5445_ _5445_/A vssd1 vssd1 vccd1 vccd1 _8073_/D sky130_fd_sc_hd__clkbuf_1
X_8233_ _8233_/CLK _8233_/D vssd1 vssd1 vccd1 vccd1 _8233_/Q sky130_fd_sc_hd__dfxtp_1
X_8164_ _8164_/CLK _8164_/D vssd1 vssd1 vccd1 vccd1 _8164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5376_ _5375_/X _8101_/Q _5376_/S vssd1 vssd1 vccd1 vccd1 _5377_/A sky130_fd_sc_hd__mux2_1
X_4327_ _4327_/A vssd1 vssd1 vccd1 vccd1 _8306_/D sky130_fd_sc_hd__clkbuf_1
X_8095_ _8095_/CLK _8095_/D vssd1 vssd1 vccd1 vccd1 _8095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4258_ _4273_/S vssd1 vssd1 vccd1 vccd1 _4267_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7046_ _7052_/A vssd1 vssd1 vccd1 vccd1 _7046_/X sky130_fd_sc_hd__buf_1
XFILLER_59_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4189_ _4189_/A vssd1 vssd1 vccd1 vccd1 _8390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7948_ _7948_/CLK _7948_/D vssd1 vssd1 vccd1 vccd1 _7948_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7879_ _8345_/CLK _7879_/D vssd1 vssd1 vccd1 vccd1 _7879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7175__94 _7176__95/A vssd1 vssd1 vccd1 vccd1 _8321_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5230_ _5230_/A vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5161_ _7842_/Q _8050_/Q _8329_/Q _8077_/Q _5273_/S _5068_/X vssd1 vssd1 vccd1 vccd1
+ _5161_/X sky130_fd_sc_hd__mux4_1
X_4112_ _4035_/X _8403_/Q _4112_/S vssd1 vssd1 vccd1 vccd1 _4113_/A sky130_fd_sc_hd__mux2_1
X_5092_ _5092_/A vssd1 vssd1 vccd1 vccd1 _5092_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8560__258 vssd1 vssd1 vccd1 vccd1 partID[14] _8560__258/LO sky130_fd_sc_hd__conb_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4043_ _4011_/X _8433_/Q _4049_/S vssd1 vssd1 vccd1 vccd1 _4044_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5994_ _5994_/A vssd1 vssd1 vccd1 vccd1 _5994_/X sky130_fd_sc_hd__clkbuf_1
X_7802_ _8531_/CLK _7802_/D vssd1 vssd1 vccd1 vccd1 _7802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7733_ _8540_/Q _7717_/X _7732_/X _7719_/X vssd1 vssd1 vccd1 vccd1 _8540_/D sky130_fd_sc_hd__o211a_1
XFILLER_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4945_ _7008_/C _4945_/B _4945_/C vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__and3_1
X_7037__483 _7038__484/A vssd1 vssd1 vccd1 vccd1 _8210_/CLK sky130_fd_sc_hd__inv_2
X_4876_ _4876_/A vssd1 vssd1 vccd1 vccd1 _4901_/S sky130_fd_sc_hd__buf_2
X_7664_ _7664_/A vssd1 vssd1 vccd1 vccd1 _7664_/X sky130_fd_sc_hd__buf_1
XFILLER_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7595_ _6812_/A _7588_/X _7547_/X _6814_/B vssd1 vssd1 vccd1 vccd1 _7596_/B sky130_fd_sc_hd__o22a_1
X_6615_ _8183_/Q _6621_/B vssd1 vssd1 vccd1 vccd1 _6616_/A sky130_fd_sc_hd__and2_1
X_6546_ _6552_/A vssd1 vssd1 vccd1 vccd1 _6546_/X sky130_fd_sc_hd__buf_1
XFILLER_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3258_ clkbuf_0__3258_/X vssd1 vssd1 vccd1 vccd1 _6601__285/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6477_ _6477_/A vssd1 vssd1 vccd1 vccd1 _7881_/D sky130_fd_sc_hd__clkbuf_1
X_5428_ _5428_/A _5787_/B vssd1 vssd1 vccd1 vccd1 _5444_/S sky130_fd_sc_hd__or2_2
X_8216_ _8216_/CLK _8216_/D vssd1 vssd1 vccd1 vccd1 _8216_/Q sky130_fd_sc_hd__dfxtp_1
X_6983__442 _6983__442/A vssd1 vssd1 vccd1 vccd1 _8166_/CLK sky130_fd_sc_hd__inv_2
X_7475__10 _7474__9/A vssd1 vssd1 vccd1 vccd1 _8442_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8147_ _8147_/CLK _8147_/D vssd1 vssd1 vccd1 vccd1 _8147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5359_ _5281_/S _5348_/X _5358_/Y vssd1 vssd1 vccd1 vccd1 _8114_/D sky130_fd_sc_hd__a21oi_1
X_8078_ _8078_/CLK _8078_/D vssd1 vssd1 vccd1 vccd1 _8078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7079__517 _7079__517/A vssd1 vssd1 vccd1 vccd1 _8244_/CLK sky130_fd_sc_hd__inv_2
XINSDIODE2_2 _7821_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3088_ _6298_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3088_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3474_ clkbuf_0__3474_/X vssd1 vssd1 vccd1 vccd1 _7176__95/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7148__72 _7149__73/A vssd1 vssd1 vccd1 vccd1 _8299_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4730_ _7827_/Q _7947_/Q _7963_/Q _7931_/Q _4729_/X _4716_/A vssd1 vssd1 vccd1 vccd1
+ _4731_/B sky130_fd_sc_hd__mux4_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4661_ _4654_/X _4657_/X _4951_/B vssd1 vssd1 vccd1 vccd1 _4661_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6400_ _7860_/Q _6328_/A _6233_/X vssd1 vssd1 vccd1 vccd1 _6400_/X sky130_fd_sc_hd__a21o_1
X_7380_ _8130_/Q _7364_/A _7366_/A _7379_/X _7371_/X vssd1 vssd1 vccd1 vccd1 _8367_/D
+ sky130_fd_sc_hd__o311a_1
X_4592_ _4428_/X _8202_/Q _4596_/S vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__mux2_1
X_6331_ _6331_/A vssd1 vssd1 vccd1 vccd1 _6331_/X sky130_fd_sc_hd__clkbuf_2
X_6262_ _7644_/A _7817_/Q _6264_/S vssd1 vssd1 vccd1 vccd1 _6263_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5213_ _5193_/X _5211_/X _5212_/X vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__o21a_1
X_8001_ _8540_/CLK _8001_/D vssd1 vssd1 vccd1 vccd1 _8001_/Q sky130_fd_sc_hd__dfxtp_1
X_6193_ _6466_/A _6272_/B vssd1 vssd1 vccd1 vccd1 _6239_/A sky130_fd_sc_hd__or2_4
X_5144_ _5055_/A _5141_/X _5143_/X vssd1 vssd1 vccd1 vccd1 _5144_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5075_ _5182_/B vssd1 vssd1 vccd1 vccd1 _5215_/S sky130_fd_sc_hd__buf_4
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4026_ _8490_/Q vssd1 vssd1 vccd1 vccd1 _4292_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5977_ _6010_/A vssd1 vssd1 vccd1 vccd1 _5986_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6757__351 _6766__354/A vssd1 vssd1 vccd1 vccd1 _8061_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3775_ _7664_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3775_/X sky130_fd_sc_hd__clkbuf_16
X_7716_ _7728_/C vssd1 vssd1 vccd1 vccd1 _7717_/A sky130_fd_sc_hd__clkbuf_2
X_4928_ _4944_/A _4944_/B vssd1 vssd1 vccd1 vccd1 _4945_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7647_ _7647_/A vssd1 vssd1 vccd1 vccd1 _8495_/D sky130_fd_sc_hd__clkbuf_1
X_4859_ _7991_/Q _8099_/Q _4873_/S vssd1 vssd1 vccd1 vccd1 _4859_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7578_ _7585_/A _7578_/B vssd1 vssd1 vccd1 vccd1 _8468_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6868__368 _6870__370/A vssd1 vssd1 vccd1 vccd1 _8082_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3457_ clkbuf_0__3457_/X vssd1 vssd1 vccd1 vccd1 _7114_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_109 _5969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7422__142 _7422__142/A vssd1 vssd1 vccd1 vccd1 _8399_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5900_ _5969_/B vssd1 vssd1 vccd1 vccd1 _5910_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5831_ _7826_/Q _5399_/A _5833_/S vssd1 vssd1 vccd1 vccd1 _5832_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5762_ _5762_/A vssd1 vssd1 vccd1 vccd1 _7905_/D sky130_fd_sc_hd__clkbuf_1
X_8550_ _8550_/CLK _8550_/D vssd1 vssd1 vccd1 vccd1 _8550_/Q sky130_fd_sc_hd__dfxtp_4
X_6637__300 _6637__300/A vssd1 vssd1 vccd1 vccd1 _7986_/CLK sky130_fd_sc_hd__inv_2
X_7501_ _8460_/Q _7550_/C vssd1 vssd1 vccd1 vccd1 _7541_/A sky130_fd_sc_hd__nand2_1
X_4713_ _4713_/A vssd1 vssd1 vccd1 vccd1 _4713_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_6_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _8527_/CLK sky130_fd_sc_hd__clkbuf_16
X_5693_ _7935_/Q _5596_/X _5695_/S vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__mux2_1
X_8481_ _8486_/CLK _8481_/D vssd1 vssd1 vccd1 vccd1 _8481_/Q sky130_fd_sc_hd__dfxtp_1
X_7432_ _7432_/A vssd1 vssd1 vccd1 vccd1 _7432_/X sky130_fd_sc_hd__buf_1
X_4644_ _4766_/B vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4575_ _3969_/X _8209_/Q _4577_/S vssd1 vssd1 vccd1 vccd1 _4576_/A sky130_fd_sc_hd__mux2_1
X_7363_ _7363_/A vssd1 vssd1 vccd1 vccd1 _7364_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7294_ _7389_/A vssd1 vssd1 vccd1 vccd1 _7294_/X sky130_fd_sc_hd__buf_1
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3026_ clkbuf_0__3026_/X vssd1 vssd1 vccd1 vccd1 _6183__190/A sky130_fd_sc_hd__clkbuf_4
X_7142__67 _7142__67/A vssd1 vssd1 vccd1 vccd1 _8294_/CLK sky130_fd_sc_hd__inv_2
X_6245_ _8020_/Q _6188_/X _6202_/A _6213_/A _7809_/Q vssd1 vssd1 vccd1 vccd1 _7809_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_103_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6644__304 _6645__305/A vssd1 vssd1 vccd1 vccd1 _7990_/CLK sky130_fd_sc_hd__inv_2
X_5127_ _8510_/Q _8259_/Q _8243_/Q _8283_/Q _5087_/X _5061_/A vssd1 vssd1 vccd1 vccd1
+ _5128_/B sky130_fd_sc_hd__mux4_2
Xclkbuf_1_0_0__3311_ clkbuf_0__3311_/X vssd1 vssd1 vccd1 vccd1 _6740__338/A sky130_fd_sc_hd__clkbuf_4
X_5058_ _5231_/S vssd1 vssd1 vccd1 vccd1 _5284_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4009_ _4009_/A vssd1 vssd1 vccd1 vccd1 _8442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6996__452 _6999__455/A vssd1 vssd1 vccd1 vccd1 _8177_/CLK sky130_fd_sc_hd__inv_2
X_6287__192 _6290__195/A vssd1 vssd1 vccd1 vccd1 _7822_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6183__190 _6183__190/A vssd1 vssd1 vccd1 vccd1 _7777_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4360_ _4280_/X _8291_/Q _4366_/S vssd1 vssd1 vccd1 vccd1 _4361_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4291_ _4291_/A vssd1 vssd1 vccd1 vccd1 _8320_/D sky130_fd_sc_hd__clkbuf_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6708__312 _6711__315/A vssd1 vssd1 vccd1 vccd1 _8022_/CLK sky130_fd_sc_hd__inv_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _8017_/Q _6030_/B vssd1 vssd1 vccd1 vccd1 _6031_/A sky130_fd_sc_hd__and2_4
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7981_ _7981_/CLK _7981_/D vssd1 vssd1 vccd1 vccd1 _7981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6932_ _6932_/A vssd1 vssd1 vccd1 vccd1 _6932_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__3644_ clkbuf_0__3644_/X vssd1 vssd1 vccd1 vccd1 _7431__150/A sky130_fd_sc_hd__clkbuf_4
X_6863_ _8478_/Q vssd1 vssd1 vccd1 vccd1 _6865_/A sky130_fd_sc_hd__inv_2
X_5814_ _5814_/A vssd1 vssd1 vccd1 vccd1 _7834_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3575_ clkbuf_0__3575_/X vssd1 vssd1 vccd1 vccd1 _7388__115/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6794_ _6818_/A vssd1 vssd1 vccd1 vccd1 _6830_/A sky130_fd_sc_hd__buf_2
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7429__148 _7429__148/A vssd1 vssd1 vccd1 vccd1 _8405_/CLK sky130_fd_sc_hd__inv_2
X_5745_ _7912_/Q _5569_/A _5749_/S vssd1 vssd1 vccd1 vccd1 _5746_/A sky130_fd_sc_hd__mux2_1
X_8533_ _8548_/CLK _8533_/D vssd1 vssd1 vccd1 vccd1 _8533_/Q sky130_fd_sc_hd__dfxtp_1
X_5676_ _5676_/A vssd1 vssd1 vccd1 vccd1 _7943_/D sky130_fd_sc_hd__clkbuf_1
X_8464_ _8487_/CLK _8464_/D vssd1 vssd1 vccd1 vccd1 _8464_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3474_ _7171_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3474_/X sky130_fd_sc_hd__clkbuf_16
X_4627_ _4622_/X _4627_/B _4627_/C _4627_/D vssd1 vssd1 vccd1 vccd1 _6605_/B sky130_fd_sc_hd__and4b_2
X_8395_ _8395_/CLK _8395_/D vssd1 vssd1 vccd1 vccd1 _8395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4558_ _4558_/A vssd1 vssd1 vccd1 vccd1 _8217_/D sky130_fd_sc_hd__clkbuf_1
X_7346_ _7348_/A _7346_/B vssd1 vssd1 vccd1 vccd1 _8357_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4489_ _4489_/A vssd1 vssd1 vccd1 vccd1 _8245_/D sky130_fd_sc_hd__clkbuf_1
X_7277_ _7275_/X _7277_/B _7277_/C _7277_/D vssd1 vssd1 vccd1 vccd1 _7284_/C sky130_fd_sc_hd__and4b_1
X_6228_ _6225_/X _8009_/Q _6227_/X _6221_/X _7798_/Q vssd1 vssd1 vccd1 vccd1 _7798_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_106_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6466_/A vssd1 vssd1 vccd1 vccd1 _7689_/A sky130_fd_sc_hd__inv_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3087_ clkbuf_0__3087_/X vssd1 vssd1 vccd1 vccd1 _6310_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7657__35 _7657__35/A vssd1 vssd1 vccd1 vccd1 _8504_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3860_ _3860_/A _3860_/B _3860_/C _3860_/D vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__or4_1
XFILLER_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ _5379_/X _8032_/Q _5534_/S vssd1 vssd1 vccd1 vccd1 _5531_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7031__478 _7033__480/A vssd1 vssd1 vccd1 vccd1 _8205_/CLK sky130_fd_sc_hd__inv_2
X_5461_ _5461_/A vssd1 vssd1 vccd1 vccd1 _8066_/D sky130_fd_sc_hd__clkbuf_1
X_4412_ _4391_/X _8271_/Q _4416_/S vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7200_ _8358_/Q _7344_/A vssd1 vssd1 vccd1 vccd1 _7201_/B sky130_fd_sc_hd__xor2_1
X_8180_ _8180_/CLK _8180_/D vssd1 vssd1 vccd1 vccd1 _8180_/Q sky130_fd_sc_hd__dfxtp_1
X_5392_ _5361_/X _8097_/Q _5402_/S vssd1 vssd1 vccd1 vccd1 _5393_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4343_ _4343_/A vssd1 vssd1 vccd1 vccd1 _8299_/D sky130_fd_sc_hd__clkbuf_1
X_4274_ _4274_/A vssd1 vssd1 vccd1 vccd1 _8325_/D sky130_fd_sc_hd__clkbuf_1
X_6013_ _8009_/Q _6019_/B vssd1 vssd1 vccd1 vccd1 _6014_/A sky130_fd_sc_hd__and2_1
XFILLER_113_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7435__152 _7436__153/A vssd1 vssd1 vccd1 vccd1 _8409_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7964_ _7964_/CLK _7964_/D vssd1 vssd1 vccd1 vccd1 _7964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7895_ _8520_/CLK _7895_/D vssd1 vssd1 vccd1 vccd1 _7895_/Q sky130_fd_sc_hd__dfxtp_1
X_6846_ _8464_/Q vssd1 vssd1 vccd1 vccd1 _6847_/A sky130_fd_sc_hd__inv_2
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _3989_/A vssd1 vssd1 vccd1 vccd1 _8450_/D sky130_fd_sc_hd__clkbuf_1
X_8516_ _8516_/CLK _8516_/D vssd1 vssd1 vccd1 vccd1 _8516_/Q sky130_fd_sc_hd__dfxtp_1
X_5728_ _5728_/A vssd1 vssd1 vccd1 vccd1 _7920_/D sky130_fd_sc_hd__clkbuf_1
X_8447_ _8447_/CLK _8447_/D vssd1 vssd1 vccd1 vccd1 _8447_/Q sky130_fd_sc_hd__dfxtp_1
X_5659_ _7950_/Q _5599_/X _5659_/S vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__mux2_1
X_8378_ _8378_/CLK _8378_/D vssd1 vssd1 vccd1 vccd1 _8378_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__3457_ _7089_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3457_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_117_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3774_ clkbuf_0__3774_/X vssd1 vssd1 vccd1 vccd1 _7663__40/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7329_ _7329_/A _7329_/B vssd1 vssd1 vccd1 vccd1 _7329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_wb_clk_i _6163_/A vssd1 vssd1 vccd1 vccd1 _8540_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4961_ _8166_/Q _4465_/X _4969_/S vssd1 vssd1 vccd1 vccd1 _4962_/A sky130_fd_sc_hd__mux2_1
X_3912_ _3911_/X _8512_/Q _3912_/S vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__mux2_1
X_4892_ _7990_/Q _8098_/Q _4909_/S vssd1 vssd1 vccd1 vccd1 _4892_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6700_ _8018_/Q _5963_/A _6700_/S vssd1 vssd1 vccd1 vccd1 _6701_/A sky130_fd_sc_hd__mux2_1
X_7680_ _7680_/A _7680_/B vssd1 vssd1 vccd1 vccd1 _8523_/D sky130_fd_sc_hd__nor2_1
X_3843_ _8120_/Q _8115_/Q vssd1 vssd1 vccd1 vccd1 _5034_/B sky130_fd_sc_hd__xnor2_1
X_7474__9 _7474__9/A vssd1 vssd1 vccd1 vccd1 _8441_/CLK sky130_fd_sc_hd__inv_2
X_8301_ _8301_/CLK _8301_/D vssd1 vssd1 vccd1 vccd1 _8301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3274_ clkbuf_0__3274_/X vssd1 vssd1 vccd1 vccd1 _6651__310/A sky130_fd_sc_hd__clkbuf_4
X_5513_ _5513_/A vssd1 vssd1 vccd1 vccd1 _8040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6493_ _6493_/A vssd1 vssd1 vccd1 vccd1 _7888_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3311_ _6737_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3311_/X sky130_fd_sc_hd__clkbuf_16
X_5444_ _3981_/X _8073_/Q _5444_/S vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__mux2_1
X_8232_ _8232_/CLK _8232_/D vssd1 vssd1 vccd1 vccd1 _8232_/Q sky130_fd_sc_hd__dfxtp_1
X_8163_ _8163_/CLK _8163_/D vssd1 vssd1 vccd1 vccd1 _8163_/Q sky130_fd_sc_hd__dfxtp_1
X_7114_ _7114_/A vssd1 vssd1 vccd1 vccd1 _7114_/X sky130_fd_sc_hd__buf_1
X_5375_ _5566_/A vssd1 vssd1 vccd1 vccd1 _5375_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4326_ _4283_/X _8306_/Q _4330_/S vssd1 vssd1 vccd1 vccd1 _4327_/A sky130_fd_sc_hd__mux2_1
X_8094_ _8094_/CLK _8094_/D vssd1 vssd1 vccd1 vccd1 _8094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4257_ _5500_/B _5787_/B vssd1 vssd1 vccd1 vccd1 _4273_/S sky130_fd_sc_hd__nor2_2
XFILLER_101_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4188_ _8390_/Q _4187_/X _4188_/S vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7947_ _7947_/CLK _7947_/D vssd1 vssd1 vccd1 vccd1 _7947_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _8345_/CLK _7878_/D vssd1 vssd1 vccd1 vccd1 _7878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6829_ _6822_/Y _6823_/X _6827_/Y _6828_/X vssd1 vssd1 vccd1 vccd1 _6855_/B sky130_fd_sc_hd__o211a_1
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5160_ _5055_/X _5157_/X _5159_/X vssd1 vssd1 vccd1 vccd1 _5160_/X sky130_fd_sc_hd__a21o_1
X_4111_ _4111_/A vssd1 vssd1 vccd1 vccd1 _8404_/D sky130_fd_sc_hd__clkbuf_1
X_5091_ _5091_/A vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__clkbuf_2
X_4042_ _4042_/A vssd1 vssd1 vccd1 vccd1 _8434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5993_ _5993_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5994_/A sky130_fd_sc_hd__and2_1
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7801_ _8531_/CLK _7801_/D vssd1 vssd1 vccd1 vccd1 _7801_/Q sky130_fd_sc_hd__dfxtp_1
X_7732_ _5926_/A _7731_/X _7723_/X vssd1 vssd1 vccd1 vccd1 _7732_/X sky130_fd_sc_hd__a21bo_1
X_4944_ _4944_/A _4944_/B vssd1 vssd1 vccd1 vccd1 _4945_/C sky130_fd_sc_hd__or2_1
X_4875_ _4770_/X _4873_/X _4874_/X vssd1 vssd1 vccd1 vccd1 _4875_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7594_ _7600_/A _7594_/B vssd1 vssd1 vccd1 vccd1 _8474_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6614_ _6614_/A vssd1 vssd1 vccd1 vccd1 _7969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3257_ clkbuf_0__3257_/X vssd1 vssd1 vccd1 vccd1 _6594__279/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8215_ _8215_/CLK _8215_/D vssd1 vssd1 vccd1 vccd1 _8215_/Q sky130_fd_sc_hd__dfxtp_1
X_6476_ _5984_/A _7881_/Q _6476_/S vssd1 vssd1 vccd1 vccd1 _6477_/A sky130_fd_sc_hd__mux2_1
X_5427_ _5427_/A vssd1 vssd1 vccd1 vccd1 _8082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8146_ _8146_/CLK _8146_/D vssd1 vssd1 vccd1 vccd1 _8146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5358_ _5281_/S _5356_/A _5343_/A vssd1 vssd1 vccd1 vccd1 _5358_/Y sky130_fd_sc_hd__o21ai_1
X_8077_ _8077_/CLK _8077_/D vssd1 vssd1 vccd1 vccd1 _8077_/Q sky130_fd_sc_hd__dfxtp_1
X_4309_ _4309_/A vssd1 vssd1 vccd1 vccd1 _8314_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_3 _7821_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5289_ _5230_/X _5287_/X _5288_/X vssd1 vssd1 vccd1 vccd1 _5293_/B sky130_fd_sc_hd__o21ai_1
XFILLER_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7028_ _7040_/A vssd1 vssd1 vccd1 vccd1 _7028_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3087_ _6297_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3087_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__3473_ clkbuf_0__3473_/X vssd1 vssd1 vccd1 vccd1 _7169__89/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4694_/A vssd1 vssd1 vccd1 vccd1 _4951_/B sky130_fd_sc_hd__buf_2
X_6555__248 _6557__250/A vssd1 vssd1 vccd1 vccd1 _7926_/CLK sky130_fd_sc_hd__inv_2
X_6330_ _7742_/B vssd1 vssd1 vccd1 vccd1 _6331_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4591_ _4591_/A vssd1 vssd1 vccd1 vccd1 _8203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7154__76 _7156__78/A vssd1 vssd1 vccd1 vccd1 _8303_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6261_ _6261_/A vssd1 vssd1 vccd1 vccd1 _7816_/D sky130_fd_sc_hd__clkbuf_1
X_5212_ _8414_/Q _5196_/X _5207_/A _8406_/Q _5167_/S vssd1 vssd1 vccd1 vccd1 _5212_/X
+ sky130_fd_sc_hd__o221a_1
X_6192_ _7820_/Q _7819_/Q vssd1 vssd1 vccd1 vccd1 _6272_/B sky130_fd_sc_hd__or2b_4
X_8000_ _8540_/CLK _8000_/D vssd1 vssd1 vccd1 vccd1 _8000_/Q sky130_fd_sc_hd__dfxtp_1
X_5143_ _5079_/X _5142_/X _5131_/X vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _5055_/X _5062_/X _5073_/X vssd1 vssd1 vccd1 vccd1 _5074_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4025_ _4025_/A vssd1 vssd1 vccd1 vccd1 _8438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5976_ _5976_/A vssd1 vssd1 vccd1 vccd1 _5976_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3774_ _7658_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3774_/X sky130_fd_sc_hd__clkbuf_16
X_7715_ _8063_/Q _7747_/B vssd1 vssd1 vccd1 vccd1 _7728_/C sky130_fd_sc_hd__and2_1
X_4927_ _8176_/Q vssd1 vssd1 vccd1 vccd1 _5014_/B sky130_fd_sc_hd__clkbuf_4
X_4858_ _4438_/X _4629_/X _4856_/X _4857_/X vssd1 vssd1 vccd1 vccd1 _8181_/D sky130_fd_sc_hd__o211a_1
X_7646_ _7646_/A _7646_/B _7646_/C vssd1 vssd1 vccd1 vccd1 _7647_/A sky130_fd_sc_hd__and3_1
X_7085__522 _7087__524/A vssd1 vssd1 vccd1 vccd1 _8249_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3309_ clkbuf_0__3309_/X vssd1 vssd1 vccd1 vccd1 _6727__327/A sky130_fd_sc_hd__clkbuf_4
X_4789_ _8248_/Q _4781_/X _4782_/X _4788_/X vssd1 vssd1 vccd1 vccd1 _4789_/X sky130_fd_sc_hd__o211a_1
X_7577_ _7574_/Y _7570_/X _7575_/X _7576_/Y vssd1 vssd1 vccd1 vccd1 _7578_/B sky130_fd_sc_hd__o22a_1
XFILLER_118_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6528_ _6540_/A vssd1 vssd1 vccd1 vccd1 _6528_/X sky130_fd_sc_hd__buf_1
XFILLER_107_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6459_ _8535_/Q vssd1 vssd1 vccd1 vccd1 _6462_/A sky130_fd_sc_hd__inv_2
XFILLER_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8129_ _8129_/CLK _8129_/D vssd1 vssd1 vccd1 vccd1 _8129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3456_ clkbuf_0__3456_/X vssd1 vssd1 vccd1 vccd1 _7088__525/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6561__252 _6563__254/A vssd1 vssd1 vccd1 vccd1 _7930_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5830_ _5830_/A vssd1 vssd1 vccd1 vccd1 _7827_/D sky130_fd_sc_hd__clkbuf_1
X_6299__201 _6299__201/A vssd1 vssd1 vccd1 vccd1 _7831_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761_ _7905_/Q _5566_/A _5761_/S vssd1 vssd1 vccd1 vccd1 _5762_/A sky130_fd_sc_hd__mux2_1
X_7500_ _8459_/Q vssd1 vssd1 vccd1 vccd1 _7550_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_8480_ _8480_/CLK _8480_/D vssd1 vssd1 vccd1 vccd1 _8480_/Q sky130_fd_sc_hd__dfxtp_1
X_4712_ _4712_/A vssd1 vssd1 vccd1 vccd1 _4712_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5692_ _5692_/A vssd1 vssd1 vccd1 vccd1 _7936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4643_ _4677_/S vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__clkbuf_2
X_4574_ _4574_/A vssd1 vssd1 vccd1 vccd1 _8210_/D sky130_fd_sc_hd__clkbuf_1
X_7362_ _8361_/Q _7286_/A _7357_/X _7361_/Y vssd1 vssd1 vccd1 vccd1 _8361_/D sky130_fd_sc_hd__a31o_1
XFILLER_116_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__3025_ clkbuf_0__3025_/X vssd1 vssd1 vccd1 vccd1 _6175__183/A sky130_fd_sc_hd__clkbuf_4
X_6244_ _8019_/Q _6238_/X _6202_/A _6239_/X _7808_/Q vssd1 vssd1 vccd1 vccd1 _7808_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5126_ _5123_/X _5124_/X _5205_/S vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3310_ clkbuf_0__3310_/X vssd1 vssd1 vccd1 vccd1 _6733__332/A sky130_fd_sc_hd__clkbuf_4
X_5057_ _5252_/S vssd1 vssd1 vccd1 vccd1 _5231_/S sky130_fd_sc_hd__clkbuf_4
X_4008_ _4005_/X _8442_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4009_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5959_ _5959_/A _5965_/B vssd1 vssd1 vccd1 vccd1 _5960_/A sky130_fd_sc_hd__or2_1
XFILLER_111_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6874__373 _6876__375/A vssd1 vssd1 vccd1 vccd1 _8087_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6915__392 _6918__395/A vssd1 vssd1 vccd1 vccd1 _8114_/CLK sky130_fd_sc_hd__inv_2
X_7629_ _8487_/Q _7601_/X vssd1 vssd1 vccd1 vccd1 _7629_/X sky130_fd_sc_hd__or2b_1
XFILLER_119_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3439_ clkbuf_0__3439_/X vssd1 vssd1 vccd1 vccd1 _6998__454/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4290_ _4289_/X _8320_/Q _4290_/S vssd1 vssd1 vccd1 vccd1 _4291_/A sky130_fd_sc_hd__mux2_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7980_ _7980_/CLK _7980_/D vssd1 vssd1 vccd1 vccd1 _7980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__3643_ clkbuf_0__3643_/X vssd1 vssd1 vccd1 vccd1 _7425__145/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6862_ _7614_/A vssd1 vssd1 vccd1 vccd1 _7613_/A sky130_fd_sc_hd__clkbuf_2
X_5813_ _3969_/X _7834_/Q _5815_/S vssd1 vssd1 vccd1 vccd1 _5814_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3574_ clkbuf_0__3574_/X vssd1 vssd1 vccd1 vccd1 _7293__110/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6793_ _7528_/A _6793_/B vssd1 vssd1 vccd1 vccd1 _6808_/A sky130_fd_sc_hd__xor2_1
X_8532_ _8548_/CLK _8532_/D vssd1 vssd1 vccd1 vccd1 _8532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5744_ _5744_/A vssd1 vssd1 vccd1 vccd1 _7913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5675_ _5572_/X _7943_/Q _5677_/S vssd1 vssd1 vccd1 vccd1 _5676_/A sky130_fd_sc_hd__mux2_1
X_8463_ _8487_/CLK _8463_/D vssd1 vssd1 vccd1 vccd1 _8463_/Q sky130_fd_sc_hd__dfxtp_1
X_8394_ _8394_/CLK _8394_/D vssd1 vssd1 vccd1 vccd1 _8394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7414_ _7420_/A vssd1 vssd1 vccd1 vccd1 _7414_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3473_ _7165_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3473_/X sky130_fd_sc_hd__clkbuf_16
X_4626_ _4217_/B _4810_/S _4125_/A vssd1 vssd1 vccd1 vccd1 _4627_/D sky130_fd_sc_hd__a21oi_1
X_7345_ _8357_/Q _7334_/X _7310_/A _7344_/Y vssd1 vssd1 vccd1 vccd1 _7346_/B sky130_fd_sc_hd__o2bb2a_1
X_4557_ _4432_/X _8217_/Q _4559_/S vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4488_ _8245_/Q _4487_/X _4488_/S vssd1 vssd1 vccd1 vccd1 _4489_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7276_ _7234_/Y _7235_/X _7261_/B _7514_/A _7262_/B vssd1 vssd1 vccd1 vccd1 _7277_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6227_ _6272_/A vssd1 vssd1 vccd1 vccd1 _6227_/X sky130_fd_sc_hd__clkbuf_2
X_6568__258 _6568__258/A vssd1 vssd1 vccd1 vccd1 _7936_/CLK sky130_fd_sc_hd__inv_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6247_/A vssd1 vssd1 vccd1 vccd1 _6466_/A sky130_fd_sc_hd__buf_2
XFILLER_111_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5109_/A vssd1 vssd1 vccd1 vccd1 _6941_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_73_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6089_ _6138_/A vssd1 vssd1 vccd1 vccd1 _6105_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3086_ clkbuf_0__3086_/X vssd1 vssd1 vccd1 vccd1 _6296__200/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7098__532 _7099__533/A vssd1 vssd1 vccd1 vccd1 _8259_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5460_ _8066_/Q _4193_/X _5462_/S vssd1 vssd1 vccd1 vccd1 _5461_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4411_ _4411_/A vssd1 vssd1 vccd1 vccd1 _8272_/D sky130_fd_sc_hd__clkbuf_1
X_5391_ _5408_/S vssd1 vssd1 vccd1 vccd1 _5402_/S sky130_fd_sc_hd__buf_2
XFILLER_98_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4342_ _4280_/X _8299_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4343_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4273_ _8325_/Q _4196_/X _4273_/S vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6012_ _6012_/A vssd1 vssd1 vccd1 vccd1 _6012_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
.ends

